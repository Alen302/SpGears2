// Generator : SpinalHDL v1.7.0b    git head : 541894e01cf6b5ef03f924225e4f769fb167dea8
// Component : arraySlice
// Git hash  : c54a5c8a6bc169e2fb8b3189591cb8f780d9540c

`timescale 1ns/1ps

module arraySlice (
  input               inputStreamArrayData_valid,
  output reg          inputStreamArrayData_ready,
  input      [31:0]   inputStreamArrayData_payload,
  input      [6:0]    inputFeatureMapWidth,
  input      [6:0]    inputFeatureMapHeight,
  input      [3:0]    outputFeatureMapHeight,
  input      [3:0]    outputFeatureMapWidth,
  output reg          outputStreamArrayData_0_valid,
  input               outputStreamArrayData_0_ready,
  output reg [31:0]   outputStreamArrayData_0_payload,
  output reg          outputStreamArrayData_1_valid,
  input               outputStreamArrayData_1_ready,
  output reg [31:0]   outputStreamArrayData_1_payload,
  output reg          outputStreamArrayData_2_valid,
  input               outputStreamArrayData_2_ready,
  output reg [31:0]   outputStreamArrayData_2_payload,
  output reg          outputStreamArrayData_3_valid,
  input               outputStreamArrayData_3_ready,
  output reg [31:0]   outputStreamArrayData_3_payload,
  output reg          outputStreamArrayData_4_valid,
  input               outputStreamArrayData_4_ready,
  output reg [31:0]   outputStreamArrayData_4_payload,
  output reg          outputStreamArrayData_5_valid,
  input               outputStreamArrayData_5_ready,
  output reg [31:0]   outputStreamArrayData_5_payload,
  output reg          outputStreamArrayData_6_valid,
  input               outputStreamArrayData_6_ready,
  output reg [31:0]   outputStreamArrayData_6_payload,
  output reg          outputStreamArrayData_7_valid,
  input               outputStreamArrayData_7_ready,
  output reg [31:0]   outputStreamArrayData_7_payload,
  input               clk,
  input               resetn
);
  localparam arraySliceStateMachine_enumDef_BOOT = 2'd0;
  localparam arraySliceStateMachine_enumDef_writeDataOnly = 2'd1;
  localparam arraySliceStateMachine_enumDef_readDataOnly = 2'd2;
  localparam arraySliceStateMachine_enumDef_readWriteData = 2'd3;

  reg                 fifoGroup_0_io_push_valid;
  reg        [31:0]   fifoGroup_0_io_push_payload;
  reg                 fifoGroup_0_io_pop_ready;
  reg                 fifoGroup_1_io_push_valid;
  reg        [31:0]   fifoGroup_1_io_push_payload;
  reg                 fifoGroup_1_io_pop_ready;
  reg                 fifoGroup_2_io_push_valid;
  reg        [31:0]   fifoGroup_2_io_push_payload;
  reg                 fifoGroup_2_io_pop_ready;
  reg                 fifoGroup_3_io_push_valid;
  reg        [31:0]   fifoGroup_3_io_push_payload;
  reg                 fifoGroup_3_io_pop_ready;
  reg                 fifoGroup_4_io_push_valid;
  reg        [31:0]   fifoGroup_4_io_push_payload;
  reg                 fifoGroup_4_io_pop_ready;
  reg                 fifoGroup_5_io_push_valid;
  reg        [31:0]   fifoGroup_5_io_push_payload;
  reg                 fifoGroup_5_io_pop_ready;
  reg                 fifoGroup_6_io_push_valid;
  reg        [31:0]   fifoGroup_6_io_push_payload;
  reg                 fifoGroup_6_io_pop_ready;
  reg                 fifoGroup_7_io_push_valid;
  reg        [31:0]   fifoGroup_7_io_push_payload;
  reg                 fifoGroup_7_io_pop_ready;
  reg                 fifoGroup_8_io_push_valid;
  reg        [31:0]   fifoGroup_8_io_push_payload;
  reg                 fifoGroup_8_io_pop_ready;
  reg                 fifoGroup_9_io_push_valid;
  reg        [31:0]   fifoGroup_9_io_push_payload;
  reg                 fifoGroup_9_io_pop_ready;
  reg                 fifoGroup_10_io_push_valid;
  reg        [31:0]   fifoGroup_10_io_push_payload;
  reg                 fifoGroup_10_io_pop_ready;
  reg                 fifoGroup_11_io_push_valid;
  reg        [31:0]   fifoGroup_11_io_push_payload;
  reg                 fifoGroup_11_io_pop_ready;
  reg                 fifoGroup_12_io_push_valid;
  reg        [31:0]   fifoGroup_12_io_push_payload;
  reg                 fifoGroup_12_io_pop_ready;
  reg                 fifoGroup_13_io_push_valid;
  reg        [31:0]   fifoGroup_13_io_push_payload;
  reg                 fifoGroup_13_io_pop_ready;
  reg                 fifoGroup_14_io_push_valid;
  reg        [31:0]   fifoGroup_14_io_push_payload;
  reg                 fifoGroup_14_io_pop_ready;
  reg                 fifoGroup_15_io_push_valid;
  reg        [31:0]   fifoGroup_15_io_push_payload;
  reg                 fifoGroup_15_io_pop_ready;
  reg                 fifoGroup_16_io_push_valid;
  reg        [31:0]   fifoGroup_16_io_push_payload;
  reg                 fifoGroup_16_io_pop_ready;
  reg                 fifoGroup_17_io_push_valid;
  reg        [31:0]   fifoGroup_17_io_push_payload;
  reg                 fifoGroup_17_io_pop_ready;
  reg                 fifoGroup_18_io_push_valid;
  reg        [31:0]   fifoGroup_18_io_push_payload;
  reg                 fifoGroup_18_io_pop_ready;
  reg                 fifoGroup_19_io_push_valid;
  reg        [31:0]   fifoGroup_19_io_push_payload;
  reg                 fifoGroup_19_io_pop_ready;
  reg                 fifoGroup_20_io_push_valid;
  reg        [31:0]   fifoGroup_20_io_push_payload;
  reg                 fifoGroup_20_io_pop_ready;
  reg                 fifoGroup_21_io_push_valid;
  reg        [31:0]   fifoGroup_21_io_push_payload;
  reg                 fifoGroup_21_io_pop_ready;
  reg                 fifoGroup_22_io_push_valid;
  reg        [31:0]   fifoGroup_22_io_push_payload;
  reg                 fifoGroup_22_io_pop_ready;
  reg                 fifoGroup_23_io_push_valid;
  reg        [31:0]   fifoGroup_23_io_push_payload;
  reg                 fifoGroup_23_io_pop_ready;
  reg                 fifoGroup_24_io_push_valid;
  reg        [31:0]   fifoGroup_24_io_push_payload;
  reg                 fifoGroup_24_io_pop_ready;
  reg                 fifoGroup_25_io_push_valid;
  reg        [31:0]   fifoGroup_25_io_push_payload;
  reg                 fifoGroup_25_io_pop_ready;
  reg                 fifoGroup_26_io_push_valid;
  reg        [31:0]   fifoGroup_26_io_push_payload;
  reg                 fifoGroup_26_io_pop_ready;
  reg                 fifoGroup_27_io_push_valid;
  reg        [31:0]   fifoGroup_27_io_push_payload;
  reg                 fifoGroup_27_io_pop_ready;
  reg                 fifoGroup_28_io_push_valid;
  reg        [31:0]   fifoGroup_28_io_push_payload;
  reg                 fifoGroup_28_io_pop_ready;
  reg                 fifoGroup_29_io_push_valid;
  reg        [31:0]   fifoGroup_29_io_push_payload;
  reg                 fifoGroup_29_io_pop_ready;
  reg                 fifoGroup_30_io_push_valid;
  reg        [31:0]   fifoGroup_30_io_push_payload;
  reg                 fifoGroup_30_io_pop_ready;
  reg                 fifoGroup_31_io_push_valid;
  reg        [31:0]   fifoGroup_31_io_push_payload;
  reg                 fifoGroup_31_io_pop_ready;
  reg                 fifoGroup_32_io_push_valid;
  reg        [31:0]   fifoGroup_32_io_push_payload;
  reg                 fifoGroup_32_io_pop_ready;
  reg                 fifoGroup_33_io_push_valid;
  reg        [31:0]   fifoGroup_33_io_push_payload;
  reg                 fifoGroup_33_io_pop_ready;
  reg                 fifoGroup_34_io_push_valid;
  reg        [31:0]   fifoGroup_34_io_push_payload;
  reg                 fifoGroup_34_io_pop_ready;
  reg                 fifoGroup_35_io_push_valid;
  reg        [31:0]   fifoGroup_35_io_push_payload;
  reg                 fifoGroup_35_io_pop_ready;
  reg                 fifoGroup_36_io_push_valid;
  reg        [31:0]   fifoGroup_36_io_push_payload;
  reg                 fifoGroup_36_io_pop_ready;
  reg                 fifoGroup_37_io_push_valid;
  reg        [31:0]   fifoGroup_37_io_push_payload;
  reg                 fifoGroup_37_io_pop_ready;
  reg                 fifoGroup_38_io_push_valid;
  reg        [31:0]   fifoGroup_38_io_push_payload;
  reg                 fifoGroup_38_io_pop_ready;
  reg                 fifoGroup_39_io_push_valid;
  reg        [31:0]   fifoGroup_39_io_push_payload;
  reg                 fifoGroup_39_io_pop_ready;
  reg                 fifoGroup_40_io_push_valid;
  reg        [31:0]   fifoGroup_40_io_push_payload;
  reg                 fifoGroup_40_io_pop_ready;
  reg                 fifoGroup_41_io_push_valid;
  reg        [31:0]   fifoGroup_41_io_push_payload;
  reg                 fifoGroup_41_io_pop_ready;
  reg                 fifoGroup_42_io_push_valid;
  reg        [31:0]   fifoGroup_42_io_push_payload;
  reg                 fifoGroup_42_io_pop_ready;
  reg                 fifoGroup_43_io_push_valid;
  reg        [31:0]   fifoGroup_43_io_push_payload;
  reg                 fifoGroup_43_io_pop_ready;
  reg                 fifoGroup_44_io_push_valid;
  reg        [31:0]   fifoGroup_44_io_push_payload;
  reg                 fifoGroup_44_io_pop_ready;
  reg                 fifoGroup_45_io_push_valid;
  reg        [31:0]   fifoGroup_45_io_push_payload;
  reg                 fifoGroup_45_io_pop_ready;
  reg                 fifoGroup_46_io_push_valid;
  reg        [31:0]   fifoGroup_46_io_push_payload;
  reg                 fifoGroup_46_io_pop_ready;
  reg                 fifoGroup_47_io_push_valid;
  reg        [31:0]   fifoGroup_47_io_push_payload;
  reg                 fifoGroup_47_io_pop_ready;
  reg                 fifoGroup_48_io_push_valid;
  reg        [31:0]   fifoGroup_48_io_push_payload;
  reg                 fifoGroup_48_io_pop_ready;
  reg                 fifoGroup_49_io_push_valid;
  reg        [31:0]   fifoGroup_49_io_push_payload;
  reg                 fifoGroup_49_io_pop_ready;
  reg                 fifoGroup_50_io_push_valid;
  reg        [31:0]   fifoGroup_50_io_push_payload;
  reg                 fifoGroup_50_io_pop_ready;
  reg                 fifoGroup_51_io_push_valid;
  reg        [31:0]   fifoGroup_51_io_push_payload;
  reg                 fifoGroup_51_io_pop_ready;
  reg                 fifoGroup_52_io_push_valid;
  reg        [31:0]   fifoGroup_52_io_push_payload;
  reg                 fifoGroup_52_io_pop_ready;
  reg                 fifoGroup_53_io_push_valid;
  reg        [31:0]   fifoGroup_53_io_push_payload;
  reg                 fifoGroup_53_io_pop_ready;
  reg                 fifoGroup_54_io_push_valid;
  reg        [31:0]   fifoGroup_54_io_push_payload;
  reg                 fifoGroup_54_io_pop_ready;
  reg                 fifoGroup_55_io_push_valid;
  reg        [31:0]   fifoGroup_55_io_push_payload;
  reg                 fifoGroup_55_io_pop_ready;
  reg                 fifoGroup_56_io_push_valid;
  reg        [31:0]   fifoGroup_56_io_push_payload;
  reg                 fifoGroup_56_io_pop_ready;
  reg                 fifoGroup_57_io_push_valid;
  reg        [31:0]   fifoGroup_57_io_push_payload;
  reg                 fifoGroup_57_io_pop_ready;
  reg                 fifoGroup_58_io_push_valid;
  reg        [31:0]   fifoGroup_58_io_push_payload;
  reg                 fifoGroup_58_io_pop_ready;
  reg                 fifoGroup_59_io_push_valid;
  reg        [31:0]   fifoGroup_59_io_push_payload;
  reg                 fifoGroup_59_io_pop_ready;
  reg                 fifoGroup_60_io_push_valid;
  reg        [31:0]   fifoGroup_60_io_push_payload;
  reg                 fifoGroup_60_io_pop_ready;
  reg                 fifoGroup_61_io_push_valid;
  reg        [31:0]   fifoGroup_61_io_push_payload;
  reg                 fifoGroup_61_io_pop_ready;
  reg                 fifoGroup_62_io_push_valid;
  reg        [31:0]   fifoGroup_62_io_push_payload;
  reg                 fifoGroup_62_io_pop_ready;
  reg                 fifoGroup_63_io_push_valid;
  reg        [31:0]   fifoGroup_63_io_push_payload;
  reg                 fifoGroup_63_io_pop_ready;
  reg                 fifoGroup_64_io_push_valid;
  reg        [31:0]   fifoGroup_64_io_push_payload;
  reg                 fifoGroup_64_io_pop_ready;
  reg                 fifoGroup_65_io_push_valid;
  reg        [31:0]   fifoGroup_65_io_push_payload;
  reg                 fifoGroup_65_io_pop_ready;
  reg                 fifoGroup_66_io_push_valid;
  reg        [31:0]   fifoGroup_66_io_push_payload;
  reg                 fifoGroup_66_io_pop_ready;
  reg                 fifoGroup_67_io_push_valid;
  reg        [31:0]   fifoGroup_67_io_push_payload;
  reg                 fifoGroup_67_io_pop_ready;
  reg                 fifoGroup_68_io_push_valid;
  reg        [31:0]   fifoGroup_68_io_push_payload;
  reg                 fifoGroup_68_io_pop_ready;
  reg                 fifoGroup_69_io_push_valid;
  reg        [31:0]   fifoGroup_69_io_push_payload;
  reg                 fifoGroup_69_io_pop_ready;
  reg                 fifoGroup_70_io_push_valid;
  reg        [31:0]   fifoGroup_70_io_push_payload;
  reg                 fifoGroup_70_io_pop_ready;
  reg                 fifoGroup_71_io_push_valid;
  reg        [31:0]   fifoGroup_71_io_push_payload;
  reg                 fifoGroup_71_io_pop_ready;
  reg                 fifoGroup_72_io_push_valid;
  reg        [31:0]   fifoGroup_72_io_push_payload;
  reg                 fifoGroup_72_io_pop_ready;
  reg                 fifoGroup_73_io_push_valid;
  reg        [31:0]   fifoGroup_73_io_push_payload;
  reg                 fifoGroup_73_io_pop_ready;
  reg                 fifoGroup_74_io_push_valid;
  reg        [31:0]   fifoGroup_74_io_push_payload;
  reg                 fifoGroup_74_io_pop_ready;
  reg                 fifoGroup_75_io_push_valid;
  reg        [31:0]   fifoGroup_75_io_push_payload;
  reg                 fifoGroup_75_io_pop_ready;
  reg                 fifoGroup_76_io_push_valid;
  reg        [31:0]   fifoGroup_76_io_push_payload;
  reg                 fifoGroup_76_io_pop_ready;
  reg                 fifoGroup_77_io_push_valid;
  reg        [31:0]   fifoGroup_77_io_push_payload;
  reg                 fifoGroup_77_io_pop_ready;
  reg                 fifoGroup_78_io_push_valid;
  reg        [31:0]   fifoGroup_78_io_push_payload;
  reg                 fifoGroup_78_io_pop_ready;
  reg                 fifoGroup_79_io_push_valid;
  reg        [31:0]   fifoGroup_79_io_push_payload;
  reg                 fifoGroup_79_io_pop_ready;
  reg                 fifoGroup_80_io_push_valid;
  reg        [31:0]   fifoGroup_80_io_push_payload;
  reg                 fifoGroup_80_io_pop_ready;
  reg                 fifoGroup_81_io_push_valid;
  reg        [31:0]   fifoGroup_81_io_push_payload;
  reg                 fifoGroup_81_io_pop_ready;
  reg                 fifoGroup_82_io_push_valid;
  reg        [31:0]   fifoGroup_82_io_push_payload;
  reg                 fifoGroup_82_io_pop_ready;
  reg                 fifoGroup_83_io_push_valid;
  reg        [31:0]   fifoGroup_83_io_push_payload;
  reg                 fifoGroup_83_io_pop_ready;
  reg                 fifoGroup_84_io_push_valid;
  reg        [31:0]   fifoGroup_84_io_push_payload;
  reg                 fifoGroup_84_io_pop_ready;
  reg                 fifoGroup_85_io_push_valid;
  reg        [31:0]   fifoGroup_85_io_push_payload;
  reg                 fifoGroup_85_io_pop_ready;
  reg                 fifoGroup_86_io_push_valid;
  reg        [31:0]   fifoGroup_86_io_push_payload;
  reg                 fifoGroup_86_io_pop_ready;
  reg                 fifoGroup_87_io_push_valid;
  reg        [31:0]   fifoGroup_87_io_push_payload;
  reg                 fifoGroup_87_io_pop_ready;
  reg                 fifoGroup_88_io_push_valid;
  reg        [31:0]   fifoGroup_88_io_push_payload;
  reg                 fifoGroup_88_io_pop_ready;
  reg                 fifoGroup_89_io_push_valid;
  reg        [31:0]   fifoGroup_89_io_push_payload;
  reg                 fifoGroup_89_io_pop_ready;
  reg                 fifoGroup_90_io_push_valid;
  reg        [31:0]   fifoGroup_90_io_push_payload;
  reg                 fifoGroup_90_io_pop_ready;
  reg                 fifoGroup_91_io_push_valid;
  reg        [31:0]   fifoGroup_91_io_push_payload;
  reg                 fifoGroup_91_io_pop_ready;
  reg                 fifoGroup_92_io_push_valid;
  reg        [31:0]   fifoGroup_92_io_push_payload;
  reg                 fifoGroup_92_io_pop_ready;
  reg                 fifoGroup_93_io_push_valid;
  reg        [31:0]   fifoGroup_93_io_push_payload;
  reg                 fifoGroup_93_io_pop_ready;
  reg                 fifoGroup_94_io_push_valid;
  reg        [31:0]   fifoGroup_94_io_push_payload;
  reg                 fifoGroup_94_io_pop_ready;
  reg                 fifoGroup_95_io_push_valid;
  reg        [31:0]   fifoGroup_95_io_push_payload;
  reg                 fifoGroup_95_io_pop_ready;
  reg                 fifoGroup_96_io_push_valid;
  reg        [31:0]   fifoGroup_96_io_push_payload;
  reg                 fifoGroup_96_io_pop_ready;
  reg                 fifoGroup_97_io_push_valid;
  reg        [31:0]   fifoGroup_97_io_push_payload;
  reg                 fifoGroup_97_io_pop_ready;
  reg                 fifoGroup_98_io_push_valid;
  reg        [31:0]   fifoGroup_98_io_push_payload;
  reg                 fifoGroup_98_io_pop_ready;
  reg                 fifoGroup_99_io_push_valid;
  reg        [31:0]   fifoGroup_99_io_push_payload;
  reg                 fifoGroup_99_io_pop_ready;
  reg                 fifoGroup_100_io_push_valid;
  reg        [31:0]   fifoGroup_100_io_push_payload;
  reg                 fifoGroup_100_io_pop_ready;
  reg                 fifoGroup_101_io_push_valid;
  reg        [31:0]   fifoGroup_101_io_push_payload;
  reg                 fifoGroup_101_io_pop_ready;
  reg                 fifoGroup_102_io_push_valid;
  reg        [31:0]   fifoGroup_102_io_push_payload;
  reg                 fifoGroup_102_io_pop_ready;
  reg                 fifoGroup_103_io_push_valid;
  reg        [31:0]   fifoGroup_103_io_push_payload;
  reg                 fifoGroup_103_io_pop_ready;
  reg                 fifoGroup_104_io_push_valid;
  reg        [31:0]   fifoGroup_104_io_push_payload;
  reg                 fifoGroup_104_io_pop_ready;
  reg                 fifoGroup_105_io_push_valid;
  reg        [31:0]   fifoGroup_105_io_push_payload;
  reg                 fifoGroup_105_io_pop_ready;
  reg                 fifoGroup_106_io_push_valid;
  reg        [31:0]   fifoGroup_106_io_push_payload;
  reg                 fifoGroup_106_io_pop_ready;
  reg                 fifoGroup_107_io_push_valid;
  reg        [31:0]   fifoGroup_107_io_push_payload;
  reg                 fifoGroup_107_io_pop_ready;
  reg                 fifoGroup_108_io_push_valid;
  reg        [31:0]   fifoGroup_108_io_push_payload;
  reg                 fifoGroup_108_io_pop_ready;
  reg                 fifoGroup_109_io_push_valid;
  reg        [31:0]   fifoGroup_109_io_push_payload;
  reg                 fifoGroup_109_io_pop_ready;
  wire                fifoGroup_0_io_push_ready;
  wire                fifoGroup_0_io_pop_valid;
  wire       [31:0]   fifoGroup_0_io_pop_payload;
  wire       [6:0]    fifoGroup_0_io_occupancy;
  wire       [6:0]    fifoGroup_0_io_availability;
  wire                fifoGroup_1_io_push_ready;
  wire                fifoGroup_1_io_pop_valid;
  wire       [31:0]   fifoGroup_1_io_pop_payload;
  wire       [6:0]    fifoGroup_1_io_occupancy;
  wire       [6:0]    fifoGroup_1_io_availability;
  wire                fifoGroup_2_io_push_ready;
  wire                fifoGroup_2_io_pop_valid;
  wire       [31:0]   fifoGroup_2_io_pop_payload;
  wire       [6:0]    fifoGroup_2_io_occupancy;
  wire       [6:0]    fifoGroup_2_io_availability;
  wire                fifoGroup_3_io_push_ready;
  wire                fifoGroup_3_io_pop_valid;
  wire       [31:0]   fifoGroup_3_io_pop_payload;
  wire       [6:0]    fifoGroup_3_io_occupancy;
  wire       [6:0]    fifoGroup_3_io_availability;
  wire                fifoGroup_4_io_push_ready;
  wire                fifoGroup_4_io_pop_valid;
  wire       [31:0]   fifoGroup_4_io_pop_payload;
  wire       [6:0]    fifoGroup_4_io_occupancy;
  wire       [6:0]    fifoGroup_4_io_availability;
  wire                fifoGroup_5_io_push_ready;
  wire                fifoGroup_5_io_pop_valid;
  wire       [31:0]   fifoGroup_5_io_pop_payload;
  wire       [6:0]    fifoGroup_5_io_occupancy;
  wire       [6:0]    fifoGroup_5_io_availability;
  wire                fifoGroup_6_io_push_ready;
  wire                fifoGroup_6_io_pop_valid;
  wire       [31:0]   fifoGroup_6_io_pop_payload;
  wire       [6:0]    fifoGroup_6_io_occupancy;
  wire       [6:0]    fifoGroup_6_io_availability;
  wire                fifoGroup_7_io_push_ready;
  wire                fifoGroup_7_io_pop_valid;
  wire       [31:0]   fifoGroup_7_io_pop_payload;
  wire       [6:0]    fifoGroup_7_io_occupancy;
  wire       [6:0]    fifoGroup_7_io_availability;
  wire                fifoGroup_8_io_push_ready;
  wire                fifoGroup_8_io_pop_valid;
  wire       [31:0]   fifoGroup_8_io_pop_payload;
  wire       [6:0]    fifoGroup_8_io_occupancy;
  wire       [6:0]    fifoGroup_8_io_availability;
  wire                fifoGroup_9_io_push_ready;
  wire                fifoGroup_9_io_pop_valid;
  wire       [31:0]   fifoGroup_9_io_pop_payload;
  wire       [6:0]    fifoGroup_9_io_occupancy;
  wire       [6:0]    fifoGroup_9_io_availability;
  wire                fifoGroup_10_io_push_ready;
  wire                fifoGroup_10_io_pop_valid;
  wire       [31:0]   fifoGroup_10_io_pop_payload;
  wire       [6:0]    fifoGroup_10_io_occupancy;
  wire       [6:0]    fifoGroup_10_io_availability;
  wire                fifoGroup_11_io_push_ready;
  wire                fifoGroup_11_io_pop_valid;
  wire       [31:0]   fifoGroup_11_io_pop_payload;
  wire       [6:0]    fifoGroup_11_io_occupancy;
  wire       [6:0]    fifoGroup_11_io_availability;
  wire                fifoGroup_12_io_push_ready;
  wire                fifoGroup_12_io_pop_valid;
  wire       [31:0]   fifoGroup_12_io_pop_payload;
  wire       [6:0]    fifoGroup_12_io_occupancy;
  wire       [6:0]    fifoGroup_12_io_availability;
  wire                fifoGroup_13_io_push_ready;
  wire                fifoGroup_13_io_pop_valid;
  wire       [31:0]   fifoGroup_13_io_pop_payload;
  wire       [6:0]    fifoGroup_13_io_occupancy;
  wire       [6:0]    fifoGroup_13_io_availability;
  wire                fifoGroup_14_io_push_ready;
  wire                fifoGroup_14_io_pop_valid;
  wire       [31:0]   fifoGroup_14_io_pop_payload;
  wire       [6:0]    fifoGroup_14_io_occupancy;
  wire       [6:0]    fifoGroup_14_io_availability;
  wire                fifoGroup_15_io_push_ready;
  wire                fifoGroup_15_io_pop_valid;
  wire       [31:0]   fifoGroup_15_io_pop_payload;
  wire       [6:0]    fifoGroup_15_io_occupancy;
  wire       [6:0]    fifoGroup_15_io_availability;
  wire                fifoGroup_16_io_push_ready;
  wire                fifoGroup_16_io_pop_valid;
  wire       [31:0]   fifoGroup_16_io_pop_payload;
  wire       [6:0]    fifoGroup_16_io_occupancy;
  wire       [6:0]    fifoGroup_16_io_availability;
  wire                fifoGroup_17_io_push_ready;
  wire                fifoGroup_17_io_pop_valid;
  wire       [31:0]   fifoGroup_17_io_pop_payload;
  wire       [6:0]    fifoGroup_17_io_occupancy;
  wire       [6:0]    fifoGroup_17_io_availability;
  wire                fifoGroup_18_io_push_ready;
  wire                fifoGroup_18_io_pop_valid;
  wire       [31:0]   fifoGroup_18_io_pop_payload;
  wire       [6:0]    fifoGroup_18_io_occupancy;
  wire       [6:0]    fifoGroup_18_io_availability;
  wire                fifoGroup_19_io_push_ready;
  wire                fifoGroup_19_io_pop_valid;
  wire       [31:0]   fifoGroup_19_io_pop_payload;
  wire       [6:0]    fifoGroup_19_io_occupancy;
  wire       [6:0]    fifoGroup_19_io_availability;
  wire                fifoGroup_20_io_push_ready;
  wire                fifoGroup_20_io_pop_valid;
  wire       [31:0]   fifoGroup_20_io_pop_payload;
  wire       [6:0]    fifoGroup_20_io_occupancy;
  wire       [6:0]    fifoGroup_20_io_availability;
  wire                fifoGroup_21_io_push_ready;
  wire                fifoGroup_21_io_pop_valid;
  wire       [31:0]   fifoGroup_21_io_pop_payload;
  wire       [6:0]    fifoGroup_21_io_occupancy;
  wire       [6:0]    fifoGroup_21_io_availability;
  wire                fifoGroup_22_io_push_ready;
  wire                fifoGroup_22_io_pop_valid;
  wire       [31:0]   fifoGroup_22_io_pop_payload;
  wire       [6:0]    fifoGroup_22_io_occupancy;
  wire       [6:0]    fifoGroup_22_io_availability;
  wire                fifoGroup_23_io_push_ready;
  wire                fifoGroup_23_io_pop_valid;
  wire       [31:0]   fifoGroup_23_io_pop_payload;
  wire       [6:0]    fifoGroup_23_io_occupancy;
  wire       [6:0]    fifoGroup_23_io_availability;
  wire                fifoGroup_24_io_push_ready;
  wire                fifoGroup_24_io_pop_valid;
  wire       [31:0]   fifoGroup_24_io_pop_payload;
  wire       [6:0]    fifoGroup_24_io_occupancy;
  wire       [6:0]    fifoGroup_24_io_availability;
  wire                fifoGroup_25_io_push_ready;
  wire                fifoGroup_25_io_pop_valid;
  wire       [31:0]   fifoGroup_25_io_pop_payload;
  wire       [6:0]    fifoGroup_25_io_occupancy;
  wire       [6:0]    fifoGroup_25_io_availability;
  wire                fifoGroup_26_io_push_ready;
  wire                fifoGroup_26_io_pop_valid;
  wire       [31:0]   fifoGroup_26_io_pop_payload;
  wire       [6:0]    fifoGroup_26_io_occupancy;
  wire       [6:0]    fifoGroup_26_io_availability;
  wire                fifoGroup_27_io_push_ready;
  wire                fifoGroup_27_io_pop_valid;
  wire       [31:0]   fifoGroup_27_io_pop_payload;
  wire       [6:0]    fifoGroup_27_io_occupancy;
  wire       [6:0]    fifoGroup_27_io_availability;
  wire                fifoGroup_28_io_push_ready;
  wire                fifoGroup_28_io_pop_valid;
  wire       [31:0]   fifoGroup_28_io_pop_payload;
  wire       [6:0]    fifoGroup_28_io_occupancy;
  wire       [6:0]    fifoGroup_28_io_availability;
  wire                fifoGroup_29_io_push_ready;
  wire                fifoGroup_29_io_pop_valid;
  wire       [31:0]   fifoGroup_29_io_pop_payload;
  wire       [6:0]    fifoGroup_29_io_occupancy;
  wire       [6:0]    fifoGroup_29_io_availability;
  wire                fifoGroup_30_io_push_ready;
  wire                fifoGroup_30_io_pop_valid;
  wire       [31:0]   fifoGroup_30_io_pop_payload;
  wire       [6:0]    fifoGroup_30_io_occupancy;
  wire       [6:0]    fifoGroup_30_io_availability;
  wire                fifoGroup_31_io_push_ready;
  wire                fifoGroup_31_io_pop_valid;
  wire       [31:0]   fifoGroup_31_io_pop_payload;
  wire       [6:0]    fifoGroup_31_io_occupancy;
  wire       [6:0]    fifoGroup_31_io_availability;
  wire                fifoGroup_32_io_push_ready;
  wire                fifoGroup_32_io_pop_valid;
  wire       [31:0]   fifoGroup_32_io_pop_payload;
  wire       [6:0]    fifoGroup_32_io_occupancy;
  wire       [6:0]    fifoGroup_32_io_availability;
  wire                fifoGroup_33_io_push_ready;
  wire                fifoGroup_33_io_pop_valid;
  wire       [31:0]   fifoGroup_33_io_pop_payload;
  wire       [6:0]    fifoGroup_33_io_occupancy;
  wire       [6:0]    fifoGroup_33_io_availability;
  wire                fifoGroup_34_io_push_ready;
  wire                fifoGroup_34_io_pop_valid;
  wire       [31:0]   fifoGroup_34_io_pop_payload;
  wire       [6:0]    fifoGroup_34_io_occupancy;
  wire       [6:0]    fifoGroup_34_io_availability;
  wire                fifoGroup_35_io_push_ready;
  wire                fifoGroup_35_io_pop_valid;
  wire       [31:0]   fifoGroup_35_io_pop_payload;
  wire       [6:0]    fifoGroup_35_io_occupancy;
  wire       [6:0]    fifoGroup_35_io_availability;
  wire                fifoGroup_36_io_push_ready;
  wire                fifoGroup_36_io_pop_valid;
  wire       [31:0]   fifoGroup_36_io_pop_payload;
  wire       [6:0]    fifoGroup_36_io_occupancy;
  wire       [6:0]    fifoGroup_36_io_availability;
  wire                fifoGroup_37_io_push_ready;
  wire                fifoGroup_37_io_pop_valid;
  wire       [31:0]   fifoGroup_37_io_pop_payload;
  wire       [6:0]    fifoGroup_37_io_occupancy;
  wire       [6:0]    fifoGroup_37_io_availability;
  wire                fifoGroup_38_io_push_ready;
  wire                fifoGroup_38_io_pop_valid;
  wire       [31:0]   fifoGroup_38_io_pop_payload;
  wire       [6:0]    fifoGroup_38_io_occupancy;
  wire       [6:0]    fifoGroup_38_io_availability;
  wire                fifoGroup_39_io_push_ready;
  wire                fifoGroup_39_io_pop_valid;
  wire       [31:0]   fifoGroup_39_io_pop_payload;
  wire       [6:0]    fifoGroup_39_io_occupancy;
  wire       [6:0]    fifoGroup_39_io_availability;
  wire                fifoGroup_40_io_push_ready;
  wire                fifoGroup_40_io_pop_valid;
  wire       [31:0]   fifoGroup_40_io_pop_payload;
  wire       [6:0]    fifoGroup_40_io_occupancy;
  wire       [6:0]    fifoGroup_40_io_availability;
  wire                fifoGroup_41_io_push_ready;
  wire                fifoGroup_41_io_pop_valid;
  wire       [31:0]   fifoGroup_41_io_pop_payload;
  wire       [6:0]    fifoGroup_41_io_occupancy;
  wire       [6:0]    fifoGroup_41_io_availability;
  wire                fifoGroup_42_io_push_ready;
  wire                fifoGroup_42_io_pop_valid;
  wire       [31:0]   fifoGroup_42_io_pop_payload;
  wire       [6:0]    fifoGroup_42_io_occupancy;
  wire       [6:0]    fifoGroup_42_io_availability;
  wire                fifoGroup_43_io_push_ready;
  wire                fifoGroup_43_io_pop_valid;
  wire       [31:0]   fifoGroup_43_io_pop_payload;
  wire       [6:0]    fifoGroup_43_io_occupancy;
  wire       [6:0]    fifoGroup_43_io_availability;
  wire                fifoGroup_44_io_push_ready;
  wire                fifoGroup_44_io_pop_valid;
  wire       [31:0]   fifoGroup_44_io_pop_payload;
  wire       [6:0]    fifoGroup_44_io_occupancy;
  wire       [6:0]    fifoGroup_44_io_availability;
  wire                fifoGroup_45_io_push_ready;
  wire                fifoGroup_45_io_pop_valid;
  wire       [31:0]   fifoGroup_45_io_pop_payload;
  wire       [6:0]    fifoGroup_45_io_occupancy;
  wire       [6:0]    fifoGroup_45_io_availability;
  wire                fifoGroup_46_io_push_ready;
  wire                fifoGroup_46_io_pop_valid;
  wire       [31:0]   fifoGroup_46_io_pop_payload;
  wire       [6:0]    fifoGroup_46_io_occupancy;
  wire       [6:0]    fifoGroup_46_io_availability;
  wire                fifoGroup_47_io_push_ready;
  wire                fifoGroup_47_io_pop_valid;
  wire       [31:0]   fifoGroup_47_io_pop_payload;
  wire       [6:0]    fifoGroup_47_io_occupancy;
  wire       [6:0]    fifoGroup_47_io_availability;
  wire                fifoGroup_48_io_push_ready;
  wire                fifoGroup_48_io_pop_valid;
  wire       [31:0]   fifoGroup_48_io_pop_payload;
  wire       [6:0]    fifoGroup_48_io_occupancy;
  wire       [6:0]    fifoGroup_48_io_availability;
  wire                fifoGroup_49_io_push_ready;
  wire                fifoGroup_49_io_pop_valid;
  wire       [31:0]   fifoGroup_49_io_pop_payload;
  wire       [6:0]    fifoGroup_49_io_occupancy;
  wire       [6:0]    fifoGroup_49_io_availability;
  wire                fifoGroup_50_io_push_ready;
  wire                fifoGroup_50_io_pop_valid;
  wire       [31:0]   fifoGroup_50_io_pop_payload;
  wire       [6:0]    fifoGroup_50_io_occupancy;
  wire       [6:0]    fifoGroup_50_io_availability;
  wire                fifoGroup_51_io_push_ready;
  wire                fifoGroup_51_io_pop_valid;
  wire       [31:0]   fifoGroup_51_io_pop_payload;
  wire       [6:0]    fifoGroup_51_io_occupancy;
  wire       [6:0]    fifoGroup_51_io_availability;
  wire                fifoGroup_52_io_push_ready;
  wire                fifoGroup_52_io_pop_valid;
  wire       [31:0]   fifoGroup_52_io_pop_payload;
  wire       [6:0]    fifoGroup_52_io_occupancy;
  wire       [6:0]    fifoGroup_52_io_availability;
  wire                fifoGroup_53_io_push_ready;
  wire                fifoGroup_53_io_pop_valid;
  wire       [31:0]   fifoGroup_53_io_pop_payload;
  wire       [6:0]    fifoGroup_53_io_occupancy;
  wire       [6:0]    fifoGroup_53_io_availability;
  wire                fifoGroup_54_io_push_ready;
  wire                fifoGroup_54_io_pop_valid;
  wire       [31:0]   fifoGroup_54_io_pop_payload;
  wire       [6:0]    fifoGroup_54_io_occupancy;
  wire       [6:0]    fifoGroup_54_io_availability;
  wire                fifoGroup_55_io_push_ready;
  wire                fifoGroup_55_io_pop_valid;
  wire       [31:0]   fifoGroup_55_io_pop_payload;
  wire       [6:0]    fifoGroup_55_io_occupancy;
  wire       [6:0]    fifoGroup_55_io_availability;
  wire                fifoGroup_56_io_push_ready;
  wire                fifoGroup_56_io_pop_valid;
  wire       [31:0]   fifoGroup_56_io_pop_payload;
  wire       [6:0]    fifoGroup_56_io_occupancy;
  wire       [6:0]    fifoGroup_56_io_availability;
  wire                fifoGroup_57_io_push_ready;
  wire                fifoGroup_57_io_pop_valid;
  wire       [31:0]   fifoGroup_57_io_pop_payload;
  wire       [6:0]    fifoGroup_57_io_occupancy;
  wire       [6:0]    fifoGroup_57_io_availability;
  wire                fifoGroup_58_io_push_ready;
  wire                fifoGroup_58_io_pop_valid;
  wire       [31:0]   fifoGroup_58_io_pop_payload;
  wire       [6:0]    fifoGroup_58_io_occupancy;
  wire       [6:0]    fifoGroup_58_io_availability;
  wire                fifoGroup_59_io_push_ready;
  wire                fifoGroup_59_io_pop_valid;
  wire       [31:0]   fifoGroup_59_io_pop_payload;
  wire       [6:0]    fifoGroup_59_io_occupancy;
  wire       [6:0]    fifoGroup_59_io_availability;
  wire                fifoGroup_60_io_push_ready;
  wire                fifoGroup_60_io_pop_valid;
  wire       [31:0]   fifoGroup_60_io_pop_payload;
  wire       [6:0]    fifoGroup_60_io_occupancy;
  wire       [6:0]    fifoGroup_60_io_availability;
  wire                fifoGroup_61_io_push_ready;
  wire                fifoGroup_61_io_pop_valid;
  wire       [31:0]   fifoGroup_61_io_pop_payload;
  wire       [6:0]    fifoGroup_61_io_occupancy;
  wire       [6:0]    fifoGroup_61_io_availability;
  wire                fifoGroup_62_io_push_ready;
  wire                fifoGroup_62_io_pop_valid;
  wire       [31:0]   fifoGroup_62_io_pop_payload;
  wire       [6:0]    fifoGroup_62_io_occupancy;
  wire       [6:0]    fifoGroup_62_io_availability;
  wire                fifoGroup_63_io_push_ready;
  wire                fifoGroup_63_io_pop_valid;
  wire       [31:0]   fifoGroup_63_io_pop_payload;
  wire       [6:0]    fifoGroup_63_io_occupancy;
  wire       [6:0]    fifoGroup_63_io_availability;
  wire                fifoGroup_64_io_push_ready;
  wire                fifoGroup_64_io_pop_valid;
  wire       [31:0]   fifoGroup_64_io_pop_payload;
  wire       [6:0]    fifoGroup_64_io_occupancy;
  wire       [6:0]    fifoGroup_64_io_availability;
  wire                fifoGroup_65_io_push_ready;
  wire                fifoGroup_65_io_pop_valid;
  wire       [31:0]   fifoGroup_65_io_pop_payload;
  wire       [6:0]    fifoGroup_65_io_occupancy;
  wire       [6:0]    fifoGroup_65_io_availability;
  wire                fifoGroup_66_io_push_ready;
  wire                fifoGroup_66_io_pop_valid;
  wire       [31:0]   fifoGroup_66_io_pop_payload;
  wire       [6:0]    fifoGroup_66_io_occupancy;
  wire       [6:0]    fifoGroup_66_io_availability;
  wire                fifoGroup_67_io_push_ready;
  wire                fifoGroup_67_io_pop_valid;
  wire       [31:0]   fifoGroup_67_io_pop_payload;
  wire       [6:0]    fifoGroup_67_io_occupancy;
  wire       [6:0]    fifoGroup_67_io_availability;
  wire                fifoGroup_68_io_push_ready;
  wire                fifoGroup_68_io_pop_valid;
  wire       [31:0]   fifoGroup_68_io_pop_payload;
  wire       [6:0]    fifoGroup_68_io_occupancy;
  wire       [6:0]    fifoGroup_68_io_availability;
  wire                fifoGroup_69_io_push_ready;
  wire                fifoGroup_69_io_pop_valid;
  wire       [31:0]   fifoGroup_69_io_pop_payload;
  wire       [6:0]    fifoGroup_69_io_occupancy;
  wire       [6:0]    fifoGroup_69_io_availability;
  wire                fifoGroup_70_io_push_ready;
  wire                fifoGroup_70_io_pop_valid;
  wire       [31:0]   fifoGroup_70_io_pop_payload;
  wire       [6:0]    fifoGroup_70_io_occupancy;
  wire       [6:0]    fifoGroup_70_io_availability;
  wire                fifoGroup_71_io_push_ready;
  wire                fifoGroup_71_io_pop_valid;
  wire       [31:0]   fifoGroup_71_io_pop_payload;
  wire       [6:0]    fifoGroup_71_io_occupancy;
  wire       [6:0]    fifoGroup_71_io_availability;
  wire                fifoGroup_72_io_push_ready;
  wire                fifoGroup_72_io_pop_valid;
  wire       [31:0]   fifoGroup_72_io_pop_payload;
  wire       [6:0]    fifoGroup_72_io_occupancy;
  wire       [6:0]    fifoGroup_72_io_availability;
  wire                fifoGroup_73_io_push_ready;
  wire                fifoGroup_73_io_pop_valid;
  wire       [31:0]   fifoGroup_73_io_pop_payload;
  wire       [6:0]    fifoGroup_73_io_occupancy;
  wire       [6:0]    fifoGroup_73_io_availability;
  wire                fifoGroup_74_io_push_ready;
  wire                fifoGroup_74_io_pop_valid;
  wire       [31:0]   fifoGroup_74_io_pop_payload;
  wire       [6:0]    fifoGroup_74_io_occupancy;
  wire       [6:0]    fifoGroup_74_io_availability;
  wire                fifoGroup_75_io_push_ready;
  wire                fifoGroup_75_io_pop_valid;
  wire       [31:0]   fifoGroup_75_io_pop_payload;
  wire       [6:0]    fifoGroup_75_io_occupancy;
  wire       [6:0]    fifoGroup_75_io_availability;
  wire                fifoGroup_76_io_push_ready;
  wire                fifoGroup_76_io_pop_valid;
  wire       [31:0]   fifoGroup_76_io_pop_payload;
  wire       [6:0]    fifoGroup_76_io_occupancy;
  wire       [6:0]    fifoGroup_76_io_availability;
  wire                fifoGroup_77_io_push_ready;
  wire                fifoGroup_77_io_pop_valid;
  wire       [31:0]   fifoGroup_77_io_pop_payload;
  wire       [6:0]    fifoGroup_77_io_occupancy;
  wire       [6:0]    fifoGroup_77_io_availability;
  wire                fifoGroup_78_io_push_ready;
  wire                fifoGroup_78_io_pop_valid;
  wire       [31:0]   fifoGroup_78_io_pop_payload;
  wire       [6:0]    fifoGroup_78_io_occupancy;
  wire       [6:0]    fifoGroup_78_io_availability;
  wire                fifoGroup_79_io_push_ready;
  wire                fifoGroup_79_io_pop_valid;
  wire       [31:0]   fifoGroup_79_io_pop_payload;
  wire       [6:0]    fifoGroup_79_io_occupancy;
  wire       [6:0]    fifoGroup_79_io_availability;
  wire                fifoGroup_80_io_push_ready;
  wire                fifoGroup_80_io_pop_valid;
  wire       [31:0]   fifoGroup_80_io_pop_payload;
  wire       [6:0]    fifoGroup_80_io_occupancy;
  wire       [6:0]    fifoGroup_80_io_availability;
  wire                fifoGroup_81_io_push_ready;
  wire                fifoGroup_81_io_pop_valid;
  wire       [31:0]   fifoGroup_81_io_pop_payload;
  wire       [6:0]    fifoGroup_81_io_occupancy;
  wire       [6:0]    fifoGroup_81_io_availability;
  wire                fifoGroup_82_io_push_ready;
  wire                fifoGroup_82_io_pop_valid;
  wire       [31:0]   fifoGroup_82_io_pop_payload;
  wire       [6:0]    fifoGroup_82_io_occupancy;
  wire       [6:0]    fifoGroup_82_io_availability;
  wire                fifoGroup_83_io_push_ready;
  wire                fifoGroup_83_io_pop_valid;
  wire       [31:0]   fifoGroup_83_io_pop_payload;
  wire       [6:0]    fifoGroup_83_io_occupancy;
  wire       [6:0]    fifoGroup_83_io_availability;
  wire                fifoGroup_84_io_push_ready;
  wire                fifoGroup_84_io_pop_valid;
  wire       [31:0]   fifoGroup_84_io_pop_payload;
  wire       [6:0]    fifoGroup_84_io_occupancy;
  wire       [6:0]    fifoGroup_84_io_availability;
  wire                fifoGroup_85_io_push_ready;
  wire                fifoGroup_85_io_pop_valid;
  wire       [31:0]   fifoGroup_85_io_pop_payload;
  wire       [6:0]    fifoGroup_85_io_occupancy;
  wire       [6:0]    fifoGroup_85_io_availability;
  wire                fifoGroup_86_io_push_ready;
  wire                fifoGroup_86_io_pop_valid;
  wire       [31:0]   fifoGroup_86_io_pop_payload;
  wire       [6:0]    fifoGroup_86_io_occupancy;
  wire       [6:0]    fifoGroup_86_io_availability;
  wire                fifoGroup_87_io_push_ready;
  wire                fifoGroup_87_io_pop_valid;
  wire       [31:0]   fifoGroup_87_io_pop_payload;
  wire       [6:0]    fifoGroup_87_io_occupancy;
  wire       [6:0]    fifoGroup_87_io_availability;
  wire                fifoGroup_88_io_push_ready;
  wire                fifoGroup_88_io_pop_valid;
  wire       [31:0]   fifoGroup_88_io_pop_payload;
  wire       [6:0]    fifoGroup_88_io_occupancy;
  wire       [6:0]    fifoGroup_88_io_availability;
  wire                fifoGroup_89_io_push_ready;
  wire                fifoGroup_89_io_pop_valid;
  wire       [31:0]   fifoGroup_89_io_pop_payload;
  wire       [6:0]    fifoGroup_89_io_occupancy;
  wire       [6:0]    fifoGroup_89_io_availability;
  wire                fifoGroup_90_io_push_ready;
  wire                fifoGroup_90_io_pop_valid;
  wire       [31:0]   fifoGroup_90_io_pop_payload;
  wire       [6:0]    fifoGroup_90_io_occupancy;
  wire       [6:0]    fifoGroup_90_io_availability;
  wire                fifoGroup_91_io_push_ready;
  wire                fifoGroup_91_io_pop_valid;
  wire       [31:0]   fifoGroup_91_io_pop_payload;
  wire       [6:0]    fifoGroup_91_io_occupancy;
  wire       [6:0]    fifoGroup_91_io_availability;
  wire                fifoGroup_92_io_push_ready;
  wire                fifoGroup_92_io_pop_valid;
  wire       [31:0]   fifoGroup_92_io_pop_payload;
  wire       [6:0]    fifoGroup_92_io_occupancy;
  wire       [6:0]    fifoGroup_92_io_availability;
  wire                fifoGroup_93_io_push_ready;
  wire                fifoGroup_93_io_pop_valid;
  wire       [31:0]   fifoGroup_93_io_pop_payload;
  wire       [6:0]    fifoGroup_93_io_occupancy;
  wire       [6:0]    fifoGroup_93_io_availability;
  wire                fifoGroup_94_io_push_ready;
  wire                fifoGroup_94_io_pop_valid;
  wire       [31:0]   fifoGroup_94_io_pop_payload;
  wire       [6:0]    fifoGroup_94_io_occupancy;
  wire       [6:0]    fifoGroup_94_io_availability;
  wire                fifoGroup_95_io_push_ready;
  wire                fifoGroup_95_io_pop_valid;
  wire       [31:0]   fifoGroup_95_io_pop_payload;
  wire       [6:0]    fifoGroup_95_io_occupancy;
  wire       [6:0]    fifoGroup_95_io_availability;
  wire                fifoGroup_96_io_push_ready;
  wire                fifoGroup_96_io_pop_valid;
  wire       [31:0]   fifoGroup_96_io_pop_payload;
  wire       [6:0]    fifoGroup_96_io_occupancy;
  wire       [6:0]    fifoGroup_96_io_availability;
  wire                fifoGroup_97_io_push_ready;
  wire                fifoGroup_97_io_pop_valid;
  wire       [31:0]   fifoGroup_97_io_pop_payload;
  wire       [6:0]    fifoGroup_97_io_occupancy;
  wire       [6:0]    fifoGroup_97_io_availability;
  wire                fifoGroup_98_io_push_ready;
  wire                fifoGroup_98_io_pop_valid;
  wire       [31:0]   fifoGroup_98_io_pop_payload;
  wire       [6:0]    fifoGroup_98_io_occupancy;
  wire       [6:0]    fifoGroup_98_io_availability;
  wire                fifoGroup_99_io_push_ready;
  wire                fifoGroup_99_io_pop_valid;
  wire       [31:0]   fifoGroup_99_io_pop_payload;
  wire       [6:0]    fifoGroup_99_io_occupancy;
  wire       [6:0]    fifoGroup_99_io_availability;
  wire                fifoGroup_100_io_push_ready;
  wire                fifoGroup_100_io_pop_valid;
  wire       [31:0]   fifoGroup_100_io_pop_payload;
  wire       [6:0]    fifoGroup_100_io_occupancy;
  wire       [6:0]    fifoGroup_100_io_availability;
  wire                fifoGroup_101_io_push_ready;
  wire                fifoGroup_101_io_pop_valid;
  wire       [31:0]   fifoGroup_101_io_pop_payload;
  wire       [6:0]    fifoGroup_101_io_occupancy;
  wire       [6:0]    fifoGroup_101_io_availability;
  wire                fifoGroup_102_io_push_ready;
  wire                fifoGroup_102_io_pop_valid;
  wire       [31:0]   fifoGroup_102_io_pop_payload;
  wire       [6:0]    fifoGroup_102_io_occupancy;
  wire       [6:0]    fifoGroup_102_io_availability;
  wire                fifoGroup_103_io_push_ready;
  wire                fifoGroup_103_io_pop_valid;
  wire       [31:0]   fifoGroup_103_io_pop_payload;
  wire       [6:0]    fifoGroup_103_io_occupancy;
  wire       [6:0]    fifoGroup_103_io_availability;
  wire                fifoGroup_104_io_push_ready;
  wire                fifoGroup_104_io_pop_valid;
  wire       [31:0]   fifoGroup_104_io_pop_payload;
  wire       [6:0]    fifoGroup_104_io_occupancy;
  wire       [6:0]    fifoGroup_104_io_availability;
  wire                fifoGroup_105_io_push_ready;
  wire                fifoGroup_105_io_pop_valid;
  wire       [31:0]   fifoGroup_105_io_pop_payload;
  wire       [6:0]    fifoGroup_105_io_occupancy;
  wire       [6:0]    fifoGroup_105_io_availability;
  wire                fifoGroup_106_io_push_ready;
  wire                fifoGroup_106_io_pop_valid;
  wire       [31:0]   fifoGroup_106_io_pop_payload;
  wire       [6:0]    fifoGroup_106_io_occupancy;
  wire       [6:0]    fifoGroup_106_io_availability;
  wire                fifoGroup_107_io_push_ready;
  wire                fifoGroup_107_io_pop_valid;
  wire       [31:0]   fifoGroup_107_io_pop_payload;
  wire       [6:0]    fifoGroup_107_io_occupancy;
  wire       [6:0]    fifoGroup_107_io_availability;
  wire                fifoGroup_108_io_push_ready;
  wire                fifoGroup_108_io_pop_valid;
  wire       [31:0]   fifoGroup_108_io_pop_payload;
  wire       [6:0]    fifoGroup_108_io_occupancy;
  wire       [6:0]    fifoGroup_108_io_availability;
  wire                fifoGroup_109_io_push_ready;
  wire                fifoGroup_109_io_pop_valid;
  wire       [31:0]   fifoGroup_109_io_pop_payload;
  wire       [6:0]    fifoGroup_109_io_occupancy;
  wire       [6:0]    fifoGroup_109_io_availability;
  wire       [12:0]   _zz_handshakeTimes_0_valueNext;
  wire       [0:0]    _zz_handshakeTimes_0_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_1_valueNext;
  wire       [0:0]    _zz_handshakeTimes_1_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_2_valueNext;
  wire       [0:0]    _zz_handshakeTimes_2_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_3_valueNext;
  wire       [0:0]    _zz_handshakeTimes_3_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_4_valueNext;
  wire       [0:0]    _zz_handshakeTimes_4_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_5_valueNext;
  wire       [0:0]    _zz_handshakeTimes_5_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_6_valueNext;
  wire       [0:0]    _zz_handshakeTimes_6_valueNext_1;
  wire       [12:0]   _zz_handshakeTimes_7_valueNext;
  wire       [0:0]    _zz_handshakeTimes_7_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_0_valueNext;
  wire       [0:0]    _zz_outSliceNumb_0_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_1_valueNext;
  wire       [0:0]    _zz_outSliceNumb_1_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_2_valueNext;
  wire       [0:0]    _zz_outSliceNumb_2_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_3_valueNext;
  wire       [0:0]    _zz_outSliceNumb_3_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_4_valueNext;
  wire       [0:0]    _zz_outSliceNumb_4_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_5_valueNext;
  wire       [0:0]    _zz_outSliceNumb_5_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_6_valueNext;
  wire       [0:0]    _zz_outSliceNumb_6_valueNext_1;
  wire       [6:0]    _zz_outSliceNumb_7_valueNext;
  wire       [0:0]    _zz_outSliceNumb_7_valueNext_1;
  reg        [6:0]    _zz_when_ArraySlice_l204;
  reg                 _zz_inputStreamArrayData_ready;
  reg        [6:0]    _zz_when_ArraySlice_l208;
  wire       [6:0]    _zz_when_ArraySlice_l208_1;
  wire       [6:0]    _zz_when_ArraySlice_l209;
  wire       [7:0]    _zz_when_ArraySlice_l158;
  wire       [7:0]    _zz_when_ArraySlice_l158_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_3;
  wire       [7:0]    _zz_when_ArraySlice_l159;
  wire       [7:0]    _zz_when_ArraySlice_l159_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_5;
  wire       [7:0]    _zz__zz_realValue_0;
  wire       [7:0]    _zz__zz_realValue_0_1;
  wire       [7:0]    _zz_realValue_0_416;
  wire       [7:0]    _zz_realValue_0_417;
  wire       [7:0]    _zz_realValue_0_418;
  wire       [7:0]    _zz_when_ArraySlice_l166;
  wire       [7:0]    _zz_when_ArraySlice_l166_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l158_1_2;
  wire       [4:0]    _zz_when_ArraySlice_l158_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l158_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l159_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_1_5;
  wire       [7:0]    _zz_when_ArraySlice_l159_1_6;
  wire       [4:0]    _zz_when_ArraySlice_l159_1_7;
  wire       [7:0]    _zz__zz_realValue_0_1_1;
  wire       [7:0]    _zz__zz_realValue_0_1_2;
  wire       [7:0]    _zz_realValue_0_1_1;
  wire       [7:0]    _zz_realValue_0_1_2;
  wire       [7:0]    _zz_realValue_0_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l166_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_6;
  wire       [4:0]    _zz_when_ArraySlice_l166_1_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_1_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l158_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l158_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l158_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l159_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_2_5;
  wire       [7:0]    _zz_when_ArraySlice_l159_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l159_2_7;
  wire       [7:0]    _zz__zz_realValue_0_2;
  wire       [7:0]    _zz__zz_realValue_0_2_1;
  wire       [7:0]    _zz_realValue_0_2_1;
  wire       [7:0]    _zz_realValue_0_2_2;
  wire       [7:0]    _zz_realValue_0_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l166_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_6;
  wire       [5:0]    _zz_when_ArraySlice_l166_2_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_2_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l158_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l158_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l158_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l159_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_3_5;
  wire       [7:0]    _zz_when_ArraySlice_l159_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l159_3_7;
  wire       [7:0]    _zz__zz_realValue_0_3;
  wire       [7:0]    _zz__zz_realValue_0_3_1;
  wire       [7:0]    _zz_realValue_0_3_1;
  wire       [7:0]    _zz_realValue_0_3_2;
  wire       [7:0]    _zz_realValue_0_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l166_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_6;
  wire       [5:0]    _zz_when_ArraySlice_l166_3_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_3_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_4;
  wire       [7:0]    _zz_when_ArraySlice_l158_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l159_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_4_5;
  wire       [7:0]    _zz_when_ArraySlice_l159_4_6;
  wire       [6:0]    _zz_when_ArraySlice_l159_4_7;
  wire       [7:0]    _zz__zz_realValue_0_4;
  wire       [7:0]    _zz__zz_realValue_0_4_1;
  wire       [7:0]    _zz_realValue_0_4_1;
  wire       [7:0]    _zz_realValue_0_4_2;
  wire       [7:0]    _zz_realValue_0_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l166_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_6;
  wire       [6:0]    _zz_when_ArraySlice_l166_4_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_4_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l159_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_5_5;
  wire       [7:0]    _zz_when_ArraySlice_l159_5_6;
  wire       [6:0]    _zz_when_ArraySlice_l159_5_7;
  wire       [7:0]    _zz__zz_realValue_0_5;
  wire       [7:0]    _zz__zz_realValue_0_5_1;
  wire       [7:0]    _zz_realValue_0_5_1;
  wire       [7:0]    _zz_realValue_0_5_2;
  wire       [7:0]    _zz_realValue_0_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_6;
  wire       [6:0]    _zz_when_ArraySlice_l166_5_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_5_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_6;
  wire       [5:0]    _zz_when_ArraySlice_l159_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_6_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_6_6;
  wire       [7:0]    _zz__zz_realValue_0_6;
  wire       [7:0]    _zz__zz_realValue_0_6_1;
  wire       [7:0]    _zz_realValue_0_6_1;
  wire       [7:0]    _zz_realValue_0_6_2;
  wire       [7:0]    _zz_realValue_0_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_1;
  wire       [5:0]    _zz_when_ArraySlice_l166_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_6;
  wire       [6:0]    _zz_when_ArraySlice_l166_6_7;
  wire       [7:0]    _zz_when_ArraySlice_l166_6_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_7;
  wire       [4:0]    _zz_when_ArraySlice_l159_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_7_6;
  wire       [7:0]    _zz__zz_realValue_0_7;
  wire       [7:0]    _zz__zz_realValue_0_7_1;
  wire       [7:0]    _zz_realValue_0_7_1;
  wire       [7:0]    _zz_realValue_0_7_2;
  wire       [7:0]    _zz_realValue_0_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_7;
  wire       [4:0]    _zz_when_ArraySlice_l166_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_7_7;
  wire       [7:0]    _zz_when_ArraySlice_l376;
  wire       [7:0]    _zz_when_ArraySlice_l376_1;
  wire       [3:0]    _zz_when_ArraySlice_l376_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_3;
  reg        [6:0]    _zz_when_ArraySlice_l377;
  wire       [6:0]    _zz_when_ArraySlice_l377_1;
  wire       [7:0]    _zz_when_ArraySlice_l377_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_3;
  wire       [3:0]    _zz_when_ArraySlice_l377_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_0_valid;
  wire       [3:0]    _zz__zz_outputStreamArrayData_0_valid_1;
  wire       [6:0]    _zz__zz_3;
  reg                 _zz_outputStreamArrayData_0_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_0_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_0_payload;
  wire       [6:0]    _zz_outputStreamArrayData_0_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383;
  wire       [6:0]    _zz_when_ArraySlice_l383_1;
  wire       [7:0]    _zz_when_ArraySlice_l383_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_3;
  wire       [3:0]    _zz_when_ArraySlice_l383_4;
  wire       [12:0]   _zz_when_ArraySlice_l384;
  wire       [7:0]    _zz_when_ArraySlice_l384_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_2;
  wire       [7:0]    _zz_selectReadFifo_0;
  wire       [7:0]    _zz_selectReadFifo_0_1;
  wire       [12:0]   _zz_when_ArraySlice_l387;
  wire       [12:0]   _zz_when_ArraySlice_l387_1;
  reg        [6:0]    _zz_when_ArraySlice_l392;
  wire       [6:0]    _zz_when_ArraySlice_l392_1;
  wire       [7:0]    _zz_when_ArraySlice_l392_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_3;
  wire       [3:0]    _zz_when_ArraySlice_l392_4;
  wire       [12:0]   _zz_when_ArraySlice_l393;
  wire       [7:0]    _zz_when_ArraySlice_l393_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_2;
  wire       [7:0]    _zz__zz_realValue1_0;
  wire       [7:0]    _zz__zz_realValue1_0_1;
  wire       [7:0]    _zz_realValue1_0_48;
  wire       [7:0]    _zz_realValue1_0_49;
  wire       [7:0]    _zz_realValue1_0_50;
  wire       [7:0]    _zz_when_ArraySlice_l395;
  wire       [6:0]    _zz_when_ArraySlice_l395_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_2;
  wire       [7:0]    _zz_selectReadFifo_0_2;
  wire       [7:0]    _zz_selectReadFifo_0_3;
  wire       [7:0]    _zz_selectReadFifo_0_4;
  wire       [0:0]    _zz_selectReadFifo_0_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_8;
  wire       [7:0]    _zz_when_ArraySlice_l158_8_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_8_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_8_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_8;
  wire       [7:0]    _zz_when_ArraySlice_l159_8_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_8_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_8_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_8_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_8_5;
  wire       [7:0]    _zz__zz_realValue_0_8;
  wire       [7:0]    _zz__zz_realValue_0_8_1;
  wire       [7:0]    _zz_realValue_0_8_1;
  wire       [7:0]    _zz_realValue_0_8_2;
  wire       [7:0]    _zz_realValue_0_8_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_8;
  wire       [7:0]    _zz_when_ArraySlice_l166_8_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_8_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_8_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_8_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_8_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_8_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_9;
  wire       [7:0]    _zz_when_ArraySlice_l158_9_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_9_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_9_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_9;
  wire       [6:0]    _zz_when_ArraySlice_l159_9_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_9_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_9_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_9_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_9_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_9_6;
  wire       [7:0]    _zz__zz_realValue_0_9;
  wire       [7:0]    _zz__zz_realValue_0_9_1;
  wire       [7:0]    _zz_realValue_0_9_1;
  wire       [7:0]    _zz_realValue_0_9_2;
  wire       [7:0]    _zz_realValue_0_9_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_9;
  wire       [6:0]    _zz_when_ArraySlice_l166_9_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_9_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_9_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_9_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_9_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_9_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_9_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_10_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_10_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_10_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_10;
  wire       [6:0]    _zz_when_ArraySlice_l159_10_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_10_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_10_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_10_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_10_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_10_6;
  wire       [7:0]    _zz__zz_realValue_0_10;
  wire       [7:0]    _zz__zz_realValue_0_10_1;
  wire       [7:0]    _zz_realValue_0_10_1;
  wire       [7:0]    _zz_realValue_0_10_2;
  wire       [7:0]    _zz_realValue_0_10_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_10;
  wire       [6:0]    _zz_when_ArraySlice_l166_10_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_10_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_10_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_10_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_10_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_10_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_10_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_11;
  wire       [7:0]    _zz_when_ArraySlice_l158_11_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_11_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_11_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_11;
  wire       [6:0]    _zz_when_ArraySlice_l159_11_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_11_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_11_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_11_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_11_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_11_6;
  wire       [7:0]    _zz__zz_realValue_0_11;
  wire       [7:0]    _zz__zz_realValue_0_11_1;
  wire       [7:0]    _zz_realValue_0_11_1;
  wire       [7:0]    _zz_realValue_0_11_2;
  wire       [7:0]    _zz_realValue_0_11_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_11;
  wire       [6:0]    _zz_when_ArraySlice_l166_11_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_11_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_11_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_11_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_11_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_11_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_11_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_12;
  wire       [7:0]    _zz_when_ArraySlice_l158_12_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_12_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_12_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_12;
  wire       [6:0]    _zz_when_ArraySlice_l159_12_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_12_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_12_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_12_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_12_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_12_6;
  wire       [7:0]    _zz__zz_realValue_0_12;
  wire       [7:0]    _zz__zz_realValue_0_12_1;
  wire       [7:0]    _zz_realValue_0_12_1;
  wire       [7:0]    _zz_realValue_0_12_2;
  wire       [7:0]    _zz_realValue_0_12_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_12;
  wire       [6:0]    _zz_when_ArraySlice_l166_12_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_12_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_12_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_12_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_12_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_12_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_12_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_13;
  wire       [7:0]    _zz_when_ArraySlice_l158_13_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_13_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_13_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_13;
  wire       [5:0]    _zz_when_ArraySlice_l159_13_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_13_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_13_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_13_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_13_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_13_6;
  wire       [7:0]    _zz__zz_realValue_0_13;
  wire       [7:0]    _zz__zz_realValue_0_13_1;
  wire       [7:0]    _zz_realValue_0_13_1;
  wire       [7:0]    _zz_realValue_0_13_2;
  wire       [7:0]    _zz_realValue_0_13_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_13;
  wire       [5:0]    _zz_when_ArraySlice_l166_13_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_13_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_13_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_13_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_13_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_13_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_13_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_14;
  wire       [7:0]    _zz_when_ArraySlice_l158_14_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_14_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_14_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_14;
  wire       [5:0]    _zz_when_ArraySlice_l159_14_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_14_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_14_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_14_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_14_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_14_6;
  wire       [7:0]    _zz__zz_realValue_0_14;
  wire       [7:0]    _zz__zz_realValue_0_14_1;
  wire       [7:0]    _zz_realValue_0_14_1;
  wire       [7:0]    _zz_realValue_0_14_2;
  wire       [7:0]    _zz_realValue_0_14_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_14;
  wire       [5:0]    _zz_when_ArraySlice_l166_14_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_14_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_14_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_14_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_14_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_14_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_14_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_15_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_15_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_15_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_15;
  wire       [4:0]    _zz_when_ArraySlice_l159_15_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_15_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_15_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_15_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_15_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_15_6;
  wire       [7:0]    _zz__zz_realValue_0_15;
  wire       [7:0]    _zz__zz_realValue_0_15_1;
  wire       [7:0]    _zz_realValue_0_15_1;
  wire       [7:0]    _zz_realValue_0_15_2;
  wire       [7:0]    _zz_realValue_0_15_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_15;
  wire       [4:0]    _zz_when_ArraySlice_l166_15_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_15_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_15_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_15_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_15_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_15_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_15_7;
  wire                _zz_when_ArraySlice_l400;
  wire                _zz_when_ArraySlice_l400_1;
  wire                _zz_when_ArraySlice_l400_2;
  wire                _zz_when_ArraySlice_l400_3;
  wire                _zz_when_ArraySlice_l400_4;
  wire                _zz_when_ArraySlice_l400_5;
  wire                _zz_when_ArraySlice_l400_6;
  wire                _zz_when_ArraySlice_l400_7;
  wire                _zz_when_ArraySlice_l400_8;
  wire                _zz_when_ArraySlice_l400_9;
  wire       [7:0]    _zz_when_ArraySlice_l403;
  wire       [7:0]    _zz_when_ArraySlice_l403_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_4;
  wire       [6:0]    _zz_when_ArraySlice_l403_5;
  wire       [7:0]    _zz_when_ArraySlice_l403_6;
  wire       [3:0]    _zz_when_ArraySlice_l403_7;
  wire       [7:0]    _zz_when_ArraySlice_l406;
  wire       [7:0]    _zz_when_ArraySlice_l406_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_3;
  wire       [6:0]    _zz_when_ArraySlice_l406_4;
  wire       [7:0]    _zz_selectReadFifo_0_6;
  wire       [7:0]    _zz_selectReadFifo_0_7;
  wire       [6:0]    _zz_selectReadFifo_0_8;
  wire       [12:0]   _zz_when_ArraySlice_l413;
  wire       [12:0]   _zz_when_ArraySlice_l413_1;
  reg        [6:0]    _zz_when_ArraySlice_l417;
  wire       [6:0]    _zz_when_ArraySlice_l417_1;
  wire       [7:0]    _zz_when_ArraySlice_l417_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_3;
  wire       [3:0]    _zz_when_ArraySlice_l417_4;
  wire       [12:0]   _zz_when_ArraySlice_l418;
  wire       [7:0]    _zz_when_ArraySlice_l418_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_3;
  wire       [0:0]    _zz_when_ArraySlice_l418_4;
  wire       [7:0]    _zz__zz_realValue1_0_1_1;
  wire       [7:0]    _zz__zz_realValue1_0_1_2;
  wire       [7:0]    _zz_realValue1_0_1_1;
  wire       [7:0]    _zz_realValue1_0_1_2;
  wire       [7:0]    _zz_realValue1_0_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l420;
  wire       [6:0]    _zz_when_ArraySlice_l420_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_2;
  wire       [7:0]    _zz_selectReadFifo_0_9;
  wire       [7:0]    _zz_selectReadFifo_0_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_16;
  wire       [7:0]    _zz_when_ArraySlice_l158_16_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_16_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_16_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_16;
  wire       [7:0]    _zz_when_ArraySlice_l159_16_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_16_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_16_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_16_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_16_5;
  wire       [7:0]    _zz__zz_realValue_0_16;
  wire       [7:0]    _zz__zz_realValue_0_16_1;
  wire       [7:0]    _zz_realValue_0_16_1;
  wire       [7:0]    _zz_realValue_0_16_2;
  wire       [7:0]    _zz_realValue_0_16_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_16;
  wire       [7:0]    _zz_when_ArraySlice_l166_16_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_16_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_16_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_16_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_16_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_16_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_17;
  wire       [7:0]    _zz_when_ArraySlice_l158_17_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_17_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_17_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_17;
  wire       [6:0]    _zz_when_ArraySlice_l159_17_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_17_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_17_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_17_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_17_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_17_6;
  wire       [7:0]    _zz__zz_realValue_0_17;
  wire       [7:0]    _zz__zz_realValue_0_17_1;
  wire       [7:0]    _zz_realValue_0_17_1;
  wire       [7:0]    _zz_realValue_0_17_2;
  wire       [7:0]    _zz_realValue_0_17_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_17;
  wire       [6:0]    _zz_when_ArraySlice_l166_17_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_17_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_17_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_17_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_17_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_17_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_17_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_18;
  wire       [7:0]    _zz_when_ArraySlice_l158_18_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_18_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_18_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_18;
  wire       [6:0]    _zz_when_ArraySlice_l159_18_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_18_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_18_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_18_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_18_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_18_6;
  wire       [7:0]    _zz__zz_realValue_0_18;
  wire       [7:0]    _zz__zz_realValue_0_18_1;
  wire       [7:0]    _zz_realValue_0_18_1;
  wire       [7:0]    _zz_realValue_0_18_2;
  wire       [7:0]    _zz_realValue_0_18_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_18;
  wire       [6:0]    _zz_when_ArraySlice_l166_18_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_18_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_18_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_18_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_18_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_18_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_18_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_19;
  wire       [7:0]    _zz_when_ArraySlice_l158_19_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_19_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_19_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_19;
  wire       [6:0]    _zz_when_ArraySlice_l159_19_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_19_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_19_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_19_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_19_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_19_6;
  wire       [7:0]    _zz__zz_realValue_0_19;
  wire       [7:0]    _zz__zz_realValue_0_19_1;
  wire       [7:0]    _zz_realValue_0_19_1;
  wire       [7:0]    _zz_realValue_0_19_2;
  wire       [7:0]    _zz_realValue_0_19_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_19;
  wire       [6:0]    _zz_when_ArraySlice_l166_19_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_19_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_19_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_19_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_19_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_19_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_19_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_20;
  wire       [7:0]    _zz_when_ArraySlice_l158_20_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_20_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_20_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_20;
  wire       [6:0]    _zz_when_ArraySlice_l159_20_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_20_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_20_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_20_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_20_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_20_6;
  wire       [7:0]    _zz__zz_realValue_0_20;
  wire       [7:0]    _zz__zz_realValue_0_20_1;
  wire       [7:0]    _zz_realValue_0_20_1;
  wire       [7:0]    _zz_realValue_0_20_2;
  wire       [7:0]    _zz_realValue_0_20_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_20;
  wire       [6:0]    _zz_when_ArraySlice_l166_20_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_20_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_20_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_20_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_20_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_20_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_20_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_21_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_21_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_21_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_21;
  wire       [5:0]    _zz_when_ArraySlice_l159_21_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_21_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_21_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_21_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_21_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_21_6;
  wire       [7:0]    _zz__zz_realValue_0_21;
  wire       [7:0]    _zz__zz_realValue_0_21_1;
  wire       [7:0]    _zz_realValue_0_21_1;
  wire       [7:0]    _zz_realValue_0_21_2;
  wire       [7:0]    _zz_realValue_0_21_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_21;
  wire       [5:0]    _zz_when_ArraySlice_l166_21_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_21_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_21_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_21_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_21_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_21_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_21_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_22;
  wire       [7:0]    _zz_when_ArraySlice_l158_22_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_22_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_22_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_22;
  wire       [5:0]    _zz_when_ArraySlice_l159_22_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_22_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_22_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_22_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_22_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_22_6;
  wire       [7:0]    _zz__zz_realValue_0_22;
  wire       [7:0]    _zz__zz_realValue_0_22_1;
  wire       [7:0]    _zz_realValue_0_22_1;
  wire       [7:0]    _zz_realValue_0_22_2;
  wire       [7:0]    _zz_realValue_0_22_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_22;
  wire       [5:0]    _zz_when_ArraySlice_l166_22_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_22_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_22_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_22_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_22_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_22_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_22_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_23;
  wire       [7:0]    _zz_when_ArraySlice_l158_23_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_23_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_23_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_23;
  wire       [4:0]    _zz_when_ArraySlice_l159_23_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_23_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_23_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_23_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_23_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_23_6;
  wire       [7:0]    _zz__zz_realValue_0_23;
  wire       [7:0]    _zz__zz_realValue_0_23_1;
  wire       [7:0]    _zz_realValue_0_23_1;
  wire       [7:0]    _zz_realValue_0_23_2;
  wire       [7:0]    _zz_realValue_0_23_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_23;
  wire       [4:0]    _zz_when_ArraySlice_l166_23_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_23_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_23_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_23_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_23_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_23_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_23_7;
  wire                _zz_when_ArraySlice_l425;
  wire                _zz_when_ArraySlice_l425_1;
  wire                _zz_when_ArraySlice_l425_2;
  wire                _zz_when_ArraySlice_l425_3;
  wire                _zz_when_ArraySlice_l425_4;
  wire                _zz_when_ArraySlice_l425_5;
  wire       [7:0]    _zz_when_ArraySlice_l428;
  wire       [7:0]    _zz_when_ArraySlice_l428_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_4;
  wire       [6:0]    _zz_when_ArraySlice_l428_5;
  wire       [7:0]    _zz_when_ArraySlice_l428_6;
  wire       [3:0]    _zz_when_ArraySlice_l428_7;
  wire       [7:0]    _zz_when_ArraySlice_l431;
  wire       [7:0]    _zz_when_ArraySlice_l431_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_3;
  wire       [6:0]    _zz_when_ArraySlice_l431_4;
  wire       [7:0]    _zz_selectReadFifo_0_11;
  wire       [7:0]    _zz_selectReadFifo_0_12;
  wire       [6:0]    _zz_selectReadFifo_0_13;
  wire       [12:0]   _zz_when_ArraySlice_l438;
  wire       [12:0]   _zz_when_ArraySlice_l438_1;
  wire       [12:0]   _zz_when_ArraySlice_l449;
  wire       [7:0]    _zz_when_ArraySlice_l449_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_2;
  wire       [7:0]    _zz__zz_realValue1_0_2;
  wire       [7:0]    _zz__zz_realValue1_0_2_1;
  wire       [7:0]    _zz_realValue1_0_2_1;
  wire       [7:0]    _zz_realValue1_0_2_2;
  wire       [7:0]    _zz_realValue1_0_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l450;
  wire       [6:0]    _zz_when_ArraySlice_l450_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_2;
  wire       [7:0]    _zz_selectReadFifo_0_14;
  wire       [7:0]    _zz_selectReadFifo_0_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_24;
  wire       [7:0]    _zz_when_ArraySlice_l158_24_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_24_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_24_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_24;
  wire       [7:0]    _zz_when_ArraySlice_l159_24_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_24_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_24_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_24_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_24_5;
  wire       [7:0]    _zz__zz_realValue_0_24;
  wire       [7:0]    _zz__zz_realValue_0_24_1;
  wire       [7:0]    _zz_realValue_0_24_1;
  wire       [7:0]    _zz_realValue_0_24_2;
  wire       [7:0]    _zz_realValue_0_24_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_24;
  wire       [7:0]    _zz_when_ArraySlice_l166_24_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_24_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_24_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_24_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_24_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_24_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_25;
  wire       [7:0]    _zz_when_ArraySlice_l158_25_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_25_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_25_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_25;
  wire       [6:0]    _zz_when_ArraySlice_l159_25_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_25_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_25_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_25_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_25_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_25_6;
  wire       [7:0]    _zz__zz_realValue_0_25;
  wire       [7:0]    _zz__zz_realValue_0_25_1;
  wire       [7:0]    _zz_realValue_0_25_1;
  wire       [7:0]    _zz_realValue_0_25_2;
  wire       [7:0]    _zz_realValue_0_25_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_25;
  wire       [6:0]    _zz_when_ArraySlice_l166_25_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_25_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_25_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_25_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_25_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_25_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_25_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_26_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_26_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_26_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_26;
  wire       [6:0]    _zz_when_ArraySlice_l159_26_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_26_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_26_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_26_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_26_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_26_6;
  wire       [7:0]    _zz__zz_realValue_0_26;
  wire       [7:0]    _zz__zz_realValue_0_26_1;
  wire       [7:0]    _zz_realValue_0_26_1;
  wire       [7:0]    _zz_realValue_0_26_2;
  wire       [7:0]    _zz_realValue_0_26_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_26;
  wire       [6:0]    _zz_when_ArraySlice_l166_26_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_26_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_26_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_26_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_26_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_26_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_26_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_27;
  wire       [7:0]    _zz_when_ArraySlice_l158_27_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_27_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_27_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_27;
  wire       [6:0]    _zz_when_ArraySlice_l159_27_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_27_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_27_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_27_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_27_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_27_6;
  wire       [7:0]    _zz__zz_realValue_0_27;
  wire       [7:0]    _zz__zz_realValue_0_27_1;
  wire       [7:0]    _zz_realValue_0_27_1;
  wire       [7:0]    _zz_realValue_0_27_2;
  wire       [7:0]    _zz_realValue_0_27_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_27;
  wire       [6:0]    _zz_when_ArraySlice_l166_27_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_27_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_27_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_27_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_27_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_27_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_27_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_28;
  wire       [7:0]    _zz_when_ArraySlice_l158_28_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_28_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_28_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_28;
  wire       [6:0]    _zz_when_ArraySlice_l159_28_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_28_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_28_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_28_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_28_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_28_6;
  wire       [7:0]    _zz__zz_realValue_0_28;
  wire       [7:0]    _zz__zz_realValue_0_28_1;
  wire       [7:0]    _zz_realValue_0_28_1;
  wire       [7:0]    _zz_realValue_0_28_2;
  wire       [7:0]    _zz_realValue_0_28_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_28;
  wire       [6:0]    _zz_when_ArraySlice_l166_28_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_28_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_28_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_28_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_28_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_28_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_28_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_29;
  wire       [7:0]    _zz_when_ArraySlice_l158_29_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_29_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_29_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_29;
  wire       [5:0]    _zz_when_ArraySlice_l159_29_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_29_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_29_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_29_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_29_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_29_6;
  wire       [7:0]    _zz__zz_realValue_0_29;
  wire       [7:0]    _zz__zz_realValue_0_29_1;
  wire       [7:0]    _zz_realValue_0_29_1;
  wire       [7:0]    _zz_realValue_0_29_2;
  wire       [7:0]    _zz_realValue_0_29_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_29;
  wire       [5:0]    _zz_when_ArraySlice_l166_29_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_29_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_29_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_29_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_29_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_29_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_29_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_30;
  wire       [7:0]    _zz_when_ArraySlice_l158_30_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_30_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_30_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_30;
  wire       [5:0]    _zz_when_ArraySlice_l159_30_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_30_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_30_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_30_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_30_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_30_6;
  wire       [7:0]    _zz__zz_realValue_0_30;
  wire       [7:0]    _zz__zz_realValue_0_30_1;
  wire       [7:0]    _zz_realValue_0_30_1;
  wire       [7:0]    _zz_realValue_0_30_2;
  wire       [7:0]    _zz_realValue_0_30_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_30;
  wire       [5:0]    _zz_when_ArraySlice_l166_30_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_30_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_30_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_30_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_30_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_30_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_30_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_31_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_31_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_31_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_31;
  wire       [4:0]    _zz_when_ArraySlice_l159_31_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_31_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_31_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_31_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_31_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_31_6;
  wire       [7:0]    _zz__zz_realValue_0_31;
  wire       [7:0]    _zz__zz_realValue_0_31_1;
  wire       [7:0]    _zz_realValue_0_31_1;
  wire       [7:0]    _zz_realValue_0_31_2;
  wire       [7:0]    _zz_realValue_0_31_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_31;
  wire       [4:0]    _zz_when_ArraySlice_l166_31_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_31_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_31_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_31_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_31_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_31_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_31_7;
  wire                _zz_when_ArraySlice_l457;
  wire                _zz_when_ArraySlice_l457_1;
  wire                _zz_when_ArraySlice_l457_2;
  wire                _zz_when_ArraySlice_l457_3;
  wire                _zz_when_ArraySlice_l457_4;
  wire                _zz_when_ArraySlice_l457_5;
  wire       [12:0]   _zz_when_ArraySlice_l461;
  wire       [12:0]   _zz_when_ArraySlice_l461_1;
  wire       [7:0]    _zz_when_ArraySlice_l447;
  wire       [7:0]    _zz_when_ArraySlice_l447_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_2;
  wire       [3:0]    _zz_when_ArraySlice_l447_3;
  wire       [12:0]   _zz_when_ArraySlice_l468;
  wire       [7:0]    _zz_when_ArraySlice_l468_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l376_1_2;
  wire       [4:0]    _zz_when_ArraySlice_l376_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l376_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l377_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l377_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l377_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l377_1_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_1_valid;
  wire       [4:0]    _zz__zz_outputStreamArrayData_1_valid_1;
  wire       [6:0]    _zz__zz_4;
  reg                 _zz_outputStreamArrayData_1_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_1_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_1_payload;
  wire       [6:0]    _zz_outputStreamArrayData_1_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l383_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l383_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l383_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l384_1_3;
  wire       [7:0]    _zz_selectReadFifo_1;
  wire       [7:0]    _zz_selectReadFifo_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l392_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l392_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l392_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l393_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l393_1_3;
  wire       [7:0]    _zz__zz_realValue1_0_3;
  wire       [7:0]    _zz__zz_realValue1_0_3_1;
  wire       [7:0]    _zz_realValue1_0_3_1;
  wire       [7:0]    _zz_realValue1_0_3_2;
  wire       [7:0]    _zz_realValue1_0_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l395_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l395_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_2;
  wire       [7:0]    _zz_selectReadFifo_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_4;
  wire       [0:0]    _zz_selectReadFifo_1_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_32;
  wire       [7:0]    _zz_when_ArraySlice_l158_32_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_32_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_32_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_32;
  wire       [7:0]    _zz_when_ArraySlice_l159_32_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_32_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_32_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_32_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_32_5;
  wire       [7:0]    _zz__zz_realValue_0_32;
  wire       [7:0]    _zz__zz_realValue_0_32_1;
  wire       [7:0]    _zz_realValue_0_32_1;
  wire       [7:0]    _zz_realValue_0_32_2;
  wire       [7:0]    _zz_realValue_0_32_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_32;
  wire       [7:0]    _zz_when_ArraySlice_l166_32_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_32_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_32_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_32_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_32_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_32_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_33;
  wire       [7:0]    _zz_when_ArraySlice_l158_33_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_33_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_33_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_33;
  wire       [6:0]    _zz_when_ArraySlice_l159_33_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_33_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_33_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_33_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_33_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_33_6;
  wire       [7:0]    _zz__zz_realValue_0_33;
  wire       [7:0]    _zz__zz_realValue_0_33_1;
  wire       [7:0]    _zz_realValue_0_33_1;
  wire       [7:0]    _zz_realValue_0_33_2;
  wire       [7:0]    _zz_realValue_0_33_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_33;
  wire       [6:0]    _zz_when_ArraySlice_l166_33_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_33_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_33_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_33_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_33_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_33_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_33_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_34;
  wire       [7:0]    _zz_when_ArraySlice_l158_34_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_34_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_34_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_34;
  wire       [6:0]    _zz_when_ArraySlice_l159_34_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_34_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_34_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_34_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_34_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_34_6;
  wire       [7:0]    _zz__zz_realValue_0_34;
  wire       [7:0]    _zz__zz_realValue_0_34_1;
  wire       [7:0]    _zz_realValue_0_34_1;
  wire       [7:0]    _zz_realValue_0_34_2;
  wire       [7:0]    _zz_realValue_0_34_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_34;
  wire       [6:0]    _zz_when_ArraySlice_l166_34_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_34_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_34_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_34_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_34_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_34_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_34_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_35;
  wire       [7:0]    _zz_when_ArraySlice_l158_35_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_35_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_35_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_35;
  wire       [6:0]    _zz_when_ArraySlice_l159_35_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_35_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_35_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_35_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_35_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_35_6;
  wire       [7:0]    _zz__zz_realValue_0_35;
  wire       [7:0]    _zz__zz_realValue_0_35_1;
  wire       [7:0]    _zz_realValue_0_35_1;
  wire       [7:0]    _zz_realValue_0_35_2;
  wire       [7:0]    _zz_realValue_0_35_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_35;
  wire       [6:0]    _zz_when_ArraySlice_l166_35_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_35_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_35_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_35_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_35_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_35_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_35_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_36;
  wire       [7:0]    _zz_when_ArraySlice_l158_36_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_36_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_36_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_36;
  wire       [6:0]    _zz_when_ArraySlice_l159_36_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_36_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_36_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_36_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_36_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_36_6;
  wire       [7:0]    _zz__zz_realValue_0_36;
  wire       [7:0]    _zz__zz_realValue_0_36_1;
  wire       [7:0]    _zz_realValue_0_36_1;
  wire       [7:0]    _zz_realValue_0_36_2;
  wire       [7:0]    _zz_realValue_0_36_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_36;
  wire       [6:0]    _zz_when_ArraySlice_l166_36_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_36_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_36_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_36_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_36_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_36_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_36_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_37;
  wire       [7:0]    _zz_when_ArraySlice_l158_37_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_37_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_37_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_37;
  wire       [5:0]    _zz_when_ArraySlice_l159_37_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_37_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_37_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_37_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_37_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_37_6;
  wire       [7:0]    _zz__zz_realValue_0_37;
  wire       [7:0]    _zz__zz_realValue_0_37_1;
  wire       [7:0]    _zz_realValue_0_37_1;
  wire       [7:0]    _zz_realValue_0_37_2;
  wire       [7:0]    _zz_realValue_0_37_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_37;
  wire       [5:0]    _zz_when_ArraySlice_l166_37_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_37_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_37_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_37_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_37_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_37_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_37_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_38;
  wire       [7:0]    _zz_when_ArraySlice_l158_38_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_38_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_38_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_38;
  wire       [5:0]    _zz_when_ArraySlice_l159_38_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_38_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_38_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_38_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_38_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_38_6;
  wire       [7:0]    _zz__zz_realValue_0_38;
  wire       [7:0]    _zz__zz_realValue_0_38_1;
  wire       [7:0]    _zz_realValue_0_38_1;
  wire       [7:0]    _zz_realValue_0_38_2;
  wire       [7:0]    _zz_realValue_0_38_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_38;
  wire       [5:0]    _zz_when_ArraySlice_l166_38_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_38_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_38_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_38_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_38_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_38_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_38_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_39;
  wire       [7:0]    _zz_when_ArraySlice_l158_39_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_39_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_39_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_39;
  wire       [4:0]    _zz_when_ArraySlice_l159_39_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_39_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_39_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_39_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_39_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_39_6;
  wire       [7:0]    _zz__zz_realValue_0_39;
  wire       [7:0]    _zz__zz_realValue_0_39_1;
  wire       [7:0]    _zz_realValue_0_39_1;
  wire       [7:0]    _zz_realValue_0_39_2;
  wire       [7:0]    _zz_realValue_0_39_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_39;
  wire       [4:0]    _zz_when_ArraySlice_l166_39_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_39_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_39_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_39_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_39_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_39_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_39_7;
  wire                _zz_when_ArraySlice_l400_1_1;
  wire                _zz_when_ArraySlice_l400_1_2;
  wire                _zz_when_ArraySlice_l400_1_3;
  wire                _zz_when_ArraySlice_l400_1_4;
  wire                _zz_when_ArraySlice_l400_1_5;
  wire                _zz_when_ArraySlice_l400_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_1_7;
  wire       [4:0]    _zz_when_ArraySlice_l403_1_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l406_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l406_1_5;
  wire       [7:0]    _zz_selectReadFifo_1_6;
  wire       [7:0]    _zz_selectReadFifo_1_7;
  wire       [6:0]    _zz_selectReadFifo_1_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l413_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l417_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l417_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l417_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l417_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l418_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l418_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l418_1_5;
  wire       [7:0]    _zz__zz_realValue1_0_4;
  wire       [7:0]    _zz__zz_realValue1_0_4_1;
  wire       [7:0]    _zz_realValue1_0_4_1;
  wire       [7:0]    _zz_realValue1_0_4_2;
  wire       [7:0]    _zz_realValue1_0_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l420_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l420_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_9;
  wire       [7:0]    _zz_selectReadFifo_1_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_40;
  wire       [7:0]    _zz_when_ArraySlice_l158_40_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_40_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_40_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_40;
  wire       [7:0]    _zz_when_ArraySlice_l159_40_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_40_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_40_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_40_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_40_5;
  wire       [7:0]    _zz__zz_realValue_0_40;
  wire       [7:0]    _zz__zz_realValue_0_40_1;
  wire       [7:0]    _zz_realValue_0_40_1;
  wire       [7:0]    _zz_realValue_0_40_2;
  wire       [7:0]    _zz_realValue_0_40_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_40;
  wire       [7:0]    _zz_when_ArraySlice_l166_40_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_40_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_40_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_40_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_40_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_40_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_41;
  wire       [7:0]    _zz_when_ArraySlice_l158_41_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_41_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_41_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_41;
  wire       [6:0]    _zz_when_ArraySlice_l159_41_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_41_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_41_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_41_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_41_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_41_6;
  wire       [7:0]    _zz__zz_realValue_0_41;
  wire       [7:0]    _zz__zz_realValue_0_41_1;
  wire       [7:0]    _zz_realValue_0_41_1;
  wire       [7:0]    _zz_realValue_0_41_2;
  wire       [7:0]    _zz_realValue_0_41_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_41;
  wire       [6:0]    _zz_when_ArraySlice_l166_41_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_41_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_41_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_41_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_41_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_41_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_41_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_42;
  wire       [7:0]    _zz_when_ArraySlice_l158_42_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_42_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_42_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_42;
  wire       [6:0]    _zz_when_ArraySlice_l159_42_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_42_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_42_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_42_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_42_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_42_6;
  wire       [7:0]    _zz__zz_realValue_0_42;
  wire       [7:0]    _zz__zz_realValue_0_42_1;
  wire       [7:0]    _zz_realValue_0_42_1;
  wire       [7:0]    _zz_realValue_0_42_2;
  wire       [7:0]    _zz_realValue_0_42_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_42;
  wire       [6:0]    _zz_when_ArraySlice_l166_42_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_42_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_42_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_42_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_42_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_42_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_42_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_43;
  wire       [7:0]    _zz_when_ArraySlice_l158_43_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_43_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_43_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_43;
  wire       [6:0]    _zz_when_ArraySlice_l159_43_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_43_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_43_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_43_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_43_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_43_6;
  wire       [7:0]    _zz__zz_realValue_0_43;
  wire       [7:0]    _zz__zz_realValue_0_43_1;
  wire       [7:0]    _zz_realValue_0_43_1;
  wire       [7:0]    _zz_realValue_0_43_2;
  wire       [7:0]    _zz_realValue_0_43_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_43;
  wire       [6:0]    _zz_when_ArraySlice_l166_43_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_43_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_43_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_43_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_43_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_43_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_43_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_44;
  wire       [7:0]    _zz_when_ArraySlice_l158_44_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_44_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_44_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_44;
  wire       [6:0]    _zz_when_ArraySlice_l159_44_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_44_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_44_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_44_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_44_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_44_6;
  wire       [7:0]    _zz__zz_realValue_0_44;
  wire       [7:0]    _zz__zz_realValue_0_44_1;
  wire       [7:0]    _zz_realValue_0_44_1;
  wire       [7:0]    _zz_realValue_0_44_2;
  wire       [7:0]    _zz_realValue_0_44_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_44;
  wire       [6:0]    _zz_when_ArraySlice_l166_44_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_44_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_44_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_44_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_44_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_44_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_44_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_45;
  wire       [7:0]    _zz_when_ArraySlice_l158_45_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_45_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_45_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_45;
  wire       [5:0]    _zz_when_ArraySlice_l159_45_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_45_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_45_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_45_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_45_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_45_6;
  wire       [7:0]    _zz__zz_realValue_0_45;
  wire       [7:0]    _zz__zz_realValue_0_45_1;
  wire       [7:0]    _zz_realValue_0_45_1;
  wire       [7:0]    _zz_realValue_0_45_2;
  wire       [7:0]    _zz_realValue_0_45_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_45;
  wire       [5:0]    _zz_when_ArraySlice_l166_45_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_45_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_45_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_45_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_45_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_45_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_45_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_46;
  wire       [7:0]    _zz_when_ArraySlice_l158_46_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_46_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_46_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_46;
  wire       [5:0]    _zz_when_ArraySlice_l159_46_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_46_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_46_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_46_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_46_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_46_6;
  wire       [7:0]    _zz__zz_realValue_0_46;
  wire       [7:0]    _zz__zz_realValue_0_46_1;
  wire       [7:0]    _zz_realValue_0_46_1;
  wire       [7:0]    _zz_realValue_0_46_2;
  wire       [7:0]    _zz_realValue_0_46_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_46;
  wire       [5:0]    _zz_when_ArraySlice_l166_46_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_46_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_46_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_46_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_46_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_46_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_46_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_47;
  wire       [7:0]    _zz_when_ArraySlice_l158_47_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_47_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_47_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_47;
  wire       [4:0]    _zz_when_ArraySlice_l159_47_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_47_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_47_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_47_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_47_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_47_6;
  wire       [7:0]    _zz__zz_realValue_0_47;
  wire       [7:0]    _zz__zz_realValue_0_47_1;
  wire       [7:0]    _zz_realValue_0_47_1;
  wire       [7:0]    _zz_realValue_0_47_2;
  wire       [7:0]    _zz_realValue_0_47_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_47;
  wire       [4:0]    _zz_when_ArraySlice_l166_47_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_47_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_47_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_47_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_47_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_47_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_47_7;
  wire                _zz_when_ArraySlice_l425_1_1;
  wire                _zz_when_ArraySlice_l425_1_2;
  wire                _zz_when_ArraySlice_l425_1_3;
  wire                _zz_when_ArraySlice_l425_1_4;
  wire                _zz_when_ArraySlice_l425_1_5;
  wire                _zz_when_ArraySlice_l425_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_1_7;
  wire       [4:0]    _zz_when_ArraySlice_l428_1_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l431_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l431_1_5;
  wire       [7:0]    _zz_selectReadFifo_1_11;
  wire       [7:0]    _zz_selectReadFifo_1_12;
  wire       [6:0]    _zz_selectReadFifo_1_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l438_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l449_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l449_1_3;
  wire       [7:0]    _zz__zz_realValue1_0_5;
  wire       [7:0]    _zz__zz_realValue1_0_5_1;
  wire       [7:0]    _zz_realValue1_0_5_1;
  wire       [7:0]    _zz_realValue1_0_5_2;
  wire       [7:0]    _zz_realValue1_0_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l450_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l450_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_14;
  wire       [7:0]    _zz_selectReadFifo_1_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_48;
  wire       [7:0]    _zz_when_ArraySlice_l158_48_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_48_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_48_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_48;
  wire       [7:0]    _zz_when_ArraySlice_l159_48_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_48_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_48_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_48_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_48_5;
  wire       [7:0]    _zz__zz_realValue_0_48;
  wire       [7:0]    _zz__zz_realValue_0_48_1;
  wire       [7:0]    _zz_realValue_0_48_1;
  wire       [7:0]    _zz_realValue_0_48_2;
  wire       [7:0]    _zz_realValue_0_48_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_48;
  wire       [7:0]    _zz_when_ArraySlice_l166_48_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_48_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_48_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_48_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_48_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_48_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_49;
  wire       [7:0]    _zz_when_ArraySlice_l158_49_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_49_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_49_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_49;
  wire       [6:0]    _zz_when_ArraySlice_l159_49_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_49_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_49_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_49_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_49_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_49_6;
  wire       [7:0]    _zz__zz_realValue_0_49;
  wire       [7:0]    _zz__zz_realValue_0_49_1;
  wire       [7:0]    _zz_realValue_0_49_1;
  wire       [7:0]    _zz_realValue_0_49_2;
  wire       [7:0]    _zz_realValue_0_49_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_49;
  wire       [6:0]    _zz_when_ArraySlice_l166_49_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_49_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_49_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_49_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_49_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_49_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_49_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_50;
  wire       [7:0]    _zz_when_ArraySlice_l158_50_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_50_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_50_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_50;
  wire       [6:0]    _zz_when_ArraySlice_l159_50_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_50_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_50_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_50_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_50_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_50_6;
  wire       [7:0]    _zz__zz_realValue_0_50;
  wire       [7:0]    _zz__zz_realValue_0_50_1;
  wire       [7:0]    _zz_realValue_0_50_1;
  wire       [7:0]    _zz_realValue_0_50_2;
  wire       [7:0]    _zz_realValue_0_50_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_50;
  wire       [6:0]    _zz_when_ArraySlice_l166_50_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_50_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_50_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_50_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_50_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_50_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_50_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_51;
  wire       [7:0]    _zz_when_ArraySlice_l158_51_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_51_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_51_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_51;
  wire       [6:0]    _zz_when_ArraySlice_l159_51_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_51_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_51_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_51_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_51_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_51_6;
  wire       [7:0]    _zz__zz_realValue_0_51;
  wire       [7:0]    _zz__zz_realValue_0_51_1;
  wire       [7:0]    _zz_realValue_0_51_1;
  wire       [7:0]    _zz_realValue_0_51_2;
  wire       [7:0]    _zz_realValue_0_51_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_51;
  wire       [6:0]    _zz_when_ArraySlice_l166_51_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_51_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_51_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_51_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_51_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_51_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_51_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_52;
  wire       [7:0]    _zz_when_ArraySlice_l158_52_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_52_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_52_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_52;
  wire       [6:0]    _zz_when_ArraySlice_l159_52_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_52_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_52_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_52_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_52_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_52_6;
  wire       [7:0]    _zz__zz_realValue_0_52;
  wire       [7:0]    _zz__zz_realValue_0_52_1;
  wire       [7:0]    _zz_realValue_0_52_1;
  wire       [7:0]    _zz_realValue_0_52_2;
  wire       [7:0]    _zz_realValue_0_52_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_52;
  wire       [6:0]    _zz_when_ArraySlice_l166_52_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_52_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_52_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_52_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_52_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_52_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_52_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_53;
  wire       [7:0]    _zz_when_ArraySlice_l158_53_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_53_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_53_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_53;
  wire       [5:0]    _zz_when_ArraySlice_l159_53_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_53_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_53_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_53_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_53_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_53_6;
  wire       [7:0]    _zz__zz_realValue_0_53;
  wire       [7:0]    _zz__zz_realValue_0_53_1;
  wire       [7:0]    _zz_realValue_0_53_1;
  wire       [7:0]    _zz_realValue_0_53_2;
  wire       [7:0]    _zz_realValue_0_53_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_53;
  wire       [5:0]    _zz_when_ArraySlice_l166_53_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_53_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_53_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_53_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_53_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_53_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_53_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_54;
  wire       [7:0]    _zz_when_ArraySlice_l158_54_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_54_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_54_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_54;
  wire       [5:0]    _zz_when_ArraySlice_l159_54_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_54_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_54_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_54_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_54_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_54_6;
  wire       [7:0]    _zz__zz_realValue_0_54;
  wire       [7:0]    _zz__zz_realValue_0_54_1;
  wire       [7:0]    _zz_realValue_0_54_1;
  wire       [7:0]    _zz_realValue_0_54_2;
  wire       [7:0]    _zz_realValue_0_54_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_54;
  wire       [5:0]    _zz_when_ArraySlice_l166_54_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_54_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_54_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_54_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_54_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_54_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_54_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_55;
  wire       [7:0]    _zz_when_ArraySlice_l158_55_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_55_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_55_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_55;
  wire       [4:0]    _zz_when_ArraySlice_l159_55_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_55_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_55_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_55_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_55_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_55_6;
  wire       [7:0]    _zz__zz_realValue_0_55;
  wire       [7:0]    _zz__zz_realValue_0_55_1;
  wire       [7:0]    _zz_realValue_0_55_1;
  wire       [7:0]    _zz_realValue_0_55_2;
  wire       [7:0]    _zz_realValue_0_55_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_55;
  wire       [4:0]    _zz_when_ArraySlice_l166_55_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_55_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_55_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_55_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_55_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_55_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_55_7;
  wire                _zz_when_ArraySlice_l457_1_1;
  wire                _zz_when_ArraySlice_l457_1_2;
  wire                _zz_when_ArraySlice_l457_1_3;
  wire                _zz_when_ArraySlice_l457_1_4;
  wire                _zz_when_ArraySlice_l457_1_5;
  wire                _zz_when_ArraySlice_l457_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l461_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l447_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l447_1_3;
  wire       [4:0]    _zz_when_ArraySlice_l447_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l468_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l468_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l376_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l376_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l376_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l376_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l377_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l377_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l377_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l377_2_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_2_valid;
  wire       [5:0]    _zz__zz_outputStreamArrayData_2_valid_1;
  wire       [6:0]    _zz__zz_5;
  reg                 _zz_outputStreamArrayData_2_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_2_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_2_payload;
  wire       [6:0]    _zz_outputStreamArrayData_2_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l383_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l383_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l383_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l384_2_3;
  wire       [7:0]    _zz_selectReadFifo_2;
  wire       [7:0]    _zz_selectReadFifo_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_2;
  wire       [12:0]   _zz_when_ArraySlice_l387_2_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l392_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l392_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l393_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l393_2_3;
  wire       [7:0]    _zz__zz_realValue1_0_6;
  wire       [7:0]    _zz__zz_realValue1_0_6_1;
  wire       [7:0]    _zz_realValue1_0_6_1;
  wire       [7:0]    _zz_realValue1_0_6_2;
  wire       [7:0]    _zz_realValue1_0_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l395_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l395_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_2;
  wire       [7:0]    _zz_selectReadFifo_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_4;
  wire       [0:0]    _zz_selectReadFifo_2_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_56;
  wire       [7:0]    _zz_when_ArraySlice_l158_56_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_56_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_56_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_56;
  wire       [7:0]    _zz_when_ArraySlice_l159_56_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_56_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_56_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_56_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_56_5;
  wire       [7:0]    _zz__zz_realValue_0_56;
  wire       [7:0]    _zz__zz_realValue_0_56_1;
  wire       [7:0]    _zz_realValue_0_56_1;
  wire       [7:0]    _zz_realValue_0_56_2;
  wire       [7:0]    _zz_realValue_0_56_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_56;
  wire       [7:0]    _zz_when_ArraySlice_l166_56_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_56_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_56_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_56_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_56_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_56_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_57;
  wire       [7:0]    _zz_when_ArraySlice_l158_57_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_57_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_57_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_57;
  wire       [6:0]    _zz_when_ArraySlice_l159_57_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_57_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_57_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_57_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_57_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_57_6;
  wire       [7:0]    _zz__zz_realValue_0_57;
  wire       [7:0]    _zz__zz_realValue_0_57_1;
  wire       [7:0]    _zz_realValue_0_57_1;
  wire       [7:0]    _zz_realValue_0_57_2;
  wire       [7:0]    _zz_realValue_0_57_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_57;
  wire       [6:0]    _zz_when_ArraySlice_l166_57_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_57_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_57_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_57_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_57_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_57_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_57_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_58;
  wire       [7:0]    _zz_when_ArraySlice_l158_58_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_58_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_58_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_58;
  wire       [6:0]    _zz_when_ArraySlice_l159_58_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_58_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_58_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_58_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_58_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_58_6;
  wire       [7:0]    _zz__zz_realValue_0_58;
  wire       [7:0]    _zz__zz_realValue_0_58_1;
  wire       [7:0]    _zz_realValue_0_58_1;
  wire       [7:0]    _zz_realValue_0_58_2;
  wire       [7:0]    _zz_realValue_0_58_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_58;
  wire       [6:0]    _zz_when_ArraySlice_l166_58_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_58_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_58_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_58_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_58_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_58_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_58_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_59;
  wire       [7:0]    _zz_when_ArraySlice_l158_59_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_59_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_59_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_59;
  wire       [6:0]    _zz_when_ArraySlice_l159_59_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_59_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_59_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_59_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_59_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_59_6;
  wire       [7:0]    _zz__zz_realValue_0_59;
  wire       [7:0]    _zz__zz_realValue_0_59_1;
  wire       [7:0]    _zz_realValue_0_59_1;
  wire       [7:0]    _zz_realValue_0_59_2;
  wire       [7:0]    _zz_realValue_0_59_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_59;
  wire       [6:0]    _zz_when_ArraySlice_l166_59_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_59_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_59_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_59_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_59_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_59_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_59_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_60;
  wire       [7:0]    _zz_when_ArraySlice_l158_60_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_60_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_60_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_60;
  wire       [6:0]    _zz_when_ArraySlice_l159_60_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_60_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_60_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_60_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_60_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_60_6;
  wire       [7:0]    _zz__zz_realValue_0_60;
  wire       [7:0]    _zz__zz_realValue_0_60_1;
  wire       [7:0]    _zz_realValue_0_60_1;
  wire       [7:0]    _zz_realValue_0_60_2;
  wire       [7:0]    _zz_realValue_0_60_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_60;
  wire       [6:0]    _zz_when_ArraySlice_l166_60_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_60_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_60_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_60_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_60_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_60_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_60_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_61;
  wire       [7:0]    _zz_when_ArraySlice_l158_61_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_61_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_61_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_61;
  wire       [5:0]    _zz_when_ArraySlice_l159_61_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_61_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_61_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_61_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_61_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_61_6;
  wire       [7:0]    _zz__zz_realValue_0_61;
  wire       [7:0]    _zz__zz_realValue_0_61_1;
  wire       [7:0]    _zz_realValue_0_61_1;
  wire       [7:0]    _zz_realValue_0_61_2;
  wire       [7:0]    _zz_realValue_0_61_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_61;
  wire       [5:0]    _zz_when_ArraySlice_l166_61_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_61_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_61_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_61_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_61_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_61_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_61_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_62;
  wire       [7:0]    _zz_when_ArraySlice_l158_62_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_62_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_62_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_62;
  wire       [5:0]    _zz_when_ArraySlice_l159_62_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_62_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_62_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_62_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_62_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_62_6;
  wire       [7:0]    _zz__zz_realValue_0_62;
  wire       [7:0]    _zz__zz_realValue_0_62_1;
  wire       [7:0]    _zz_realValue_0_62_1;
  wire       [7:0]    _zz_realValue_0_62_2;
  wire       [7:0]    _zz_realValue_0_62_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_62;
  wire       [5:0]    _zz_when_ArraySlice_l166_62_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_62_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_62_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_62_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_62_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_62_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_62_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_63;
  wire       [7:0]    _zz_when_ArraySlice_l158_63_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_63_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_63_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_63;
  wire       [4:0]    _zz_when_ArraySlice_l159_63_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_63_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_63_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_63_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_63_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_63_6;
  wire       [7:0]    _zz__zz_realValue_0_63;
  wire       [7:0]    _zz__zz_realValue_0_63_1;
  wire       [7:0]    _zz_realValue_0_63_1;
  wire       [7:0]    _zz_realValue_0_63_2;
  wire       [7:0]    _zz_realValue_0_63_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_63;
  wire       [4:0]    _zz_when_ArraySlice_l166_63_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_63_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_63_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_63_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_63_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_63_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_63_7;
  wire                _zz_when_ArraySlice_l400_2_1;
  wire                _zz_when_ArraySlice_l400_2_2;
  wire                _zz_when_ArraySlice_l400_2_3;
  wire                _zz_when_ArraySlice_l400_2_4;
  wire                _zz_when_ArraySlice_l400_2_5;
  wire                _zz_when_ArraySlice_l400_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_2_7;
  wire       [5:0]    _zz_when_ArraySlice_l403_2_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l406_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l406_2_5;
  wire       [7:0]    _zz_selectReadFifo_2_6;
  wire       [7:0]    _zz_selectReadFifo_2_7;
  wire       [6:0]    _zz_selectReadFifo_2_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_2;
  wire       [12:0]   _zz_when_ArraySlice_l413_2_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l417_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l417_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l417_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l418_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l418_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l418_2_5;
  wire       [7:0]    _zz__zz_realValue1_0_7;
  wire       [7:0]    _zz__zz_realValue1_0_7_1;
  wire       [7:0]    _zz_realValue1_0_7_1;
  wire       [7:0]    _zz_realValue1_0_7_2;
  wire       [7:0]    _zz_realValue1_0_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l420_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l420_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_9;
  wire       [7:0]    _zz_selectReadFifo_2_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_64;
  wire       [7:0]    _zz_when_ArraySlice_l158_64_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_64_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_64_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_64;
  wire       [7:0]    _zz_when_ArraySlice_l159_64_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_64_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_64_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_64_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_64_5;
  wire       [7:0]    _zz__zz_realValue_0_64;
  wire       [7:0]    _zz__zz_realValue_0_64_1;
  wire       [7:0]    _zz_realValue_0_64_1;
  wire       [7:0]    _zz_realValue_0_64_2;
  wire       [7:0]    _zz_realValue_0_64_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_64;
  wire       [7:0]    _zz_when_ArraySlice_l166_64_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_64_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_64_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_64_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_64_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_64_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_65;
  wire       [7:0]    _zz_when_ArraySlice_l158_65_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_65_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_65_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_65;
  wire       [6:0]    _zz_when_ArraySlice_l159_65_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_65_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_65_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_65_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_65_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_65_6;
  wire       [7:0]    _zz__zz_realValue_0_65;
  wire       [7:0]    _zz__zz_realValue_0_65_1;
  wire       [7:0]    _zz_realValue_0_65_1;
  wire       [7:0]    _zz_realValue_0_65_2;
  wire       [7:0]    _zz_realValue_0_65_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_65;
  wire       [6:0]    _zz_when_ArraySlice_l166_65_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_65_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_65_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_65_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_65_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_65_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_65_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_66;
  wire       [7:0]    _zz_when_ArraySlice_l158_66_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_66_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_66_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_66;
  wire       [6:0]    _zz_when_ArraySlice_l159_66_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_66_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_66_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_66_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_66_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_66_6;
  wire       [7:0]    _zz__zz_realValue_0_66;
  wire       [7:0]    _zz__zz_realValue_0_66_1;
  wire       [7:0]    _zz_realValue_0_66_1;
  wire       [7:0]    _zz_realValue_0_66_2;
  wire       [7:0]    _zz_realValue_0_66_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_66;
  wire       [6:0]    _zz_when_ArraySlice_l166_66_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_66_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_66_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_66_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_66_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_66_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_66_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_67;
  wire       [7:0]    _zz_when_ArraySlice_l158_67_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_67_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_67_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_67;
  wire       [6:0]    _zz_when_ArraySlice_l159_67_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_67_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_67_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_67_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_67_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_67_6;
  wire       [7:0]    _zz__zz_realValue_0_67;
  wire       [7:0]    _zz__zz_realValue_0_67_1;
  wire       [7:0]    _zz_realValue_0_67_1;
  wire       [7:0]    _zz_realValue_0_67_2;
  wire       [7:0]    _zz_realValue_0_67_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_67;
  wire       [6:0]    _zz_when_ArraySlice_l166_67_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_67_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_67_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_67_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_67_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_67_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_67_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_68;
  wire       [7:0]    _zz_when_ArraySlice_l158_68_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_68_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_68_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_68;
  wire       [6:0]    _zz_when_ArraySlice_l159_68_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_68_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_68_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_68_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_68_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_68_6;
  wire       [7:0]    _zz__zz_realValue_0_68;
  wire       [7:0]    _zz__zz_realValue_0_68_1;
  wire       [7:0]    _zz_realValue_0_68_1;
  wire       [7:0]    _zz_realValue_0_68_2;
  wire       [7:0]    _zz_realValue_0_68_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_68;
  wire       [6:0]    _zz_when_ArraySlice_l166_68_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_68_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_68_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_68_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_68_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_68_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_68_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_69;
  wire       [7:0]    _zz_when_ArraySlice_l158_69_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_69_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_69_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_69;
  wire       [5:0]    _zz_when_ArraySlice_l159_69_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_69_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_69_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_69_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_69_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_69_6;
  wire       [7:0]    _zz__zz_realValue_0_69;
  wire       [7:0]    _zz__zz_realValue_0_69_1;
  wire       [7:0]    _zz_realValue_0_69_1;
  wire       [7:0]    _zz_realValue_0_69_2;
  wire       [7:0]    _zz_realValue_0_69_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_69;
  wire       [5:0]    _zz_when_ArraySlice_l166_69_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_69_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_69_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_69_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_69_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_69_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_69_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_70;
  wire       [7:0]    _zz_when_ArraySlice_l158_70_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_70_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_70_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_70;
  wire       [5:0]    _zz_when_ArraySlice_l159_70_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_70_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_70_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_70_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_70_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_70_6;
  wire       [7:0]    _zz__zz_realValue_0_70;
  wire       [7:0]    _zz__zz_realValue_0_70_1;
  wire       [7:0]    _zz_realValue_0_70_1;
  wire       [7:0]    _zz_realValue_0_70_2;
  wire       [7:0]    _zz_realValue_0_70_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_70;
  wire       [5:0]    _zz_when_ArraySlice_l166_70_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_70_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_70_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_70_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_70_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_70_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_70_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_71;
  wire       [7:0]    _zz_when_ArraySlice_l158_71_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_71_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_71_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_71;
  wire       [4:0]    _zz_when_ArraySlice_l159_71_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_71_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_71_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_71_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_71_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_71_6;
  wire       [7:0]    _zz__zz_realValue_0_71;
  wire       [7:0]    _zz__zz_realValue_0_71_1;
  wire       [7:0]    _zz_realValue_0_71_1;
  wire       [7:0]    _zz_realValue_0_71_2;
  wire       [7:0]    _zz_realValue_0_71_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_71;
  wire       [4:0]    _zz_when_ArraySlice_l166_71_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_71_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_71_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_71_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_71_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_71_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_71_7;
  wire                _zz_when_ArraySlice_l425_2_1;
  wire                _zz_when_ArraySlice_l425_2_2;
  wire                _zz_when_ArraySlice_l425_2_3;
  wire                _zz_when_ArraySlice_l425_2_4;
  wire                _zz_when_ArraySlice_l425_2_5;
  wire                _zz_when_ArraySlice_l425_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_2_7;
  wire       [5:0]    _zz_when_ArraySlice_l428_2_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l431_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l431_2_5;
  wire       [7:0]    _zz_selectReadFifo_2_11;
  wire       [7:0]    _zz_selectReadFifo_2_12;
  wire       [6:0]    _zz_selectReadFifo_2_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_2;
  wire       [12:0]   _zz_when_ArraySlice_l438_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l449_2_3;
  wire       [7:0]    _zz__zz_realValue1_0_8;
  wire       [7:0]    _zz__zz_realValue1_0_8_1;
  wire       [7:0]    _zz_realValue1_0_8_1;
  wire       [7:0]    _zz_realValue1_0_8_2;
  wire       [7:0]    _zz_realValue1_0_8_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l450_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l450_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_14;
  wire       [7:0]    _zz_selectReadFifo_2_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_72;
  wire       [7:0]    _zz_when_ArraySlice_l158_72_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_72_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_72_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_72;
  wire       [7:0]    _zz_when_ArraySlice_l159_72_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_72_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_72_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_72_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_72_5;
  wire       [7:0]    _zz__zz_realValue_0_72;
  wire       [7:0]    _zz__zz_realValue_0_72_1;
  wire       [7:0]    _zz_realValue_0_72_1;
  wire       [7:0]    _zz_realValue_0_72_2;
  wire       [7:0]    _zz_realValue_0_72_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_72;
  wire       [7:0]    _zz_when_ArraySlice_l166_72_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_72_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_72_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_72_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_72_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_72_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_73;
  wire       [7:0]    _zz_when_ArraySlice_l158_73_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_73_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_73_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_73;
  wire       [6:0]    _zz_when_ArraySlice_l159_73_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_73_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_73_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_73_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_73_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_73_6;
  wire       [7:0]    _zz__zz_realValue_0_73;
  wire       [7:0]    _zz__zz_realValue_0_73_1;
  wire       [7:0]    _zz_realValue_0_73_1;
  wire       [7:0]    _zz_realValue_0_73_2;
  wire       [7:0]    _zz_realValue_0_73_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_73;
  wire       [6:0]    _zz_when_ArraySlice_l166_73_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_73_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_73_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_73_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_73_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_73_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_73_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_74;
  wire       [7:0]    _zz_when_ArraySlice_l158_74_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_74_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_74_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_74;
  wire       [6:0]    _zz_when_ArraySlice_l159_74_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_74_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_74_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_74_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_74_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_74_6;
  wire       [7:0]    _zz__zz_realValue_0_74;
  wire       [7:0]    _zz__zz_realValue_0_74_1;
  wire       [7:0]    _zz_realValue_0_74_1;
  wire       [7:0]    _zz_realValue_0_74_2;
  wire       [7:0]    _zz_realValue_0_74_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_74;
  wire       [6:0]    _zz_when_ArraySlice_l166_74_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_74_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_74_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_74_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_74_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_74_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_74_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_75;
  wire       [7:0]    _zz_when_ArraySlice_l158_75_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_75_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_75_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_75;
  wire       [6:0]    _zz_when_ArraySlice_l159_75_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_75_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_75_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_75_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_75_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_75_6;
  wire       [7:0]    _zz__zz_realValue_0_75;
  wire       [7:0]    _zz__zz_realValue_0_75_1;
  wire       [7:0]    _zz_realValue_0_75_1;
  wire       [7:0]    _zz_realValue_0_75_2;
  wire       [7:0]    _zz_realValue_0_75_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_75;
  wire       [6:0]    _zz_when_ArraySlice_l166_75_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_75_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_75_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_75_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_75_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_75_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_75_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_76;
  wire       [7:0]    _zz_when_ArraySlice_l158_76_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_76_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_76_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_76;
  wire       [6:0]    _zz_when_ArraySlice_l159_76_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_76_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_76_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_76_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_76_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_76_6;
  wire       [7:0]    _zz__zz_realValue_0_76;
  wire       [7:0]    _zz__zz_realValue_0_76_1;
  wire       [7:0]    _zz_realValue_0_76_1;
  wire       [7:0]    _zz_realValue_0_76_2;
  wire       [7:0]    _zz_realValue_0_76_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_76;
  wire       [6:0]    _zz_when_ArraySlice_l166_76_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_76_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_76_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_76_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_76_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_76_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_76_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_77;
  wire       [7:0]    _zz_when_ArraySlice_l158_77_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_77_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_77_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_77;
  wire       [5:0]    _zz_when_ArraySlice_l159_77_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_77_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_77_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_77_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_77_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_77_6;
  wire       [7:0]    _zz__zz_realValue_0_77;
  wire       [7:0]    _zz__zz_realValue_0_77_1;
  wire       [7:0]    _zz_realValue_0_77_1;
  wire       [7:0]    _zz_realValue_0_77_2;
  wire       [7:0]    _zz_realValue_0_77_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_77;
  wire       [5:0]    _zz_when_ArraySlice_l166_77_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_77_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_77_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_77_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_77_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_77_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_77_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_78;
  wire       [7:0]    _zz_when_ArraySlice_l158_78_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_78_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_78_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_78;
  wire       [5:0]    _zz_when_ArraySlice_l159_78_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_78_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_78_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_78_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_78_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_78_6;
  wire       [7:0]    _zz__zz_realValue_0_78;
  wire       [7:0]    _zz__zz_realValue_0_78_1;
  wire       [7:0]    _zz_realValue_0_78_1;
  wire       [7:0]    _zz_realValue_0_78_2;
  wire       [7:0]    _zz_realValue_0_78_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_78;
  wire       [5:0]    _zz_when_ArraySlice_l166_78_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_78_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_78_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_78_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_78_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_78_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_78_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_79;
  wire       [7:0]    _zz_when_ArraySlice_l158_79_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_79_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_79_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_79;
  wire       [4:0]    _zz_when_ArraySlice_l159_79_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_79_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_79_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_79_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_79_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_79_6;
  wire       [7:0]    _zz__zz_realValue_0_79;
  wire       [7:0]    _zz__zz_realValue_0_79_1;
  wire       [7:0]    _zz_realValue_0_79_1;
  wire       [7:0]    _zz_realValue_0_79_2;
  wire       [7:0]    _zz_realValue_0_79_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_79;
  wire       [4:0]    _zz_when_ArraySlice_l166_79_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_79_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_79_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_79_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_79_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_79_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_79_7;
  wire                _zz_when_ArraySlice_l457_2_1;
  wire                _zz_when_ArraySlice_l457_2_2;
  wire                _zz_when_ArraySlice_l457_2_3;
  wire                _zz_when_ArraySlice_l457_2_4;
  wire                _zz_when_ArraySlice_l457_2_5;
  wire                _zz_when_ArraySlice_l457_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_2;
  wire       [12:0]   _zz_when_ArraySlice_l461_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l447_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l447_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l468_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l468_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l376_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l376_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l376_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l376_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l377_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l377_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l377_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l377_3_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_3_valid;
  wire       [5:0]    _zz__zz_outputStreamArrayData_3_valid_1;
  wire       [6:0]    _zz__zz_6;
  reg                 _zz_outputStreamArrayData_3_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_3_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_3_payload;
  wire       [6:0]    _zz_outputStreamArrayData_3_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l383_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l383_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l383_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_3;
  wire       [7:0]    _zz_when_ArraySlice_l384_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_3_2;
  wire       [7:0]    _zz_selectReadFifo_3;
  wire       [7:0]    _zz_selectReadFifo_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_3;
  wire       [12:0]   _zz_when_ArraySlice_l387_3_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l392_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l392_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l393_3;
  wire       [7:0]    _zz_when_ArraySlice_l393_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_3_2;
  wire       [7:0]    _zz__zz_realValue1_0_9;
  wire       [7:0]    _zz__zz_realValue1_0_9_1;
  wire       [7:0]    _zz_realValue1_0_9_1;
  wire       [7:0]    _zz_realValue1_0_9_2;
  wire       [7:0]    _zz_realValue1_0_9_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_3;
  wire       [6:0]    _zz_when_ArraySlice_l395_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_3;
  wire       [7:0]    _zz_selectReadFifo_3_4;
  wire       [0:0]    _zz_selectReadFifo_3_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_80;
  wire       [7:0]    _zz_when_ArraySlice_l158_80_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_80_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_80_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_80;
  wire       [7:0]    _zz_when_ArraySlice_l159_80_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_80_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_80_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_80_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_80_5;
  wire       [7:0]    _zz__zz_realValue_0_80;
  wire       [7:0]    _zz__zz_realValue_0_80_1;
  wire       [7:0]    _zz_realValue_0_80_1;
  wire       [7:0]    _zz_realValue_0_80_2;
  wire       [7:0]    _zz_realValue_0_80_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_80;
  wire       [7:0]    _zz_when_ArraySlice_l166_80_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_80_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_80_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_80_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_80_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_80_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_81;
  wire       [7:0]    _zz_when_ArraySlice_l158_81_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_81_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_81_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_81;
  wire       [6:0]    _zz_when_ArraySlice_l159_81_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_81_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_81_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_81_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_81_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_81_6;
  wire       [7:0]    _zz__zz_realValue_0_81;
  wire       [7:0]    _zz__zz_realValue_0_81_1;
  wire       [7:0]    _zz_realValue_0_81_1;
  wire       [7:0]    _zz_realValue_0_81_2;
  wire       [7:0]    _zz_realValue_0_81_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_81;
  wire       [6:0]    _zz_when_ArraySlice_l166_81_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_81_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_81_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_81_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_81_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_81_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_81_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_82;
  wire       [7:0]    _zz_when_ArraySlice_l158_82_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_82_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_82_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_82;
  wire       [6:0]    _zz_when_ArraySlice_l159_82_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_82_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_82_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_82_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_82_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_82_6;
  wire       [7:0]    _zz__zz_realValue_0_82;
  wire       [7:0]    _zz__zz_realValue_0_82_1;
  wire       [7:0]    _zz_realValue_0_82_1;
  wire       [7:0]    _zz_realValue_0_82_2;
  wire       [7:0]    _zz_realValue_0_82_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_82;
  wire       [6:0]    _zz_when_ArraySlice_l166_82_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_82_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_82_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_82_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_82_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_82_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_82_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_83;
  wire       [7:0]    _zz_when_ArraySlice_l158_83_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_83_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_83_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_83;
  wire       [6:0]    _zz_when_ArraySlice_l159_83_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_83_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_83_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_83_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_83_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_83_6;
  wire       [7:0]    _zz__zz_realValue_0_83;
  wire       [7:0]    _zz__zz_realValue_0_83_1;
  wire       [7:0]    _zz_realValue_0_83_1;
  wire       [7:0]    _zz_realValue_0_83_2;
  wire       [7:0]    _zz_realValue_0_83_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_83;
  wire       [6:0]    _zz_when_ArraySlice_l166_83_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_83_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_83_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_83_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_83_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_83_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_83_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_84;
  wire       [7:0]    _zz_when_ArraySlice_l158_84_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_84_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_84_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_84;
  wire       [6:0]    _zz_when_ArraySlice_l159_84_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_84_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_84_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_84_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_84_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_84_6;
  wire       [7:0]    _zz__zz_realValue_0_84;
  wire       [7:0]    _zz__zz_realValue_0_84_1;
  wire       [7:0]    _zz_realValue_0_84_1;
  wire       [7:0]    _zz_realValue_0_84_2;
  wire       [7:0]    _zz_realValue_0_84_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_84;
  wire       [6:0]    _zz_when_ArraySlice_l166_84_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_84_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_84_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_84_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_84_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_84_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_84_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_85;
  wire       [7:0]    _zz_when_ArraySlice_l158_85_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_85_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_85_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_85;
  wire       [5:0]    _zz_when_ArraySlice_l159_85_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_85_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_85_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_85_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_85_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_85_6;
  wire       [7:0]    _zz__zz_realValue_0_85;
  wire       [7:0]    _zz__zz_realValue_0_85_1;
  wire       [7:0]    _zz_realValue_0_85_1;
  wire       [7:0]    _zz_realValue_0_85_2;
  wire       [7:0]    _zz_realValue_0_85_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_85;
  wire       [5:0]    _zz_when_ArraySlice_l166_85_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_85_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_85_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_85_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_85_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_85_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_85_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_86;
  wire       [7:0]    _zz_when_ArraySlice_l158_86_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_86_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_86_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_86;
  wire       [5:0]    _zz_when_ArraySlice_l159_86_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_86_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_86_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_86_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_86_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_86_6;
  wire       [7:0]    _zz__zz_realValue_0_86;
  wire       [7:0]    _zz__zz_realValue_0_86_1;
  wire       [7:0]    _zz_realValue_0_86_1;
  wire       [7:0]    _zz_realValue_0_86_2;
  wire       [7:0]    _zz_realValue_0_86_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_86;
  wire       [5:0]    _zz_when_ArraySlice_l166_86_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_86_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_86_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_86_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_86_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_86_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_86_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_87;
  wire       [7:0]    _zz_when_ArraySlice_l158_87_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_87_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_87_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_87;
  wire       [4:0]    _zz_when_ArraySlice_l159_87_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_87_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_87_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_87_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_87_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_87_6;
  wire       [7:0]    _zz__zz_realValue_0_87;
  wire       [7:0]    _zz__zz_realValue_0_87_1;
  wire       [7:0]    _zz_realValue_0_87_1;
  wire       [7:0]    _zz_realValue_0_87_2;
  wire       [7:0]    _zz_realValue_0_87_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_87;
  wire       [4:0]    _zz_when_ArraySlice_l166_87_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_87_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_87_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_87_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_87_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_87_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_87_7;
  wire                _zz_when_ArraySlice_l400_3_1;
  wire                _zz_when_ArraySlice_l400_3_2;
  wire                _zz_when_ArraySlice_l400_3_3;
  wire                _zz_when_ArraySlice_l400_3_4;
  wire                _zz_when_ArraySlice_l400_3_5;
  wire                _zz_when_ArraySlice_l400_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_3_7;
  wire       [5:0]    _zz_when_ArraySlice_l403_3_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l406_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l406_3_5;
  wire       [7:0]    _zz_selectReadFifo_3_6;
  wire       [7:0]    _zz_selectReadFifo_3_7;
  wire       [6:0]    _zz_selectReadFifo_3_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_3;
  wire       [12:0]   _zz_when_ArraySlice_l413_3_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l417_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l417_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l417_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l418_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l418_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l418_3_5;
  wire       [7:0]    _zz__zz_realValue1_0_10;
  wire       [7:0]    _zz__zz_realValue1_0_10_1;
  wire       [7:0]    _zz_realValue1_0_10_1;
  wire       [7:0]    _zz_realValue1_0_10_2;
  wire       [7:0]    _zz_realValue1_0_10_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_3;
  wire       [6:0]    _zz_when_ArraySlice_l420_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_9;
  wire       [7:0]    _zz_selectReadFifo_3_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_88;
  wire       [7:0]    _zz_when_ArraySlice_l158_88_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_88_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_88_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_88;
  wire       [7:0]    _zz_when_ArraySlice_l159_88_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_88_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_88_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_88_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_88_5;
  wire       [7:0]    _zz__zz_realValue_0_88;
  wire       [7:0]    _zz__zz_realValue_0_88_1;
  wire       [7:0]    _zz_realValue_0_88_1;
  wire       [7:0]    _zz_realValue_0_88_2;
  wire       [7:0]    _zz_realValue_0_88_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_88;
  wire       [7:0]    _zz_when_ArraySlice_l166_88_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_88_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_88_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_88_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_88_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_88_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_89;
  wire       [7:0]    _zz_when_ArraySlice_l158_89_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_89_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_89_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_89;
  wire       [6:0]    _zz_when_ArraySlice_l159_89_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_89_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_89_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_89_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_89_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_89_6;
  wire       [7:0]    _zz__zz_realValue_0_89;
  wire       [7:0]    _zz__zz_realValue_0_89_1;
  wire       [7:0]    _zz_realValue_0_89_1;
  wire       [7:0]    _zz_realValue_0_89_2;
  wire       [7:0]    _zz_realValue_0_89_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_89;
  wire       [6:0]    _zz_when_ArraySlice_l166_89_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_89_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_89_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_89_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_89_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_89_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_89_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_90;
  wire       [7:0]    _zz_when_ArraySlice_l158_90_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_90_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_90_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_90;
  wire       [6:0]    _zz_when_ArraySlice_l159_90_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_90_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_90_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_90_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_90_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_90_6;
  wire       [7:0]    _zz__zz_realValue_0_90;
  wire       [7:0]    _zz__zz_realValue_0_90_1;
  wire       [7:0]    _zz_realValue_0_90_1;
  wire       [7:0]    _zz_realValue_0_90_2;
  wire       [7:0]    _zz_realValue_0_90_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_90;
  wire       [6:0]    _zz_when_ArraySlice_l166_90_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_90_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_90_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_90_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_90_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_90_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_90_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_91;
  wire       [7:0]    _zz_when_ArraySlice_l158_91_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_91_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_91_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_91;
  wire       [6:0]    _zz_when_ArraySlice_l159_91_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_91_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_91_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_91_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_91_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_91_6;
  wire       [7:0]    _zz__zz_realValue_0_91;
  wire       [7:0]    _zz__zz_realValue_0_91_1;
  wire       [7:0]    _zz_realValue_0_91_1;
  wire       [7:0]    _zz_realValue_0_91_2;
  wire       [7:0]    _zz_realValue_0_91_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_91;
  wire       [6:0]    _zz_when_ArraySlice_l166_91_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_91_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_91_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_91_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_91_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_91_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_91_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_92;
  wire       [7:0]    _zz_when_ArraySlice_l158_92_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_92_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_92_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_92;
  wire       [6:0]    _zz_when_ArraySlice_l159_92_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_92_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_92_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_92_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_92_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_92_6;
  wire       [7:0]    _zz__zz_realValue_0_92;
  wire       [7:0]    _zz__zz_realValue_0_92_1;
  wire       [7:0]    _zz_realValue_0_92_1;
  wire       [7:0]    _zz_realValue_0_92_2;
  wire       [7:0]    _zz_realValue_0_92_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_92;
  wire       [6:0]    _zz_when_ArraySlice_l166_92_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_92_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_92_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_92_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_92_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_92_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_92_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_93;
  wire       [7:0]    _zz_when_ArraySlice_l158_93_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_93_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_93_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_93;
  wire       [5:0]    _zz_when_ArraySlice_l159_93_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_93_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_93_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_93_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_93_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_93_6;
  wire       [7:0]    _zz__zz_realValue_0_93;
  wire       [7:0]    _zz__zz_realValue_0_93_1;
  wire       [7:0]    _zz_realValue_0_93_1;
  wire       [7:0]    _zz_realValue_0_93_2;
  wire       [7:0]    _zz_realValue_0_93_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_93;
  wire       [5:0]    _zz_when_ArraySlice_l166_93_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_93_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_93_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_93_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_93_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_93_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_93_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_94;
  wire       [7:0]    _zz_when_ArraySlice_l158_94_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_94_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_94_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_94;
  wire       [5:0]    _zz_when_ArraySlice_l159_94_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_94_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_94_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_94_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_94_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_94_6;
  wire       [7:0]    _zz__zz_realValue_0_94;
  wire       [7:0]    _zz__zz_realValue_0_94_1;
  wire       [7:0]    _zz_realValue_0_94_1;
  wire       [7:0]    _zz_realValue_0_94_2;
  wire       [7:0]    _zz_realValue_0_94_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_94;
  wire       [5:0]    _zz_when_ArraySlice_l166_94_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_94_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_94_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_94_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_94_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_94_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_94_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_95;
  wire       [7:0]    _zz_when_ArraySlice_l158_95_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_95_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_95_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_95;
  wire       [4:0]    _zz_when_ArraySlice_l159_95_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_95_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_95_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_95_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_95_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_95_6;
  wire       [7:0]    _zz__zz_realValue_0_95;
  wire       [7:0]    _zz__zz_realValue_0_95_1;
  wire       [7:0]    _zz_realValue_0_95_1;
  wire       [7:0]    _zz_realValue_0_95_2;
  wire       [7:0]    _zz_realValue_0_95_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_95;
  wire       [4:0]    _zz_when_ArraySlice_l166_95_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_95_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_95_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_95_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_95_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_95_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_95_7;
  wire                _zz_when_ArraySlice_l425_3_1;
  wire                _zz_when_ArraySlice_l425_3_2;
  wire                _zz_when_ArraySlice_l425_3_3;
  wire                _zz_when_ArraySlice_l425_3_4;
  wire                _zz_when_ArraySlice_l425_3_5;
  wire                _zz_when_ArraySlice_l425_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_3_7;
  wire       [5:0]    _zz_when_ArraySlice_l428_3_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l431_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l431_3_5;
  wire       [7:0]    _zz_selectReadFifo_3_11;
  wire       [7:0]    _zz_selectReadFifo_3_12;
  wire       [6:0]    _zz_selectReadFifo_3_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_3;
  wire       [12:0]   _zz_when_ArraySlice_l438_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_3;
  wire       [7:0]    _zz_when_ArraySlice_l449_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_3_2;
  wire       [7:0]    _zz__zz_realValue1_0_11;
  wire       [7:0]    _zz__zz_realValue1_0_11_1;
  wire       [7:0]    _zz_realValue1_0_11_1;
  wire       [7:0]    _zz_realValue1_0_11_2;
  wire       [7:0]    _zz_realValue1_0_11_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_3;
  wire       [6:0]    _zz_when_ArraySlice_l450_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_14;
  wire       [7:0]    _zz_selectReadFifo_3_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_96;
  wire       [7:0]    _zz_when_ArraySlice_l158_96_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_96_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_96_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_96;
  wire       [7:0]    _zz_when_ArraySlice_l159_96_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_96_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_96_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_96_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_96_5;
  wire       [7:0]    _zz__zz_realValue_0_96;
  wire       [7:0]    _zz__zz_realValue_0_96_1;
  wire       [7:0]    _zz_realValue_0_96_1;
  wire       [7:0]    _zz_realValue_0_96_2;
  wire       [7:0]    _zz_realValue_0_96_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_96;
  wire       [7:0]    _zz_when_ArraySlice_l166_96_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_96_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_96_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_96_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_96_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_96_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_97;
  wire       [7:0]    _zz_when_ArraySlice_l158_97_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_97_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_97_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_97;
  wire       [6:0]    _zz_when_ArraySlice_l159_97_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_97_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_97_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_97_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_97_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_97_6;
  wire       [7:0]    _zz__zz_realValue_0_97;
  wire       [7:0]    _zz__zz_realValue_0_97_1;
  wire       [7:0]    _zz_realValue_0_97_1;
  wire       [7:0]    _zz_realValue_0_97_2;
  wire       [7:0]    _zz_realValue_0_97_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_97;
  wire       [6:0]    _zz_when_ArraySlice_l166_97_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_97_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_97_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_97_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_97_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_97_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_97_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_98;
  wire       [7:0]    _zz_when_ArraySlice_l158_98_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_98_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_98_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_98;
  wire       [6:0]    _zz_when_ArraySlice_l159_98_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_98_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_98_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_98_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_98_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_98_6;
  wire       [7:0]    _zz__zz_realValue_0_98;
  wire       [7:0]    _zz__zz_realValue_0_98_1;
  wire       [7:0]    _zz_realValue_0_98_1;
  wire       [7:0]    _zz_realValue_0_98_2;
  wire       [7:0]    _zz_realValue_0_98_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_98;
  wire       [6:0]    _zz_when_ArraySlice_l166_98_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_98_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_98_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_98_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_98_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_98_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_98_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_99;
  wire       [7:0]    _zz_when_ArraySlice_l158_99_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_99_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_99_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_99;
  wire       [6:0]    _zz_when_ArraySlice_l159_99_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_99_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_99_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_99_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_99_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_99_6;
  wire       [7:0]    _zz__zz_realValue_0_99;
  wire       [7:0]    _zz__zz_realValue_0_99_1;
  wire       [7:0]    _zz_realValue_0_99_1;
  wire       [7:0]    _zz_realValue_0_99_2;
  wire       [7:0]    _zz_realValue_0_99_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_99;
  wire       [6:0]    _zz_when_ArraySlice_l166_99_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_99_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_99_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_99_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_99_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_99_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_99_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_100;
  wire       [7:0]    _zz_when_ArraySlice_l158_100_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_100_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_100_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_100;
  wire       [6:0]    _zz_when_ArraySlice_l159_100_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_100_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_100_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_100_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_100_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_100_6;
  wire       [7:0]    _zz__zz_realValue_0_100;
  wire       [7:0]    _zz__zz_realValue_0_100_1;
  wire       [7:0]    _zz_realValue_0_100_1;
  wire       [7:0]    _zz_realValue_0_100_2;
  wire       [7:0]    _zz_realValue_0_100_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_100;
  wire       [6:0]    _zz_when_ArraySlice_l166_100_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_100_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_100_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_100_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_100_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_100_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_100_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_101;
  wire       [7:0]    _zz_when_ArraySlice_l158_101_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_101_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_101_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_101;
  wire       [5:0]    _zz_when_ArraySlice_l159_101_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_101_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_101_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_101_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_101_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_101_6;
  wire       [7:0]    _zz__zz_realValue_0_101;
  wire       [7:0]    _zz__zz_realValue_0_101_1;
  wire       [7:0]    _zz_realValue_0_101_1;
  wire       [7:0]    _zz_realValue_0_101_2;
  wire       [7:0]    _zz_realValue_0_101_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_101;
  wire       [5:0]    _zz_when_ArraySlice_l166_101_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_101_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_101_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_101_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_101_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_101_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_101_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_102;
  wire       [7:0]    _zz_when_ArraySlice_l158_102_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_102_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_102_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_102;
  wire       [5:0]    _zz_when_ArraySlice_l159_102_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_102_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_102_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_102_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_102_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_102_6;
  wire       [7:0]    _zz__zz_realValue_0_102;
  wire       [7:0]    _zz__zz_realValue_0_102_1;
  wire       [7:0]    _zz_realValue_0_102_1;
  wire       [7:0]    _zz_realValue_0_102_2;
  wire       [7:0]    _zz_realValue_0_102_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_102;
  wire       [5:0]    _zz_when_ArraySlice_l166_102_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_102_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_102_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_102_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_102_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_102_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_102_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_103;
  wire       [7:0]    _zz_when_ArraySlice_l158_103_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_103_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_103_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_103;
  wire       [4:0]    _zz_when_ArraySlice_l159_103_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_103_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_103_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_103_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_103_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_103_6;
  wire       [7:0]    _zz__zz_realValue_0_103;
  wire       [7:0]    _zz__zz_realValue_0_103_1;
  wire       [7:0]    _zz_realValue_0_103_1;
  wire       [7:0]    _zz_realValue_0_103_2;
  wire       [7:0]    _zz_realValue_0_103_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_103;
  wire       [4:0]    _zz_when_ArraySlice_l166_103_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_103_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_103_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_103_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_103_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_103_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_103_7;
  wire                _zz_when_ArraySlice_l457_3_1;
  wire                _zz_when_ArraySlice_l457_3_2;
  wire                _zz_when_ArraySlice_l457_3_3;
  wire                _zz_when_ArraySlice_l457_3_4;
  wire                _zz_when_ArraySlice_l457_3_5;
  wire                _zz_when_ArraySlice_l457_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_3;
  wire       [12:0]   _zz_when_ArraySlice_l461_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l447_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l447_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l468_3;
  wire       [7:0]    _zz_when_ArraySlice_l468_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_4;
  wire       [7:0]    _zz_when_ArraySlice_l376_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l376_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l377_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l377_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l377_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l377_4_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_4_valid;
  wire       [6:0]    _zz__zz_outputStreamArrayData_4_valid_1;
  wire       [6:0]    _zz__zz_7;
  reg                 _zz_outputStreamArrayData_4_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_4_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_4_payload;
  wire       [6:0]    _zz_outputStreamArrayData_4_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l383_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l383_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l383_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l384_4;
  wire       [7:0]    _zz_when_ArraySlice_l384_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_4_2;
  wire       [7:0]    _zz_selectReadFifo_4;
  wire       [7:0]    _zz_selectReadFifo_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_4;
  wire       [12:0]   _zz_when_ArraySlice_l387_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l392_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l392_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l392_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l393_4;
  wire       [7:0]    _zz_when_ArraySlice_l393_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_4_2;
  wire       [7:0]    _zz__zz_realValue1_0_12;
  wire       [7:0]    _zz__zz_realValue1_0_12_1;
  wire       [7:0]    _zz_realValue1_0_12_1;
  wire       [7:0]    _zz_realValue1_0_12_2;
  wire       [7:0]    _zz_realValue1_0_12_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_4;
  wire       [6:0]    _zz_when_ArraySlice_l395_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_3;
  wire       [7:0]    _zz_selectReadFifo_4_4;
  wire       [0:0]    _zz_selectReadFifo_4_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_104;
  wire       [7:0]    _zz_when_ArraySlice_l158_104_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_104_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_104_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_104;
  wire       [7:0]    _zz_when_ArraySlice_l159_104_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_104_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_104_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_104_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_104_5;
  wire       [7:0]    _zz__zz_realValue_0_104;
  wire       [7:0]    _zz__zz_realValue_0_104_1;
  wire       [7:0]    _zz_realValue_0_104_1;
  wire       [7:0]    _zz_realValue_0_104_2;
  wire       [7:0]    _zz_realValue_0_104_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_104;
  wire       [7:0]    _zz_when_ArraySlice_l166_104_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_104_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_104_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_104_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_104_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_104_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_105;
  wire       [7:0]    _zz_when_ArraySlice_l158_105_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_105_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_105_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_105;
  wire       [6:0]    _zz_when_ArraySlice_l159_105_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_105_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_105_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_105_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_105_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_105_6;
  wire       [7:0]    _zz__zz_realValue_0_105;
  wire       [7:0]    _zz__zz_realValue_0_105_1;
  wire       [7:0]    _zz_realValue_0_105_1;
  wire       [7:0]    _zz_realValue_0_105_2;
  wire       [7:0]    _zz_realValue_0_105_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_105;
  wire       [6:0]    _zz_when_ArraySlice_l166_105_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_105_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_105_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_105_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_105_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_105_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_105_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_106;
  wire       [7:0]    _zz_when_ArraySlice_l158_106_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_106_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_106_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_106;
  wire       [6:0]    _zz_when_ArraySlice_l159_106_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_106_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_106_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_106_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_106_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_106_6;
  wire       [7:0]    _zz__zz_realValue_0_106;
  wire       [7:0]    _zz__zz_realValue_0_106_1;
  wire       [7:0]    _zz_realValue_0_106_1;
  wire       [7:0]    _zz_realValue_0_106_2;
  wire       [7:0]    _zz_realValue_0_106_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_106;
  wire       [6:0]    _zz_when_ArraySlice_l166_106_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_106_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_106_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_106_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_106_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_106_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_106_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_107;
  wire       [7:0]    _zz_when_ArraySlice_l158_107_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_107_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_107_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_107;
  wire       [6:0]    _zz_when_ArraySlice_l159_107_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_107_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_107_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_107_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_107_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_107_6;
  wire       [7:0]    _zz__zz_realValue_0_107;
  wire       [7:0]    _zz__zz_realValue_0_107_1;
  wire       [7:0]    _zz_realValue_0_107_1;
  wire       [7:0]    _zz_realValue_0_107_2;
  wire       [7:0]    _zz_realValue_0_107_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_107;
  wire       [6:0]    _zz_when_ArraySlice_l166_107_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_107_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_107_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_107_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_107_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_107_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_107_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_108;
  wire       [7:0]    _zz_when_ArraySlice_l158_108_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_108_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_108_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_108;
  wire       [6:0]    _zz_when_ArraySlice_l159_108_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_108_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_108_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_108_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_108_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_108_6;
  wire       [7:0]    _zz__zz_realValue_0_108;
  wire       [7:0]    _zz__zz_realValue_0_108_1;
  wire       [7:0]    _zz_realValue_0_108_1;
  wire       [7:0]    _zz_realValue_0_108_2;
  wire       [7:0]    _zz_realValue_0_108_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_108;
  wire       [6:0]    _zz_when_ArraySlice_l166_108_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_108_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_108_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_108_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_108_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_108_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_108_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_109;
  wire       [7:0]    _zz_when_ArraySlice_l158_109_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_109_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_109_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_109;
  wire       [5:0]    _zz_when_ArraySlice_l159_109_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_109_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_109_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_109_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_109_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_109_6;
  wire       [7:0]    _zz__zz_realValue_0_109;
  wire       [7:0]    _zz__zz_realValue_0_109_1;
  wire       [7:0]    _zz_realValue_0_109_1;
  wire       [7:0]    _zz_realValue_0_109_2;
  wire       [7:0]    _zz_realValue_0_109_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_109;
  wire       [5:0]    _zz_when_ArraySlice_l166_109_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_109_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_109_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_109_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_109_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_109_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_109_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_110;
  wire       [7:0]    _zz_when_ArraySlice_l158_110_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_110_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_110_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_110;
  wire       [5:0]    _zz_when_ArraySlice_l159_110_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_110_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_110_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_110_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_110_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_110_6;
  wire       [7:0]    _zz__zz_realValue_0_110;
  wire       [7:0]    _zz__zz_realValue_0_110_1;
  wire       [7:0]    _zz_realValue_0_110_1;
  wire       [7:0]    _zz_realValue_0_110_2;
  wire       [7:0]    _zz_realValue_0_110_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_110;
  wire       [5:0]    _zz_when_ArraySlice_l166_110_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_110_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_110_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_110_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_110_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_110_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_110_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_111;
  wire       [7:0]    _zz_when_ArraySlice_l158_111_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_111_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_111_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_111;
  wire       [4:0]    _zz_when_ArraySlice_l159_111_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_111_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_111_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_111_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_111_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_111_6;
  wire       [7:0]    _zz__zz_realValue_0_111;
  wire       [7:0]    _zz__zz_realValue_0_111_1;
  wire       [7:0]    _zz_realValue_0_111_1;
  wire       [7:0]    _zz_realValue_0_111_2;
  wire       [7:0]    _zz_realValue_0_111_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_111;
  wire       [4:0]    _zz_when_ArraySlice_l166_111_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_111_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_111_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_111_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_111_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_111_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_111_7;
  wire                _zz_when_ArraySlice_l400_4_1;
  wire                _zz_when_ArraySlice_l400_4_2;
  wire                _zz_when_ArraySlice_l400_4_3;
  wire                _zz_when_ArraySlice_l400_4_4;
  wire                _zz_when_ArraySlice_l400_4_5;
  wire                _zz_when_ArraySlice_l400_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_4_7;
  wire       [6:0]    _zz_when_ArraySlice_l403_4_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l406_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l406_4_5;
  wire       [7:0]    _zz_selectReadFifo_4_6;
  wire       [7:0]    _zz_selectReadFifo_4_7;
  wire       [6:0]    _zz_selectReadFifo_4_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_4;
  wire       [12:0]   _zz_when_ArraySlice_l413_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l417_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l417_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l417_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l418_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l418_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l418_4_5;
  wire       [7:0]    _zz__zz_realValue1_0_13;
  wire       [7:0]    _zz__zz_realValue1_0_13_1;
  wire       [7:0]    _zz_realValue1_0_13_1;
  wire       [7:0]    _zz_realValue1_0_13_2;
  wire       [7:0]    _zz_realValue1_0_13_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_4;
  wire       [6:0]    _zz_when_ArraySlice_l420_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_9;
  wire       [7:0]    _zz_selectReadFifo_4_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_112;
  wire       [7:0]    _zz_when_ArraySlice_l158_112_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_112_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_112_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_112;
  wire       [7:0]    _zz_when_ArraySlice_l159_112_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_112_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_112_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_112_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_112_5;
  wire       [7:0]    _zz__zz_realValue_0_112;
  wire       [7:0]    _zz__zz_realValue_0_112_1;
  wire       [7:0]    _zz_realValue_0_112_1;
  wire       [7:0]    _zz_realValue_0_112_2;
  wire       [7:0]    _zz_realValue_0_112_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_112;
  wire       [7:0]    _zz_when_ArraySlice_l166_112_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_112_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_112_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_112_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_112_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_112_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_113;
  wire       [7:0]    _zz_when_ArraySlice_l158_113_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_113_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_113_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_113;
  wire       [6:0]    _zz_when_ArraySlice_l159_113_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_113_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_113_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_113_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_113_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_113_6;
  wire       [7:0]    _zz__zz_realValue_0_113;
  wire       [7:0]    _zz__zz_realValue_0_113_1;
  wire       [7:0]    _zz_realValue_0_113_1;
  wire       [7:0]    _zz_realValue_0_113_2;
  wire       [7:0]    _zz_realValue_0_113_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_113;
  wire       [6:0]    _zz_when_ArraySlice_l166_113_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_113_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_113_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_113_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_113_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_113_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_113_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_114;
  wire       [7:0]    _zz_when_ArraySlice_l158_114_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_114_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_114_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_114;
  wire       [6:0]    _zz_when_ArraySlice_l159_114_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_114_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_114_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_114_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_114_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_114_6;
  wire       [7:0]    _zz__zz_realValue_0_114;
  wire       [7:0]    _zz__zz_realValue_0_114_1;
  wire       [7:0]    _zz_realValue_0_114_1;
  wire       [7:0]    _zz_realValue_0_114_2;
  wire       [7:0]    _zz_realValue_0_114_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_114;
  wire       [6:0]    _zz_when_ArraySlice_l166_114_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_114_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_114_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_114_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_114_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_114_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_114_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_115;
  wire       [7:0]    _zz_when_ArraySlice_l158_115_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_115_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_115_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_115;
  wire       [6:0]    _zz_when_ArraySlice_l159_115_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_115_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_115_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_115_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_115_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_115_6;
  wire       [7:0]    _zz__zz_realValue_0_115;
  wire       [7:0]    _zz__zz_realValue_0_115_1;
  wire       [7:0]    _zz_realValue_0_115_1;
  wire       [7:0]    _zz_realValue_0_115_2;
  wire       [7:0]    _zz_realValue_0_115_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_115;
  wire       [6:0]    _zz_when_ArraySlice_l166_115_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_115_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_115_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_115_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_115_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_115_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_115_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_116;
  wire       [7:0]    _zz_when_ArraySlice_l158_116_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_116_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_116_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_116;
  wire       [6:0]    _zz_when_ArraySlice_l159_116_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_116_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_116_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_116_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_116_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_116_6;
  wire       [7:0]    _zz__zz_realValue_0_116;
  wire       [7:0]    _zz__zz_realValue_0_116_1;
  wire       [7:0]    _zz_realValue_0_116_1;
  wire       [7:0]    _zz_realValue_0_116_2;
  wire       [7:0]    _zz_realValue_0_116_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_116;
  wire       [6:0]    _zz_when_ArraySlice_l166_116_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_116_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_116_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_116_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_116_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_116_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_116_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_117;
  wire       [7:0]    _zz_when_ArraySlice_l158_117_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_117_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_117_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_117;
  wire       [5:0]    _zz_when_ArraySlice_l159_117_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_117_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_117_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_117_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_117_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_117_6;
  wire       [7:0]    _zz__zz_realValue_0_117;
  wire       [7:0]    _zz__zz_realValue_0_117_1;
  wire       [7:0]    _zz_realValue_0_117_1;
  wire       [7:0]    _zz_realValue_0_117_2;
  wire       [7:0]    _zz_realValue_0_117_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_117;
  wire       [5:0]    _zz_when_ArraySlice_l166_117_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_117_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_117_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_117_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_117_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_117_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_117_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_118;
  wire       [7:0]    _zz_when_ArraySlice_l158_118_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_118_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_118_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_118;
  wire       [5:0]    _zz_when_ArraySlice_l159_118_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_118_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_118_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_118_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_118_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_118_6;
  wire       [7:0]    _zz__zz_realValue_0_118;
  wire       [7:0]    _zz__zz_realValue_0_118_1;
  wire       [7:0]    _zz_realValue_0_118_1;
  wire       [7:0]    _zz_realValue_0_118_2;
  wire       [7:0]    _zz_realValue_0_118_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_118;
  wire       [5:0]    _zz_when_ArraySlice_l166_118_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_118_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_118_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_118_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_118_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_118_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_118_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_119;
  wire       [7:0]    _zz_when_ArraySlice_l158_119_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_119_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_119_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_119;
  wire       [4:0]    _zz_when_ArraySlice_l159_119_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_119_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_119_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_119_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_119_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_119_6;
  wire       [7:0]    _zz__zz_realValue_0_119;
  wire       [7:0]    _zz__zz_realValue_0_119_1;
  wire       [7:0]    _zz_realValue_0_119_1;
  wire       [7:0]    _zz_realValue_0_119_2;
  wire       [7:0]    _zz_realValue_0_119_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_119;
  wire       [4:0]    _zz_when_ArraySlice_l166_119_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_119_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_119_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_119_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_119_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_119_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_119_7;
  wire                _zz_when_ArraySlice_l425_4_1;
  wire                _zz_when_ArraySlice_l425_4_2;
  wire                _zz_when_ArraySlice_l425_4_3;
  wire                _zz_when_ArraySlice_l425_4_4;
  wire                _zz_when_ArraySlice_l425_4_5;
  wire                _zz_when_ArraySlice_l425_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_4_7;
  wire       [6:0]    _zz_when_ArraySlice_l428_4_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l431_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l431_4_5;
  wire       [7:0]    _zz_selectReadFifo_4_11;
  wire       [7:0]    _zz_selectReadFifo_4_12;
  wire       [6:0]    _zz_selectReadFifo_4_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_4;
  wire       [12:0]   _zz_when_ArraySlice_l438_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_4;
  wire       [7:0]    _zz_when_ArraySlice_l449_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_4_2;
  wire       [7:0]    _zz__zz_realValue1_0_14;
  wire       [7:0]    _zz__zz_realValue1_0_14_1;
  wire       [7:0]    _zz_realValue1_0_14_1;
  wire       [7:0]    _zz_realValue1_0_14_2;
  wire       [7:0]    _zz_realValue1_0_14_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_4;
  wire       [6:0]    _zz_when_ArraySlice_l450_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_14;
  wire       [7:0]    _zz_selectReadFifo_4_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_120;
  wire       [7:0]    _zz_when_ArraySlice_l158_120_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_120_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_120_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_120;
  wire       [7:0]    _zz_when_ArraySlice_l159_120_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_120_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_120_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_120_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_120_5;
  wire       [7:0]    _zz__zz_realValue_0_120;
  wire       [7:0]    _zz__zz_realValue_0_120_1;
  wire       [7:0]    _zz_realValue_0_120_1;
  wire       [7:0]    _zz_realValue_0_120_2;
  wire       [7:0]    _zz_realValue_0_120_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_120;
  wire       [7:0]    _zz_when_ArraySlice_l166_120_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_120_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_120_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_120_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_120_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_120_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_121;
  wire       [7:0]    _zz_when_ArraySlice_l158_121_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_121_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_121_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_121;
  wire       [6:0]    _zz_when_ArraySlice_l159_121_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_121_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_121_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_121_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_121_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_121_6;
  wire       [7:0]    _zz__zz_realValue_0_121;
  wire       [7:0]    _zz__zz_realValue_0_121_1;
  wire       [7:0]    _zz_realValue_0_121_1;
  wire       [7:0]    _zz_realValue_0_121_2;
  wire       [7:0]    _zz_realValue_0_121_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_121;
  wire       [6:0]    _zz_when_ArraySlice_l166_121_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_121_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_121_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_121_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_121_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_121_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_121_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_122;
  wire       [7:0]    _zz_when_ArraySlice_l158_122_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_122_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_122_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_122;
  wire       [6:0]    _zz_when_ArraySlice_l159_122_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_122_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_122_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_122_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_122_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_122_6;
  wire       [7:0]    _zz__zz_realValue_0_122;
  wire       [7:0]    _zz__zz_realValue_0_122_1;
  wire       [7:0]    _zz_realValue_0_122_1;
  wire       [7:0]    _zz_realValue_0_122_2;
  wire       [7:0]    _zz_realValue_0_122_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_122;
  wire       [6:0]    _zz_when_ArraySlice_l166_122_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_122_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_122_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_122_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_122_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_122_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_122_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_123;
  wire       [7:0]    _zz_when_ArraySlice_l158_123_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_123_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_123_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_123;
  wire       [6:0]    _zz_when_ArraySlice_l159_123_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_123_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_123_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_123_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_123_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_123_6;
  wire       [7:0]    _zz__zz_realValue_0_123;
  wire       [7:0]    _zz__zz_realValue_0_123_1;
  wire       [7:0]    _zz_realValue_0_123_1;
  wire       [7:0]    _zz_realValue_0_123_2;
  wire       [7:0]    _zz_realValue_0_123_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_123;
  wire       [6:0]    _zz_when_ArraySlice_l166_123_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_123_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_123_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_123_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_123_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_123_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_123_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_124;
  wire       [7:0]    _zz_when_ArraySlice_l158_124_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_124_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_124_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_124;
  wire       [6:0]    _zz_when_ArraySlice_l159_124_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_124_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_124_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_124_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_124_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_124_6;
  wire       [7:0]    _zz__zz_realValue_0_124;
  wire       [7:0]    _zz__zz_realValue_0_124_1;
  wire       [7:0]    _zz_realValue_0_124_1;
  wire       [7:0]    _zz_realValue_0_124_2;
  wire       [7:0]    _zz_realValue_0_124_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_124;
  wire       [6:0]    _zz_when_ArraySlice_l166_124_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_124_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_124_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_124_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_124_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_124_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_124_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_125;
  wire       [7:0]    _zz_when_ArraySlice_l158_125_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_125_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_125_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_125;
  wire       [5:0]    _zz_when_ArraySlice_l159_125_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_125_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_125_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_125_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_125_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_125_6;
  wire       [7:0]    _zz__zz_realValue_0_125;
  wire       [7:0]    _zz__zz_realValue_0_125_1;
  wire       [7:0]    _zz_realValue_0_125_1;
  wire       [7:0]    _zz_realValue_0_125_2;
  wire       [7:0]    _zz_realValue_0_125_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_125;
  wire       [5:0]    _zz_when_ArraySlice_l166_125_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_125_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_125_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_125_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_125_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_125_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_125_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_126;
  wire       [7:0]    _zz_when_ArraySlice_l158_126_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_126_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_126_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_126;
  wire       [5:0]    _zz_when_ArraySlice_l159_126_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_126_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_126_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_126_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_126_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_126_6;
  wire       [7:0]    _zz__zz_realValue_0_126;
  wire       [7:0]    _zz__zz_realValue_0_126_1;
  wire       [7:0]    _zz_realValue_0_126_1;
  wire       [7:0]    _zz_realValue_0_126_2;
  wire       [7:0]    _zz_realValue_0_126_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_126;
  wire       [5:0]    _zz_when_ArraySlice_l166_126_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_126_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_126_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_126_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_126_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_126_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_126_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_127;
  wire       [7:0]    _zz_when_ArraySlice_l158_127_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_127_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_127_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_127;
  wire       [4:0]    _zz_when_ArraySlice_l159_127_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_127_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_127_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_127_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_127_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_127_6;
  wire       [7:0]    _zz__zz_realValue_0_127;
  wire       [7:0]    _zz__zz_realValue_0_127_1;
  wire       [7:0]    _zz_realValue_0_127_1;
  wire       [7:0]    _zz_realValue_0_127_2;
  wire       [7:0]    _zz_realValue_0_127_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_127;
  wire       [4:0]    _zz_when_ArraySlice_l166_127_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_127_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_127_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_127_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_127_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_127_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_127_7;
  wire                _zz_when_ArraySlice_l457_4_1;
  wire                _zz_when_ArraySlice_l457_4_2;
  wire                _zz_when_ArraySlice_l457_4_3;
  wire                _zz_when_ArraySlice_l457_4_4;
  wire                _zz_when_ArraySlice_l457_4_5;
  wire                _zz_when_ArraySlice_l457_4_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_4;
  wire       [12:0]   _zz_when_ArraySlice_l461_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_4;
  wire       [7:0]    _zz_when_ArraySlice_l447_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_4_2;
  wire       [6:0]    _zz_when_ArraySlice_l447_4_3;
  wire       [12:0]   _zz_when_ArraySlice_l468_4;
  wire       [7:0]    _zz_when_ArraySlice_l468_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_5;
  wire       [7:0]    _zz_when_ArraySlice_l376_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l376_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l377_5;
  wire       [6:0]    _zz_when_ArraySlice_l377_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l377_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l377_5_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_5_valid;
  wire       [6:0]    _zz__zz_outputStreamArrayData_5_valid_1;
  wire       [6:0]    _zz__zz_8;
  reg                 _zz_outputStreamArrayData_5_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_5_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_5_payload;
  wire       [6:0]    _zz_outputStreamArrayData_5_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_5;
  wire       [6:0]    _zz_when_ArraySlice_l383_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l383_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l383_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l384_5;
  wire       [7:0]    _zz_when_ArraySlice_l384_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_5_2;
  wire       [7:0]    _zz_selectReadFifo_5;
  wire       [7:0]    _zz_selectReadFifo_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_5;
  wire       [12:0]   _zz_when_ArraySlice_l387_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_5;
  wire       [6:0]    _zz_when_ArraySlice_l392_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l392_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l393_5;
  wire       [7:0]    _zz_when_ArraySlice_l393_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_5_2;
  wire       [7:0]    _zz__zz_realValue1_0_15;
  wire       [7:0]    _zz__zz_realValue1_0_15_1;
  wire       [7:0]    _zz_realValue1_0_15_1;
  wire       [7:0]    _zz_realValue1_0_15_2;
  wire       [7:0]    _zz_realValue1_0_15_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_5;
  wire       [6:0]    _zz_when_ArraySlice_l395_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_3;
  wire       [7:0]    _zz_selectReadFifo_5_4;
  wire       [0:0]    _zz_selectReadFifo_5_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_128;
  wire       [7:0]    _zz_when_ArraySlice_l158_128_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_128_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_128_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_128;
  wire       [7:0]    _zz_when_ArraySlice_l159_128_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_128_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_128_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_128_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_128_5;
  wire       [7:0]    _zz__zz_realValue_0_128;
  wire       [7:0]    _zz__zz_realValue_0_128_1;
  wire       [7:0]    _zz_realValue_0_128_1;
  wire       [7:0]    _zz_realValue_0_128_2;
  wire       [7:0]    _zz_realValue_0_128_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_128;
  wire       [7:0]    _zz_when_ArraySlice_l166_128_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_128_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_128_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_128_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_128_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_128_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_129;
  wire       [7:0]    _zz_when_ArraySlice_l158_129_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_129_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_129_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_129;
  wire       [6:0]    _zz_when_ArraySlice_l159_129_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_129_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_129_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_129_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_129_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_129_6;
  wire       [7:0]    _zz__zz_realValue_0_129;
  wire       [7:0]    _zz__zz_realValue_0_129_1;
  wire       [7:0]    _zz_realValue_0_129_1;
  wire       [7:0]    _zz_realValue_0_129_2;
  wire       [7:0]    _zz_realValue_0_129_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_129;
  wire       [6:0]    _zz_when_ArraySlice_l166_129_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_129_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_129_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_129_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_129_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_129_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_129_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_130;
  wire       [7:0]    _zz_when_ArraySlice_l158_130_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_130_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_130_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_130;
  wire       [6:0]    _zz_when_ArraySlice_l159_130_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_130_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_130_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_130_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_130_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_130_6;
  wire       [7:0]    _zz__zz_realValue_0_130;
  wire       [7:0]    _zz__zz_realValue_0_130_1;
  wire       [7:0]    _zz_realValue_0_130_1;
  wire       [7:0]    _zz_realValue_0_130_2;
  wire       [7:0]    _zz_realValue_0_130_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_130;
  wire       [6:0]    _zz_when_ArraySlice_l166_130_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_130_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_130_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_130_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_130_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_130_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_130_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_131;
  wire       [7:0]    _zz_when_ArraySlice_l158_131_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_131_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_131_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_131;
  wire       [6:0]    _zz_when_ArraySlice_l159_131_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_131_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_131_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_131_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_131_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_131_6;
  wire       [7:0]    _zz__zz_realValue_0_131;
  wire       [7:0]    _zz__zz_realValue_0_131_1;
  wire       [7:0]    _zz_realValue_0_131_1;
  wire       [7:0]    _zz_realValue_0_131_2;
  wire       [7:0]    _zz_realValue_0_131_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_131;
  wire       [6:0]    _zz_when_ArraySlice_l166_131_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_131_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_131_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_131_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_131_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_131_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_131_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_132;
  wire       [7:0]    _zz_when_ArraySlice_l158_132_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_132_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_132_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_132;
  wire       [6:0]    _zz_when_ArraySlice_l159_132_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_132_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_132_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_132_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_132_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_132_6;
  wire       [7:0]    _zz__zz_realValue_0_132;
  wire       [7:0]    _zz__zz_realValue_0_132_1;
  wire       [7:0]    _zz_realValue_0_132_1;
  wire       [7:0]    _zz_realValue_0_132_2;
  wire       [7:0]    _zz_realValue_0_132_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_132;
  wire       [6:0]    _zz_when_ArraySlice_l166_132_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_132_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_132_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_132_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_132_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_132_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_132_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_133;
  wire       [7:0]    _zz_when_ArraySlice_l158_133_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_133_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_133_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_133;
  wire       [5:0]    _zz_when_ArraySlice_l159_133_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_133_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_133_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_133_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_133_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_133_6;
  wire       [7:0]    _zz__zz_realValue_0_133;
  wire       [7:0]    _zz__zz_realValue_0_133_1;
  wire       [7:0]    _zz_realValue_0_133_1;
  wire       [7:0]    _zz_realValue_0_133_2;
  wire       [7:0]    _zz_realValue_0_133_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_133;
  wire       [5:0]    _zz_when_ArraySlice_l166_133_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_133_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_133_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_133_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_133_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_133_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_133_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_134;
  wire       [7:0]    _zz_when_ArraySlice_l158_134_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_134_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_134_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_134;
  wire       [5:0]    _zz_when_ArraySlice_l159_134_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_134_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_134_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_134_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_134_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_134_6;
  wire       [7:0]    _zz__zz_realValue_0_134;
  wire       [7:0]    _zz__zz_realValue_0_134_1;
  wire       [7:0]    _zz_realValue_0_134_1;
  wire       [7:0]    _zz_realValue_0_134_2;
  wire       [7:0]    _zz_realValue_0_134_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_134;
  wire       [5:0]    _zz_when_ArraySlice_l166_134_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_134_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_134_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_134_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_134_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_134_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_134_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_135;
  wire       [7:0]    _zz_when_ArraySlice_l158_135_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_135_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_135_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_135;
  wire       [4:0]    _zz_when_ArraySlice_l159_135_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_135_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_135_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_135_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_135_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_135_6;
  wire       [7:0]    _zz__zz_realValue_0_135;
  wire       [7:0]    _zz__zz_realValue_0_135_1;
  wire       [7:0]    _zz_realValue_0_135_1;
  wire       [7:0]    _zz_realValue_0_135_2;
  wire       [7:0]    _zz_realValue_0_135_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_135;
  wire       [4:0]    _zz_when_ArraySlice_l166_135_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_135_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_135_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_135_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_135_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_135_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_135_7;
  wire                _zz_when_ArraySlice_l400_5_1;
  wire                _zz_when_ArraySlice_l400_5_2;
  wire                _zz_when_ArraySlice_l400_5_3;
  wire                _zz_when_ArraySlice_l400_5_4;
  wire                _zz_when_ArraySlice_l400_5_5;
  wire                _zz_when_ArraySlice_l400_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_5_7;
  wire       [6:0]    _zz_when_ArraySlice_l403_5_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_5;
  wire       [7:0]    _zz_when_ArraySlice_l406_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l406_5_4;
  wire       [7:0]    _zz_selectReadFifo_5_6;
  wire       [7:0]    _zz_selectReadFifo_5_7;
  wire       [6:0]    _zz_selectReadFifo_5_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_5;
  wire       [12:0]   _zz_when_ArraySlice_l413_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_5;
  wire       [6:0]    _zz_when_ArraySlice_l417_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l417_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l417_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l418_5;
  wire       [7:0]    _zz_when_ArraySlice_l418_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l418_5_4;
  wire       [7:0]    _zz__zz_realValue1_0_16;
  wire       [7:0]    _zz__zz_realValue1_0_16_1;
  wire       [7:0]    _zz_realValue1_0_16_1;
  wire       [7:0]    _zz_realValue1_0_16_2;
  wire       [7:0]    _zz_realValue1_0_16_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_5;
  wire       [6:0]    _zz_when_ArraySlice_l420_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_9;
  wire       [7:0]    _zz_selectReadFifo_5_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_136;
  wire       [7:0]    _zz_when_ArraySlice_l158_136_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_136_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_136_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_136;
  wire       [7:0]    _zz_when_ArraySlice_l159_136_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_136_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_136_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_136_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_136_5;
  wire       [7:0]    _zz__zz_realValue_0_136;
  wire       [7:0]    _zz__zz_realValue_0_136_1;
  wire       [7:0]    _zz_realValue_0_136_1;
  wire       [7:0]    _zz_realValue_0_136_2;
  wire       [7:0]    _zz_realValue_0_136_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_136;
  wire       [7:0]    _zz_when_ArraySlice_l166_136_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_136_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_136_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_136_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_136_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_136_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_137;
  wire       [7:0]    _zz_when_ArraySlice_l158_137_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_137_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_137_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_137;
  wire       [6:0]    _zz_when_ArraySlice_l159_137_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_137_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_137_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_137_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_137_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_137_6;
  wire       [7:0]    _zz__zz_realValue_0_137;
  wire       [7:0]    _zz__zz_realValue_0_137_1;
  wire       [7:0]    _zz_realValue_0_137_1;
  wire       [7:0]    _zz_realValue_0_137_2;
  wire       [7:0]    _zz_realValue_0_137_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_137;
  wire       [6:0]    _zz_when_ArraySlice_l166_137_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_137_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_137_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_137_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_137_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_137_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_137_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_138;
  wire       [7:0]    _zz_when_ArraySlice_l158_138_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_138_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_138_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_138;
  wire       [6:0]    _zz_when_ArraySlice_l159_138_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_138_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_138_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_138_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_138_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_138_6;
  wire       [7:0]    _zz__zz_realValue_0_138;
  wire       [7:0]    _zz__zz_realValue_0_138_1;
  wire       [7:0]    _zz_realValue_0_138_1;
  wire       [7:0]    _zz_realValue_0_138_2;
  wire       [7:0]    _zz_realValue_0_138_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_138;
  wire       [6:0]    _zz_when_ArraySlice_l166_138_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_138_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_138_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_138_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_138_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_138_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_138_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_139;
  wire       [7:0]    _zz_when_ArraySlice_l158_139_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_139_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_139_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_139;
  wire       [6:0]    _zz_when_ArraySlice_l159_139_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_139_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_139_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_139_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_139_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_139_6;
  wire       [7:0]    _zz__zz_realValue_0_139;
  wire       [7:0]    _zz__zz_realValue_0_139_1;
  wire       [7:0]    _zz_realValue_0_139_1;
  wire       [7:0]    _zz_realValue_0_139_2;
  wire       [7:0]    _zz_realValue_0_139_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_139;
  wire       [6:0]    _zz_when_ArraySlice_l166_139_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_139_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_139_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_139_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_139_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_139_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_139_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_140;
  wire       [7:0]    _zz_when_ArraySlice_l158_140_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_140_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_140_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_140;
  wire       [6:0]    _zz_when_ArraySlice_l159_140_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_140_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_140_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_140_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_140_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_140_6;
  wire       [7:0]    _zz__zz_realValue_0_140;
  wire       [7:0]    _zz__zz_realValue_0_140_1;
  wire       [7:0]    _zz_realValue_0_140_1;
  wire       [7:0]    _zz_realValue_0_140_2;
  wire       [7:0]    _zz_realValue_0_140_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_140;
  wire       [6:0]    _zz_when_ArraySlice_l166_140_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_140_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_140_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_140_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_140_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_140_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_140_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_141;
  wire       [7:0]    _zz_when_ArraySlice_l158_141_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_141_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_141_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_141;
  wire       [5:0]    _zz_when_ArraySlice_l159_141_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_141_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_141_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_141_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_141_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_141_6;
  wire       [7:0]    _zz__zz_realValue_0_141;
  wire       [7:0]    _zz__zz_realValue_0_141_1;
  wire       [7:0]    _zz_realValue_0_141_1;
  wire       [7:0]    _zz_realValue_0_141_2;
  wire       [7:0]    _zz_realValue_0_141_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_141;
  wire       [5:0]    _zz_when_ArraySlice_l166_141_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_141_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_141_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_141_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_141_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_141_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_141_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_142;
  wire       [7:0]    _zz_when_ArraySlice_l158_142_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_142_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_142_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_142;
  wire       [5:0]    _zz_when_ArraySlice_l159_142_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_142_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_142_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_142_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_142_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_142_6;
  wire       [7:0]    _zz__zz_realValue_0_142;
  wire       [7:0]    _zz__zz_realValue_0_142_1;
  wire       [7:0]    _zz_realValue_0_142_1;
  wire       [7:0]    _zz_realValue_0_142_2;
  wire       [7:0]    _zz_realValue_0_142_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_142;
  wire       [5:0]    _zz_when_ArraySlice_l166_142_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_142_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_142_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_142_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_142_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_142_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_142_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_143;
  wire       [7:0]    _zz_when_ArraySlice_l158_143_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_143_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_143_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_143;
  wire       [4:0]    _zz_when_ArraySlice_l159_143_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_143_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_143_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_143_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_143_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_143_6;
  wire       [7:0]    _zz__zz_realValue_0_143;
  wire       [7:0]    _zz__zz_realValue_0_143_1;
  wire       [7:0]    _zz_realValue_0_143_1;
  wire       [7:0]    _zz_realValue_0_143_2;
  wire       [7:0]    _zz_realValue_0_143_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_143;
  wire       [4:0]    _zz_when_ArraySlice_l166_143_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_143_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_143_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_143_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_143_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_143_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_143_7;
  wire                _zz_when_ArraySlice_l425_5_1;
  wire                _zz_when_ArraySlice_l425_5_2;
  wire                _zz_when_ArraySlice_l425_5_3;
  wire                _zz_when_ArraySlice_l425_5_4;
  wire                _zz_when_ArraySlice_l425_5_5;
  wire                _zz_when_ArraySlice_l425_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_5_7;
  wire       [6:0]    _zz_when_ArraySlice_l428_5_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_5;
  wire       [7:0]    _zz_when_ArraySlice_l431_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l431_5_4;
  wire       [7:0]    _zz_selectReadFifo_5_11;
  wire       [7:0]    _zz_selectReadFifo_5_12;
  wire       [6:0]    _zz_selectReadFifo_5_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_5;
  wire       [12:0]   _zz_when_ArraySlice_l438_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_5;
  wire       [7:0]    _zz_when_ArraySlice_l449_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_5_2;
  wire       [7:0]    _zz__zz_realValue1_0_17;
  wire       [7:0]    _zz__zz_realValue1_0_17_1;
  wire       [7:0]    _zz_realValue1_0_17_1;
  wire       [7:0]    _zz_realValue1_0_17_2;
  wire       [7:0]    _zz_realValue1_0_17_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_5;
  wire       [6:0]    _zz_when_ArraySlice_l450_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_14;
  wire       [7:0]    _zz_selectReadFifo_5_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_144;
  wire       [7:0]    _zz_when_ArraySlice_l158_144_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_144_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_144_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_144;
  wire       [7:0]    _zz_when_ArraySlice_l159_144_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_144_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_144_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_144_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_144_5;
  wire       [7:0]    _zz__zz_realValue_0_144;
  wire       [7:0]    _zz__zz_realValue_0_144_1;
  wire       [7:0]    _zz_realValue_0_144_1;
  wire       [7:0]    _zz_realValue_0_144_2;
  wire       [7:0]    _zz_realValue_0_144_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_144;
  wire       [7:0]    _zz_when_ArraySlice_l166_144_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_144_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_144_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_144_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_144_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_144_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_145;
  wire       [7:0]    _zz_when_ArraySlice_l158_145_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_145_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_145_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_145;
  wire       [6:0]    _zz_when_ArraySlice_l159_145_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_145_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_145_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_145_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_145_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_145_6;
  wire       [7:0]    _zz__zz_realValue_0_145;
  wire       [7:0]    _zz__zz_realValue_0_145_1;
  wire       [7:0]    _zz_realValue_0_145_1;
  wire       [7:0]    _zz_realValue_0_145_2;
  wire       [7:0]    _zz_realValue_0_145_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_145;
  wire       [6:0]    _zz_when_ArraySlice_l166_145_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_145_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_145_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_145_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_145_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_145_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_145_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_146;
  wire       [7:0]    _zz_when_ArraySlice_l158_146_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_146_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_146_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_146;
  wire       [6:0]    _zz_when_ArraySlice_l159_146_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_146_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_146_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_146_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_146_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_146_6;
  wire       [7:0]    _zz__zz_realValue_0_146;
  wire       [7:0]    _zz__zz_realValue_0_146_1;
  wire       [7:0]    _zz_realValue_0_146_1;
  wire       [7:0]    _zz_realValue_0_146_2;
  wire       [7:0]    _zz_realValue_0_146_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_146;
  wire       [6:0]    _zz_when_ArraySlice_l166_146_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_146_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_146_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_146_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_146_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_146_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_146_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_147;
  wire       [7:0]    _zz_when_ArraySlice_l158_147_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_147_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_147_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_147;
  wire       [6:0]    _zz_when_ArraySlice_l159_147_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_147_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_147_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_147_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_147_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_147_6;
  wire       [7:0]    _zz__zz_realValue_0_147;
  wire       [7:0]    _zz__zz_realValue_0_147_1;
  wire       [7:0]    _zz_realValue_0_147_1;
  wire       [7:0]    _zz_realValue_0_147_2;
  wire       [7:0]    _zz_realValue_0_147_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_147;
  wire       [6:0]    _zz_when_ArraySlice_l166_147_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_147_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_147_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_147_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_147_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_147_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_147_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_148;
  wire       [7:0]    _zz_when_ArraySlice_l158_148_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_148_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_148_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_148;
  wire       [6:0]    _zz_when_ArraySlice_l159_148_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_148_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_148_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_148_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_148_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_148_6;
  wire       [7:0]    _zz__zz_realValue_0_148;
  wire       [7:0]    _zz__zz_realValue_0_148_1;
  wire       [7:0]    _zz_realValue_0_148_1;
  wire       [7:0]    _zz_realValue_0_148_2;
  wire       [7:0]    _zz_realValue_0_148_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_148;
  wire       [6:0]    _zz_when_ArraySlice_l166_148_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_148_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_148_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_148_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_148_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_148_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_148_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_149;
  wire       [7:0]    _zz_when_ArraySlice_l158_149_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_149_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_149_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_149;
  wire       [5:0]    _zz_when_ArraySlice_l159_149_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_149_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_149_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_149_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_149_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_149_6;
  wire       [7:0]    _zz__zz_realValue_0_149;
  wire       [7:0]    _zz__zz_realValue_0_149_1;
  wire       [7:0]    _zz_realValue_0_149_1;
  wire       [7:0]    _zz_realValue_0_149_2;
  wire       [7:0]    _zz_realValue_0_149_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_149;
  wire       [5:0]    _zz_when_ArraySlice_l166_149_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_149_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_149_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_149_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_149_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_149_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_149_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_150;
  wire       [7:0]    _zz_when_ArraySlice_l158_150_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_150_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_150_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_150;
  wire       [5:0]    _zz_when_ArraySlice_l159_150_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_150_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_150_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_150_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_150_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_150_6;
  wire       [7:0]    _zz__zz_realValue_0_150;
  wire       [7:0]    _zz__zz_realValue_0_150_1;
  wire       [7:0]    _zz_realValue_0_150_1;
  wire       [7:0]    _zz_realValue_0_150_2;
  wire       [7:0]    _zz_realValue_0_150_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_150;
  wire       [5:0]    _zz_when_ArraySlice_l166_150_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_150_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_150_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_150_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_150_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_150_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_150_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_151;
  wire       [7:0]    _zz_when_ArraySlice_l158_151_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_151_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_151_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_151;
  wire       [4:0]    _zz_when_ArraySlice_l159_151_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_151_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_151_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_151_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_151_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_151_6;
  wire       [7:0]    _zz__zz_realValue_0_151;
  wire       [7:0]    _zz__zz_realValue_0_151_1;
  wire       [7:0]    _zz_realValue_0_151_1;
  wire       [7:0]    _zz_realValue_0_151_2;
  wire       [7:0]    _zz_realValue_0_151_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_151;
  wire       [4:0]    _zz_when_ArraySlice_l166_151_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_151_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_151_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_151_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_151_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_151_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_151_7;
  wire                _zz_when_ArraySlice_l457_5_1;
  wire                _zz_when_ArraySlice_l457_5_2;
  wire                _zz_when_ArraySlice_l457_5_3;
  wire                _zz_when_ArraySlice_l457_5_4;
  wire                _zz_when_ArraySlice_l457_5_5;
  wire                _zz_when_ArraySlice_l457_5_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_5;
  wire       [12:0]   _zz_when_ArraySlice_l461_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_5;
  wire       [7:0]    _zz_when_ArraySlice_l447_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_5_2;
  wire       [6:0]    _zz_when_ArraySlice_l447_5_3;
  wire       [12:0]   _zz_when_ArraySlice_l468_5;
  wire       [7:0]    _zz_when_ArraySlice_l468_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_6;
  wire       [7:0]    _zz_when_ArraySlice_l376_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l376_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l377_6;
  wire       [6:0]    _zz_when_ArraySlice_l377_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l377_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l377_6_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_6_valid;
  wire       [6:0]    _zz__zz_outputStreamArrayData_6_valid_1;
  wire       [6:0]    _zz__zz_9;
  reg                 _zz_outputStreamArrayData_6_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_6_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_6_payload;
  wire       [6:0]    _zz_outputStreamArrayData_6_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_6;
  wire       [6:0]    _zz_when_ArraySlice_l383_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l383_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l383_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l384_6;
  wire       [7:0]    _zz_when_ArraySlice_l384_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_6_2;
  wire       [7:0]    _zz_selectReadFifo_6;
  wire       [7:0]    _zz_selectReadFifo_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_6;
  wire       [12:0]   _zz_when_ArraySlice_l387_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_6;
  wire       [6:0]    _zz_when_ArraySlice_l392_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l392_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l393_6;
  wire       [7:0]    _zz_when_ArraySlice_l393_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_6_2;
  wire       [7:0]    _zz__zz_realValue1_0_18;
  wire       [7:0]    _zz__zz_realValue1_0_18_1;
  wire       [7:0]    _zz_realValue1_0_18_1;
  wire       [7:0]    _zz_realValue1_0_18_2;
  wire       [7:0]    _zz_realValue1_0_18_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_6;
  wire       [6:0]    _zz_when_ArraySlice_l395_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_3;
  wire       [7:0]    _zz_selectReadFifo_6_4;
  wire       [0:0]    _zz_selectReadFifo_6_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_152;
  wire       [7:0]    _zz_when_ArraySlice_l158_152_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_152_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_152_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_152;
  wire       [7:0]    _zz_when_ArraySlice_l159_152_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_152_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_152_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_152_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_152_5;
  wire       [7:0]    _zz__zz_realValue_0_152;
  wire       [7:0]    _zz__zz_realValue_0_152_1;
  wire       [7:0]    _zz_realValue_0_152_1;
  wire       [7:0]    _zz_realValue_0_152_2;
  wire       [7:0]    _zz_realValue_0_152_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_152;
  wire       [7:0]    _zz_when_ArraySlice_l166_152_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_152_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_152_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_152_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_152_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_152_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_153;
  wire       [7:0]    _zz_when_ArraySlice_l158_153_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_153_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_153_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_153;
  wire       [6:0]    _zz_when_ArraySlice_l159_153_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_153_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_153_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_153_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_153_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_153_6;
  wire       [7:0]    _zz__zz_realValue_0_153;
  wire       [7:0]    _zz__zz_realValue_0_153_1;
  wire       [7:0]    _zz_realValue_0_153_1;
  wire       [7:0]    _zz_realValue_0_153_2;
  wire       [7:0]    _zz_realValue_0_153_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_153;
  wire       [6:0]    _zz_when_ArraySlice_l166_153_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_153_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_153_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_153_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_153_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_153_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_153_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_154;
  wire       [7:0]    _zz_when_ArraySlice_l158_154_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_154_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_154_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_154;
  wire       [6:0]    _zz_when_ArraySlice_l159_154_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_154_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_154_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_154_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_154_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_154_6;
  wire       [7:0]    _zz__zz_realValue_0_154;
  wire       [7:0]    _zz__zz_realValue_0_154_1;
  wire       [7:0]    _zz_realValue_0_154_1;
  wire       [7:0]    _zz_realValue_0_154_2;
  wire       [7:0]    _zz_realValue_0_154_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_154;
  wire       [6:0]    _zz_when_ArraySlice_l166_154_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_154_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_154_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_154_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_154_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_154_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_154_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_155;
  wire       [7:0]    _zz_when_ArraySlice_l158_155_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_155_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_155_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_155;
  wire       [6:0]    _zz_when_ArraySlice_l159_155_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_155_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_155_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_155_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_155_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_155_6;
  wire       [7:0]    _zz__zz_realValue_0_155;
  wire       [7:0]    _zz__zz_realValue_0_155_1;
  wire       [7:0]    _zz_realValue_0_155_1;
  wire       [7:0]    _zz_realValue_0_155_2;
  wire       [7:0]    _zz_realValue_0_155_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_155;
  wire       [6:0]    _zz_when_ArraySlice_l166_155_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_155_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_155_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_155_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_155_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_155_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_155_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_156;
  wire       [7:0]    _zz_when_ArraySlice_l158_156_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_156_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_156_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_156;
  wire       [6:0]    _zz_when_ArraySlice_l159_156_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_156_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_156_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_156_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_156_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_156_6;
  wire       [7:0]    _zz__zz_realValue_0_156;
  wire       [7:0]    _zz__zz_realValue_0_156_1;
  wire       [7:0]    _zz_realValue_0_156_1;
  wire       [7:0]    _zz_realValue_0_156_2;
  wire       [7:0]    _zz_realValue_0_156_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_156;
  wire       [6:0]    _zz_when_ArraySlice_l166_156_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_156_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_156_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_156_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_156_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_156_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_156_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_157;
  wire       [7:0]    _zz_when_ArraySlice_l158_157_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_157_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_157_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_157;
  wire       [5:0]    _zz_when_ArraySlice_l159_157_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_157_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_157_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_157_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_157_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_157_6;
  wire       [7:0]    _zz__zz_realValue_0_157;
  wire       [7:0]    _zz__zz_realValue_0_157_1;
  wire       [7:0]    _zz_realValue_0_157_1;
  wire       [7:0]    _zz_realValue_0_157_2;
  wire       [7:0]    _zz_realValue_0_157_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_157;
  wire       [5:0]    _zz_when_ArraySlice_l166_157_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_157_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_157_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_157_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_157_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_157_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_157_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_158;
  wire       [7:0]    _zz_when_ArraySlice_l158_158_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_158_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_158_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_158;
  wire       [5:0]    _zz_when_ArraySlice_l159_158_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_158_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_158_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_158_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_158_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_158_6;
  wire       [7:0]    _zz__zz_realValue_0_158;
  wire       [7:0]    _zz__zz_realValue_0_158_1;
  wire       [7:0]    _zz_realValue_0_158_1;
  wire       [7:0]    _zz_realValue_0_158_2;
  wire       [7:0]    _zz_realValue_0_158_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_158;
  wire       [5:0]    _zz_when_ArraySlice_l166_158_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_158_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_158_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_158_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_158_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_158_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_158_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_159;
  wire       [7:0]    _zz_when_ArraySlice_l158_159_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_159_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_159_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_159;
  wire       [4:0]    _zz_when_ArraySlice_l159_159_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_159_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_159_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_159_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_159_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_159_6;
  wire       [7:0]    _zz__zz_realValue_0_159;
  wire       [7:0]    _zz__zz_realValue_0_159_1;
  wire       [7:0]    _zz_realValue_0_159_1;
  wire       [7:0]    _zz_realValue_0_159_2;
  wire       [7:0]    _zz_realValue_0_159_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_159;
  wire       [4:0]    _zz_when_ArraySlice_l166_159_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_159_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_159_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_159_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_159_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_159_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_159_7;
  wire                _zz_when_ArraySlice_l400_6_1;
  wire                _zz_when_ArraySlice_l400_6_2;
  wire                _zz_when_ArraySlice_l400_6_3;
  wire                _zz_when_ArraySlice_l400_6_4;
  wire                _zz_when_ArraySlice_l400_6_5;
  wire                _zz_when_ArraySlice_l400_6_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_6_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_6_7;
  wire       [6:0]    _zz_when_ArraySlice_l403_6_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_6;
  wire       [7:0]    _zz_when_ArraySlice_l406_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l406_6_4;
  wire       [7:0]    _zz_selectReadFifo_6_6;
  wire       [7:0]    _zz_selectReadFifo_6_7;
  wire       [6:0]    _zz_selectReadFifo_6_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_6;
  wire       [12:0]   _zz_when_ArraySlice_l413_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_6;
  wire       [6:0]    _zz_when_ArraySlice_l417_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l417_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l417_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l418_6;
  wire       [7:0]    _zz_when_ArraySlice_l418_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l418_6_4;
  wire       [7:0]    _zz__zz_realValue1_0_19;
  wire       [7:0]    _zz__zz_realValue1_0_19_1;
  wire       [7:0]    _zz_realValue1_0_19_1;
  wire       [7:0]    _zz_realValue1_0_19_2;
  wire       [7:0]    _zz_realValue1_0_19_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_6;
  wire       [6:0]    _zz_when_ArraySlice_l420_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_9;
  wire       [7:0]    _zz_selectReadFifo_6_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_160;
  wire       [7:0]    _zz_when_ArraySlice_l158_160_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_160_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_160_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_160;
  wire       [7:0]    _zz_when_ArraySlice_l159_160_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_160_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_160_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_160_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_160_5;
  wire       [7:0]    _zz__zz_realValue_0_160;
  wire       [7:0]    _zz__zz_realValue_0_160_1;
  wire       [7:0]    _zz_realValue_0_160_1;
  wire       [7:0]    _zz_realValue_0_160_2;
  wire       [7:0]    _zz_realValue_0_160_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_160;
  wire       [7:0]    _zz_when_ArraySlice_l166_160_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_160_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_160_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_160_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_160_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_160_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_161;
  wire       [7:0]    _zz_when_ArraySlice_l158_161_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_161_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_161_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_161;
  wire       [6:0]    _zz_when_ArraySlice_l159_161_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_161_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_161_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_161_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_161_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_161_6;
  wire       [7:0]    _zz__zz_realValue_0_161;
  wire       [7:0]    _zz__zz_realValue_0_161_1;
  wire       [7:0]    _zz_realValue_0_161_1;
  wire       [7:0]    _zz_realValue_0_161_2;
  wire       [7:0]    _zz_realValue_0_161_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_161;
  wire       [6:0]    _zz_when_ArraySlice_l166_161_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_161_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_161_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_161_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_161_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_161_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_161_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_162;
  wire       [7:0]    _zz_when_ArraySlice_l158_162_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_162_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_162_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_162;
  wire       [6:0]    _zz_when_ArraySlice_l159_162_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_162_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_162_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_162_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_162_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_162_6;
  wire       [7:0]    _zz__zz_realValue_0_162;
  wire       [7:0]    _zz__zz_realValue_0_162_1;
  wire       [7:0]    _zz_realValue_0_162_1;
  wire       [7:0]    _zz_realValue_0_162_2;
  wire       [7:0]    _zz_realValue_0_162_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_162;
  wire       [6:0]    _zz_when_ArraySlice_l166_162_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_162_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_162_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_162_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_162_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_162_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_162_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_163;
  wire       [7:0]    _zz_when_ArraySlice_l158_163_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_163_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_163_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_163;
  wire       [6:0]    _zz_when_ArraySlice_l159_163_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_163_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_163_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_163_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_163_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_163_6;
  wire       [7:0]    _zz__zz_realValue_0_163;
  wire       [7:0]    _zz__zz_realValue_0_163_1;
  wire       [7:0]    _zz_realValue_0_163_1;
  wire       [7:0]    _zz_realValue_0_163_2;
  wire       [7:0]    _zz_realValue_0_163_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_163;
  wire       [6:0]    _zz_when_ArraySlice_l166_163_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_163_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_163_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_163_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_163_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_163_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_163_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_164;
  wire       [7:0]    _zz_when_ArraySlice_l158_164_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_164_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_164_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_164;
  wire       [6:0]    _zz_when_ArraySlice_l159_164_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_164_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_164_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_164_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_164_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_164_6;
  wire       [7:0]    _zz__zz_realValue_0_164;
  wire       [7:0]    _zz__zz_realValue_0_164_1;
  wire       [7:0]    _zz_realValue_0_164_1;
  wire       [7:0]    _zz_realValue_0_164_2;
  wire       [7:0]    _zz_realValue_0_164_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_164;
  wire       [6:0]    _zz_when_ArraySlice_l166_164_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_164_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_164_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_164_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_164_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_164_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_164_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_165;
  wire       [7:0]    _zz_when_ArraySlice_l158_165_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_165_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_165_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_165;
  wire       [5:0]    _zz_when_ArraySlice_l159_165_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_165_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_165_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_165_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_165_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_165_6;
  wire       [7:0]    _zz__zz_realValue_0_165;
  wire       [7:0]    _zz__zz_realValue_0_165_1;
  wire       [7:0]    _zz_realValue_0_165_1;
  wire       [7:0]    _zz_realValue_0_165_2;
  wire       [7:0]    _zz_realValue_0_165_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_165;
  wire       [5:0]    _zz_when_ArraySlice_l166_165_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_165_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_165_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_165_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_165_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_165_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_165_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_166;
  wire       [7:0]    _zz_when_ArraySlice_l158_166_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_166_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_166_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_166;
  wire       [5:0]    _zz_when_ArraySlice_l159_166_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_166_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_166_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_166_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_166_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_166_6;
  wire       [7:0]    _zz__zz_realValue_0_166;
  wire       [7:0]    _zz__zz_realValue_0_166_1;
  wire       [7:0]    _zz_realValue_0_166_1;
  wire       [7:0]    _zz_realValue_0_166_2;
  wire       [7:0]    _zz_realValue_0_166_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_166;
  wire       [5:0]    _zz_when_ArraySlice_l166_166_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_166_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_166_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_166_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_166_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_166_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_166_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_167;
  wire       [7:0]    _zz_when_ArraySlice_l158_167_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_167_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_167_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_167;
  wire       [4:0]    _zz_when_ArraySlice_l159_167_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_167_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_167_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_167_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_167_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_167_6;
  wire       [7:0]    _zz__zz_realValue_0_167;
  wire       [7:0]    _zz__zz_realValue_0_167_1;
  wire       [7:0]    _zz_realValue_0_167_1;
  wire       [7:0]    _zz_realValue_0_167_2;
  wire       [7:0]    _zz_realValue_0_167_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_167;
  wire       [4:0]    _zz_when_ArraySlice_l166_167_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_167_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_167_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_167_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_167_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_167_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_167_7;
  wire                _zz_when_ArraySlice_l425_6;
  wire                _zz_when_ArraySlice_l425_6_1;
  wire                _zz_when_ArraySlice_l425_6_2;
  wire                _zz_when_ArraySlice_l425_6_3;
  wire                _zz_when_ArraySlice_l425_6_4;
  wire                _zz_when_ArraySlice_l425_6_5;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_6_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_6_7;
  wire       [6:0]    _zz_when_ArraySlice_l428_6_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_6;
  wire       [7:0]    _zz_when_ArraySlice_l431_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l431_6_4;
  wire       [7:0]    _zz_selectReadFifo_6_11;
  wire       [7:0]    _zz_selectReadFifo_6_12;
  wire       [6:0]    _zz_selectReadFifo_6_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_6;
  wire       [12:0]   _zz_when_ArraySlice_l438_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_6;
  wire       [7:0]    _zz_when_ArraySlice_l449_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_6_2;
  wire       [7:0]    _zz__zz_realValue1_0_20;
  wire       [7:0]    _zz__zz_realValue1_0_20_1;
  wire       [7:0]    _zz_realValue1_0_20_1;
  wire       [7:0]    _zz_realValue1_0_20_2;
  wire       [7:0]    _zz_realValue1_0_20_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_6;
  wire       [6:0]    _zz_when_ArraySlice_l450_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_14;
  wire       [7:0]    _zz_selectReadFifo_6_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_168;
  wire       [7:0]    _zz_when_ArraySlice_l158_168_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_168_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_168_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_168;
  wire       [7:0]    _zz_when_ArraySlice_l159_168_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_168_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_168_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_168_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_168_5;
  wire       [7:0]    _zz__zz_realValue_0_168;
  wire       [7:0]    _zz__zz_realValue_0_168_1;
  wire       [7:0]    _zz_realValue_0_168_1;
  wire       [7:0]    _zz_realValue_0_168_2;
  wire       [7:0]    _zz_realValue_0_168_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_168;
  wire       [7:0]    _zz_when_ArraySlice_l166_168_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_168_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_168_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_168_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_168_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_168_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_169;
  wire       [7:0]    _zz_when_ArraySlice_l158_169_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_169_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_169_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_169;
  wire       [6:0]    _zz_when_ArraySlice_l159_169_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_169_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_169_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_169_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_169_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_169_6;
  wire       [7:0]    _zz__zz_realValue_0_169;
  wire       [7:0]    _zz__zz_realValue_0_169_1;
  wire       [7:0]    _zz_realValue_0_169_1;
  wire       [7:0]    _zz_realValue_0_169_2;
  wire       [7:0]    _zz_realValue_0_169_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_169;
  wire       [6:0]    _zz_when_ArraySlice_l166_169_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_169_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_169_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_169_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_169_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_169_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_169_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_170;
  wire       [7:0]    _zz_when_ArraySlice_l158_170_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_170_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_170_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_170;
  wire       [6:0]    _zz_when_ArraySlice_l159_170_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_170_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_170_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_170_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_170_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_170_6;
  wire       [7:0]    _zz__zz_realValue_0_170;
  wire       [7:0]    _zz__zz_realValue_0_170_1;
  wire       [7:0]    _zz_realValue_0_170_1;
  wire       [7:0]    _zz_realValue_0_170_2;
  wire       [7:0]    _zz_realValue_0_170_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_170;
  wire       [6:0]    _zz_when_ArraySlice_l166_170_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_170_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_170_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_170_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_170_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_170_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_170_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_171;
  wire       [7:0]    _zz_when_ArraySlice_l158_171_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_171_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_171_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_171;
  wire       [6:0]    _zz_when_ArraySlice_l159_171_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_171_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_171_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_171_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_171_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_171_6;
  wire       [7:0]    _zz__zz_realValue_0_171;
  wire       [7:0]    _zz__zz_realValue_0_171_1;
  wire       [7:0]    _zz_realValue_0_171_1;
  wire       [7:0]    _zz_realValue_0_171_2;
  wire       [7:0]    _zz_realValue_0_171_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_171;
  wire       [6:0]    _zz_when_ArraySlice_l166_171_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_171_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_171_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_171_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_171_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_171_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_171_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_172;
  wire       [7:0]    _zz_when_ArraySlice_l158_172_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_172_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_172_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_172;
  wire       [6:0]    _zz_when_ArraySlice_l159_172_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_172_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_172_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_172_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_172_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_172_6;
  wire       [7:0]    _zz__zz_realValue_0_172;
  wire       [7:0]    _zz__zz_realValue_0_172_1;
  wire       [7:0]    _zz_realValue_0_172_1;
  wire       [7:0]    _zz_realValue_0_172_2;
  wire       [7:0]    _zz_realValue_0_172_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_172;
  wire       [6:0]    _zz_when_ArraySlice_l166_172_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_172_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_172_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_172_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_172_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_172_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_172_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_173;
  wire       [7:0]    _zz_when_ArraySlice_l158_173_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_173_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_173_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_173;
  wire       [5:0]    _zz_when_ArraySlice_l159_173_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_173_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_173_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_173_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_173_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_173_6;
  wire       [7:0]    _zz__zz_realValue_0_173;
  wire       [7:0]    _zz__zz_realValue_0_173_1;
  wire       [7:0]    _zz_realValue_0_173_1;
  wire       [7:0]    _zz_realValue_0_173_2;
  wire       [7:0]    _zz_realValue_0_173_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_173;
  wire       [5:0]    _zz_when_ArraySlice_l166_173_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_173_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_173_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_173_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_173_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_173_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_173_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_174;
  wire       [7:0]    _zz_when_ArraySlice_l158_174_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_174_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_174_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_174;
  wire       [5:0]    _zz_when_ArraySlice_l159_174_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_174_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_174_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_174_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_174_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_174_6;
  wire       [7:0]    _zz__zz_realValue_0_174;
  wire       [7:0]    _zz__zz_realValue_0_174_1;
  wire       [7:0]    _zz_realValue_0_174_1;
  wire       [7:0]    _zz_realValue_0_174_2;
  wire       [7:0]    _zz_realValue_0_174_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_174;
  wire       [5:0]    _zz_when_ArraySlice_l166_174_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_174_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_174_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_174_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_174_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_174_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_174_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_175;
  wire       [7:0]    _zz_when_ArraySlice_l158_175_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_175_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_175_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_175;
  wire       [4:0]    _zz_when_ArraySlice_l159_175_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_175_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_175_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_175_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_175_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_175_6;
  wire       [7:0]    _zz__zz_realValue_0_175;
  wire       [7:0]    _zz__zz_realValue_0_175_1;
  wire       [7:0]    _zz_realValue_0_175_1;
  wire       [7:0]    _zz_realValue_0_175_2;
  wire       [7:0]    _zz_realValue_0_175_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_175;
  wire       [4:0]    _zz_when_ArraySlice_l166_175_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_175_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_175_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_175_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_175_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_175_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_175_7;
  wire                _zz_when_ArraySlice_l457_6;
  wire                _zz_when_ArraySlice_l457_6_1;
  wire                _zz_when_ArraySlice_l457_6_2;
  wire                _zz_when_ArraySlice_l457_6_3;
  wire                _zz_when_ArraySlice_l457_6_4;
  wire                _zz_when_ArraySlice_l457_6_5;
  wire       [12:0]   _zz_when_ArraySlice_l461_6;
  wire       [12:0]   _zz_when_ArraySlice_l461_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_6;
  wire       [7:0]    _zz_when_ArraySlice_l447_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l447_6_3;
  wire       [12:0]   _zz_when_ArraySlice_l468_6;
  wire       [7:0]    _zz_when_ArraySlice_l468_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_7;
  wire       [7:0]    _zz_when_ArraySlice_l376_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l376_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l376_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l377_7;
  wire       [6:0]    _zz_when_ArraySlice_l377_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l377_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l377_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l377_7_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_7_valid;
  wire       [6:0]    _zz__zz_outputStreamArrayData_7_valid_1;
  wire       [6:0]    _zz__zz_10;
  reg                 _zz_outputStreamArrayData_7_valid_2;
  wire       [6:0]    _zz_outputStreamArrayData_7_valid_3;
  reg        [31:0]   _zz_outputStreamArrayData_7_payload;
  wire       [6:0]    _zz_outputStreamArrayData_7_payload_1;
  reg        [6:0]    _zz_when_ArraySlice_l383_7;
  wire       [6:0]    _zz_when_ArraySlice_l383_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l383_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l383_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l383_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l384_7;
  wire       [7:0]    _zz_when_ArraySlice_l384_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l384_7_2;
  wire       [7:0]    _zz_selectReadFifo_7;
  wire       [7:0]    _zz_selectReadFifo_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l387_7;
  wire       [12:0]   _zz_when_ArraySlice_l387_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l392_7;
  wire       [6:0]    _zz_when_ArraySlice_l392_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l392_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l392_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l392_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l393_7;
  wire       [7:0]    _zz_when_ArraySlice_l393_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l393_7_2;
  wire       [7:0]    _zz__zz_realValue1_0_21;
  wire       [7:0]    _zz__zz_realValue1_0_21_1;
  wire       [7:0]    _zz_realValue1_0_21_1;
  wire       [7:0]    _zz_realValue1_0_21_2;
  wire       [7:0]    _zz_realValue1_0_21_3;
  wire       [7:0]    _zz_when_ArraySlice_l395_7;
  wire       [6:0]    _zz_when_ArraySlice_l395_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l395_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_3;
  wire       [7:0]    _zz_selectReadFifo_7_4;
  wire       [0:0]    _zz_selectReadFifo_7_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_176;
  wire       [7:0]    _zz_when_ArraySlice_l158_176_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_176_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_176_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_176;
  wire       [7:0]    _zz_when_ArraySlice_l159_176_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_176_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_176_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_176_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_176_5;
  wire       [7:0]    _zz__zz_realValue_0_176;
  wire       [7:0]    _zz__zz_realValue_0_176_1;
  wire       [7:0]    _zz_realValue_0_176_1;
  wire       [7:0]    _zz_realValue_0_176_2;
  wire       [7:0]    _zz_realValue_0_176_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_176;
  wire       [7:0]    _zz_when_ArraySlice_l166_176_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_176_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_176_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_176_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_176_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_176_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_177;
  wire       [7:0]    _zz_when_ArraySlice_l158_177_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_177_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_177_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_177;
  wire       [6:0]    _zz_when_ArraySlice_l159_177_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_177_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_177_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_177_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_177_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_177_6;
  wire       [7:0]    _zz__zz_realValue_0_177;
  wire       [7:0]    _zz__zz_realValue_0_177_1;
  wire       [7:0]    _zz_realValue_0_177_1;
  wire       [7:0]    _zz_realValue_0_177_2;
  wire       [7:0]    _zz_realValue_0_177_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_177;
  wire       [6:0]    _zz_when_ArraySlice_l166_177_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_177_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_177_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_177_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_177_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_177_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_177_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_178;
  wire       [7:0]    _zz_when_ArraySlice_l158_178_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_178_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_178_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_178;
  wire       [6:0]    _zz_when_ArraySlice_l159_178_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_178_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_178_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_178_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_178_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_178_6;
  wire       [7:0]    _zz__zz_realValue_0_178;
  wire       [7:0]    _zz__zz_realValue_0_178_1;
  wire       [7:0]    _zz_realValue_0_178_1;
  wire       [7:0]    _zz_realValue_0_178_2;
  wire       [7:0]    _zz_realValue_0_178_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_178;
  wire       [6:0]    _zz_when_ArraySlice_l166_178_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_178_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_178_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_178_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_178_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_178_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_178_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_179;
  wire       [7:0]    _zz_when_ArraySlice_l158_179_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_179_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_179_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_179;
  wire       [6:0]    _zz_when_ArraySlice_l159_179_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_179_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_179_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_179_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_179_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_179_6;
  wire       [7:0]    _zz__zz_realValue_0_179;
  wire       [7:0]    _zz__zz_realValue_0_179_1;
  wire       [7:0]    _zz_realValue_0_179_1;
  wire       [7:0]    _zz_realValue_0_179_2;
  wire       [7:0]    _zz_realValue_0_179_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_179;
  wire       [6:0]    _zz_when_ArraySlice_l166_179_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_179_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_179_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_179_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_179_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_179_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_179_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_180;
  wire       [7:0]    _zz_when_ArraySlice_l158_180_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_180_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_180_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_180;
  wire       [6:0]    _zz_when_ArraySlice_l159_180_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_180_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_180_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_180_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_180_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_180_6;
  wire       [7:0]    _zz__zz_realValue_0_180;
  wire       [7:0]    _zz__zz_realValue_0_180_1;
  wire       [7:0]    _zz_realValue_0_180_1;
  wire       [7:0]    _zz_realValue_0_180_2;
  wire       [7:0]    _zz_realValue_0_180_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_180;
  wire       [6:0]    _zz_when_ArraySlice_l166_180_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_180_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_180_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_180_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_180_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_180_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_180_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_181;
  wire       [7:0]    _zz_when_ArraySlice_l158_181_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_181_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_181_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_181;
  wire       [5:0]    _zz_when_ArraySlice_l159_181_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_181_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_181_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_181_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_181_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_181_6;
  wire       [7:0]    _zz__zz_realValue_0_181;
  wire       [7:0]    _zz__zz_realValue_0_181_1;
  wire       [7:0]    _zz_realValue_0_181_1;
  wire       [7:0]    _zz_realValue_0_181_2;
  wire       [7:0]    _zz_realValue_0_181_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_181;
  wire       [5:0]    _zz_when_ArraySlice_l166_181_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_181_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_181_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_181_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_181_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_181_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_181_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_182;
  wire       [7:0]    _zz_when_ArraySlice_l158_182_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_182_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_182_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_182;
  wire       [5:0]    _zz_when_ArraySlice_l159_182_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_182_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_182_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_182_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_182_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_182_6;
  wire       [7:0]    _zz__zz_realValue_0_182;
  wire       [7:0]    _zz__zz_realValue_0_182_1;
  wire       [7:0]    _zz_realValue_0_182_1;
  wire       [7:0]    _zz_realValue_0_182_2;
  wire       [7:0]    _zz_realValue_0_182_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_182;
  wire       [5:0]    _zz_when_ArraySlice_l166_182_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_182_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_182_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_182_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_182_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_182_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_182_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_183;
  wire       [7:0]    _zz_when_ArraySlice_l158_183_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_183_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_183_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_183;
  wire       [4:0]    _zz_when_ArraySlice_l159_183_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_183_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_183_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_183_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_183_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_183_6;
  wire       [7:0]    _zz__zz_realValue_0_183;
  wire       [7:0]    _zz__zz_realValue_0_183_1;
  wire       [7:0]    _zz_realValue_0_183_1;
  wire       [7:0]    _zz_realValue_0_183_2;
  wire       [7:0]    _zz_realValue_0_183_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_183;
  wire       [4:0]    _zz_when_ArraySlice_l166_183_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_183_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_183_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_183_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_183_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_183_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_183_7;
  wire                _zz_when_ArraySlice_l400_7_1;
  wire                _zz_when_ArraySlice_l400_7_2;
  wire                _zz_when_ArraySlice_l400_7_3;
  wire                _zz_when_ArraySlice_l400_7_4;
  wire                _zz_when_ArraySlice_l400_7_5;
  wire                _zz_when_ArraySlice_l400_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l403_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l403_7_7;
  wire       [6:0]    _zz_when_ArraySlice_l403_7_8;
  wire       [7:0]    _zz_when_ArraySlice_l406_7;
  wire       [7:0]    _zz_when_ArraySlice_l406_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l406_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l406_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l406_7_4;
  wire       [7:0]    _zz_selectReadFifo_7_6;
  wire       [7:0]    _zz_selectReadFifo_7_7;
  wire       [6:0]    _zz_selectReadFifo_7_8;
  wire       [12:0]   _zz_when_ArraySlice_l413_7;
  wire       [12:0]   _zz_when_ArraySlice_l413_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l417_7;
  wire       [6:0]    _zz_when_ArraySlice_l417_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l417_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l417_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l417_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l418_7;
  wire       [7:0]    _zz_when_ArraySlice_l418_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l418_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l418_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l418_7_4;
  wire       [7:0]    _zz__zz_realValue1_0_22;
  wire       [7:0]    _zz__zz_realValue1_0_22_1;
  wire       [7:0]    _zz_realValue1_0_22_1;
  wire       [7:0]    _zz_realValue1_0_22_2;
  wire       [7:0]    _zz_realValue1_0_22_3;
  wire       [7:0]    _zz_when_ArraySlice_l420_7;
  wire       [6:0]    _zz_when_ArraySlice_l420_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l420_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_9;
  wire       [7:0]    _zz_selectReadFifo_7_10;
  wire       [7:0]    _zz_when_ArraySlice_l158_184;
  wire       [7:0]    _zz_when_ArraySlice_l158_184_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_184_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_184_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_184;
  wire       [7:0]    _zz_when_ArraySlice_l159_184_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_184_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_184_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_184_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_184_5;
  wire       [7:0]    _zz__zz_realValue_0_184;
  wire       [7:0]    _zz__zz_realValue_0_184_1;
  wire       [7:0]    _zz_realValue_0_184_1;
  wire       [7:0]    _zz_realValue_0_184_2;
  wire       [7:0]    _zz_realValue_0_184_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_184;
  wire       [7:0]    _zz_when_ArraySlice_l166_184_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_184_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_184_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_184_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_184_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_184_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_185;
  wire       [7:0]    _zz_when_ArraySlice_l158_185_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_185_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_185_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_185;
  wire       [6:0]    _zz_when_ArraySlice_l159_185_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_185_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_185_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_185_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_185_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_185_6;
  wire       [7:0]    _zz__zz_realValue_0_185;
  wire       [7:0]    _zz__zz_realValue_0_185_1;
  wire       [7:0]    _zz_realValue_0_185_1;
  wire       [7:0]    _zz_realValue_0_185_2;
  wire       [7:0]    _zz_realValue_0_185_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_185;
  wire       [6:0]    _zz_when_ArraySlice_l166_185_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_185_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_185_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_185_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_185_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_185_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_185_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_186;
  wire       [7:0]    _zz_when_ArraySlice_l158_186_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_186_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_186_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_186;
  wire       [6:0]    _zz_when_ArraySlice_l159_186_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_186_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_186_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_186_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_186_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_186_6;
  wire       [7:0]    _zz__zz_realValue_0_186;
  wire       [7:0]    _zz__zz_realValue_0_186_1;
  wire       [7:0]    _zz_realValue_0_186_1;
  wire       [7:0]    _zz_realValue_0_186_2;
  wire       [7:0]    _zz_realValue_0_186_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_186;
  wire       [6:0]    _zz_when_ArraySlice_l166_186_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_186_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_186_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_186_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_186_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_186_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_186_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_187;
  wire       [7:0]    _zz_when_ArraySlice_l158_187_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_187_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_187_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_187;
  wire       [6:0]    _zz_when_ArraySlice_l159_187_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_187_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_187_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_187_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_187_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_187_6;
  wire       [7:0]    _zz__zz_realValue_0_187;
  wire       [7:0]    _zz__zz_realValue_0_187_1;
  wire       [7:0]    _zz_realValue_0_187_1;
  wire       [7:0]    _zz_realValue_0_187_2;
  wire       [7:0]    _zz_realValue_0_187_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_187;
  wire       [6:0]    _zz_when_ArraySlice_l166_187_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_187_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_187_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_187_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_187_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_187_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_187_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_188;
  wire       [7:0]    _zz_when_ArraySlice_l158_188_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_188_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_188_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_188;
  wire       [6:0]    _zz_when_ArraySlice_l159_188_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_188_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_188_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_188_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_188_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_188_6;
  wire       [7:0]    _zz__zz_realValue_0_188;
  wire       [7:0]    _zz__zz_realValue_0_188_1;
  wire       [7:0]    _zz_realValue_0_188_1;
  wire       [7:0]    _zz_realValue_0_188_2;
  wire       [7:0]    _zz_realValue_0_188_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_188;
  wire       [6:0]    _zz_when_ArraySlice_l166_188_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_188_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_188_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_188_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_188_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_188_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_188_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_189;
  wire       [7:0]    _zz_when_ArraySlice_l158_189_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_189_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_189_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_189;
  wire       [5:0]    _zz_when_ArraySlice_l159_189_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_189_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_189_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_189_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_189_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_189_6;
  wire       [7:0]    _zz__zz_realValue_0_189;
  wire       [7:0]    _zz__zz_realValue_0_189_1;
  wire       [7:0]    _zz_realValue_0_189_1;
  wire       [7:0]    _zz_realValue_0_189_2;
  wire       [7:0]    _zz_realValue_0_189_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_189;
  wire       [5:0]    _zz_when_ArraySlice_l166_189_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_189_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_189_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_189_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_189_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_189_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_189_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_190;
  wire       [7:0]    _zz_when_ArraySlice_l158_190_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_190_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_190_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_190;
  wire       [5:0]    _zz_when_ArraySlice_l159_190_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_190_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_190_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_190_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_190_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_190_6;
  wire       [7:0]    _zz__zz_realValue_0_190;
  wire       [7:0]    _zz__zz_realValue_0_190_1;
  wire       [7:0]    _zz_realValue_0_190_1;
  wire       [7:0]    _zz_realValue_0_190_2;
  wire       [7:0]    _zz_realValue_0_190_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_190;
  wire       [5:0]    _zz_when_ArraySlice_l166_190_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_190_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_190_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_190_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_190_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_190_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_190_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_191;
  wire       [7:0]    _zz_when_ArraySlice_l158_191_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_191_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_191_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_191;
  wire       [4:0]    _zz_when_ArraySlice_l159_191_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_191_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_191_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_191_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_191_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_191_6;
  wire       [7:0]    _zz__zz_realValue_0_191;
  wire       [7:0]    _zz__zz_realValue_0_191_1;
  wire       [7:0]    _zz_realValue_0_191_1;
  wire       [7:0]    _zz_realValue_0_191_2;
  wire       [7:0]    _zz_realValue_0_191_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_191;
  wire       [4:0]    _zz_when_ArraySlice_l166_191_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_191_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_191_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_191_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_191_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_191_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_191_7;
  wire                _zz_when_ArraySlice_l425_7;
  wire                _zz_when_ArraySlice_l425_7_1;
  wire                _zz_when_ArraySlice_l425_7_2;
  wire                _zz_when_ArraySlice_l425_7_3;
  wire                _zz_when_ArraySlice_l425_7_4;
  wire                _zz_when_ArraySlice_l425_7_5;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l428_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l428_7_7;
  wire       [6:0]    _zz_when_ArraySlice_l428_7_8;
  wire       [7:0]    _zz_when_ArraySlice_l431_7;
  wire       [7:0]    _zz_when_ArraySlice_l431_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l431_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l431_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l431_7_4;
  wire       [7:0]    _zz_selectReadFifo_7_11;
  wire       [7:0]    _zz_selectReadFifo_7_12;
  wire       [6:0]    _zz_selectReadFifo_7_13;
  wire       [12:0]   _zz_when_ArraySlice_l438_7;
  wire       [12:0]   _zz_when_ArraySlice_l438_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l449_7;
  wire       [7:0]    _zz_when_ArraySlice_l449_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l449_7_2;
  wire       [7:0]    _zz__zz_realValue1_0_23;
  wire       [7:0]    _zz__zz_realValue1_0_23_1;
  wire       [7:0]    _zz_realValue1_0_23_1;
  wire       [7:0]    _zz_realValue1_0_23_2;
  wire       [7:0]    _zz_realValue1_0_23_3;
  wire       [7:0]    _zz_when_ArraySlice_l450_7;
  wire       [6:0]    _zz_when_ArraySlice_l450_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l450_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_14;
  wire       [7:0]    _zz_selectReadFifo_7_15;
  wire       [7:0]    _zz_when_ArraySlice_l158_192;
  wire       [7:0]    _zz_when_ArraySlice_l158_192_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_192_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_192_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_192;
  wire       [7:0]    _zz_when_ArraySlice_l159_192_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_192_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_192_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_192_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_192_5;
  wire       [7:0]    _zz__zz_realValue_0_192;
  wire       [7:0]    _zz__zz_realValue_0_192_1;
  wire       [7:0]    _zz_realValue_0_192_1;
  wire       [7:0]    _zz_realValue_0_192_2;
  wire       [7:0]    _zz_realValue_0_192_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_192;
  wire       [7:0]    _zz_when_ArraySlice_l166_192_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_192_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_192_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_192_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_192_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_192_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_193;
  wire       [7:0]    _zz_when_ArraySlice_l158_193_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_193_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_193_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_193;
  wire       [6:0]    _zz_when_ArraySlice_l159_193_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_193_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_193_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_193_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_193_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_193_6;
  wire       [7:0]    _zz__zz_realValue_0_193;
  wire       [7:0]    _zz__zz_realValue_0_193_1;
  wire       [7:0]    _zz_realValue_0_193_1;
  wire       [7:0]    _zz_realValue_0_193_2;
  wire       [7:0]    _zz_realValue_0_193_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_193;
  wire       [6:0]    _zz_when_ArraySlice_l166_193_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_193_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_193_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_193_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_193_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_193_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_193_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_194;
  wire       [7:0]    _zz_when_ArraySlice_l158_194_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_194_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_194_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_194;
  wire       [6:0]    _zz_when_ArraySlice_l159_194_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_194_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_194_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_194_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_194_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_194_6;
  wire       [7:0]    _zz__zz_realValue_0_194;
  wire       [7:0]    _zz__zz_realValue_0_194_1;
  wire       [7:0]    _zz_realValue_0_194_1;
  wire       [7:0]    _zz_realValue_0_194_2;
  wire       [7:0]    _zz_realValue_0_194_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_194;
  wire       [6:0]    _zz_when_ArraySlice_l166_194_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_194_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_194_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_194_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_194_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_194_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_194_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_195;
  wire       [7:0]    _zz_when_ArraySlice_l158_195_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_195_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_195_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_195;
  wire       [6:0]    _zz_when_ArraySlice_l159_195_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_195_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_195_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_195_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_195_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_195_6;
  wire       [7:0]    _zz__zz_realValue_0_195;
  wire       [7:0]    _zz__zz_realValue_0_195_1;
  wire       [7:0]    _zz_realValue_0_195_1;
  wire       [7:0]    _zz_realValue_0_195_2;
  wire       [7:0]    _zz_realValue_0_195_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_195;
  wire       [6:0]    _zz_when_ArraySlice_l166_195_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_195_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_195_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_195_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_195_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_195_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_195_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_196;
  wire       [7:0]    _zz_when_ArraySlice_l158_196_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_196_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_196_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_196;
  wire       [6:0]    _zz_when_ArraySlice_l159_196_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_196_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_196_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_196_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_196_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_196_6;
  wire       [7:0]    _zz__zz_realValue_0_196;
  wire       [7:0]    _zz__zz_realValue_0_196_1;
  wire       [7:0]    _zz_realValue_0_196_1;
  wire       [7:0]    _zz_realValue_0_196_2;
  wire       [7:0]    _zz_realValue_0_196_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_196;
  wire       [6:0]    _zz_when_ArraySlice_l166_196_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_196_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_196_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_196_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_196_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_196_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_196_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_197;
  wire       [7:0]    _zz_when_ArraySlice_l158_197_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_197_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_197_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_197;
  wire       [5:0]    _zz_when_ArraySlice_l159_197_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_197_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_197_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_197_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_197_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_197_6;
  wire       [7:0]    _zz__zz_realValue_0_197;
  wire       [7:0]    _zz__zz_realValue_0_197_1;
  wire       [7:0]    _zz_realValue_0_197_1;
  wire       [7:0]    _zz_realValue_0_197_2;
  wire       [7:0]    _zz_realValue_0_197_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_197;
  wire       [5:0]    _zz_when_ArraySlice_l166_197_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_197_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_197_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_197_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_197_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_197_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_197_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_198;
  wire       [7:0]    _zz_when_ArraySlice_l158_198_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_198_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_198_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_198;
  wire       [5:0]    _zz_when_ArraySlice_l159_198_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_198_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_198_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_198_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_198_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_198_6;
  wire       [7:0]    _zz__zz_realValue_0_198;
  wire       [7:0]    _zz__zz_realValue_0_198_1;
  wire       [7:0]    _zz_realValue_0_198_1;
  wire       [7:0]    _zz_realValue_0_198_2;
  wire       [7:0]    _zz_realValue_0_198_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_198;
  wire       [5:0]    _zz_when_ArraySlice_l166_198_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_198_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_198_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_198_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_198_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_198_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_198_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_199;
  wire       [7:0]    _zz_when_ArraySlice_l158_199_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_199_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_199_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_199;
  wire       [4:0]    _zz_when_ArraySlice_l159_199_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_199_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_199_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_199_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_199_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_199_6;
  wire       [7:0]    _zz__zz_realValue_0_199;
  wire       [7:0]    _zz__zz_realValue_0_199_1;
  wire       [7:0]    _zz_realValue_0_199_1;
  wire       [7:0]    _zz_realValue_0_199_2;
  wire       [7:0]    _zz_realValue_0_199_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_199;
  wire       [4:0]    _zz_when_ArraySlice_l166_199_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_199_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_199_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_199_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_199_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_199_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_199_7;
  wire                _zz_when_ArraySlice_l457_7;
  wire                _zz_when_ArraySlice_l457_7_1;
  wire                _zz_when_ArraySlice_l457_7_2;
  wire                _zz_when_ArraySlice_l457_7_3;
  wire                _zz_when_ArraySlice_l457_7_4;
  wire                _zz_when_ArraySlice_l457_7_5;
  wire       [12:0]   _zz_when_ArraySlice_l461_7;
  wire       [12:0]   _zz_when_ArraySlice_l461_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_7;
  wire       [7:0]    _zz_when_ArraySlice_l447_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l447_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l447_7_3;
  wire       [12:0]   _zz_when_ArraySlice_l468_7;
  wire       [7:0]    _zz_when_ArraySlice_l468_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l468_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_200;
  wire       [7:0]    _zz_when_ArraySlice_l158_200_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_200_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_200_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_200;
  wire       [7:0]    _zz_when_ArraySlice_l159_200_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_200_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_200_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_200_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_200_5;
  wire       [7:0]    _zz__zz_realValue_0_200;
  wire       [7:0]    _zz__zz_realValue_0_200_1;
  wire       [7:0]    _zz_realValue_0_200_1;
  wire       [7:0]    _zz_realValue_0_200_2;
  wire       [7:0]    _zz_realValue_0_200_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_200;
  wire       [7:0]    _zz_when_ArraySlice_l166_200_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_200_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_200_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_200_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_200_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_200_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_201;
  wire       [7:0]    _zz_when_ArraySlice_l158_201_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_201_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_201_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_201;
  wire       [6:0]    _zz_when_ArraySlice_l159_201_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_201_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_201_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_201_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_201_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_201_6;
  wire       [7:0]    _zz__zz_realValue_0_201;
  wire       [7:0]    _zz__zz_realValue_0_201_1;
  wire       [7:0]    _zz_realValue_0_201_1;
  wire       [7:0]    _zz_realValue_0_201_2;
  wire       [7:0]    _zz_realValue_0_201_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_201;
  wire       [6:0]    _zz_when_ArraySlice_l166_201_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_201_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_201_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_201_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_201_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_201_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_201_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_202;
  wire       [7:0]    _zz_when_ArraySlice_l158_202_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_202_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_202_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_202;
  wire       [6:0]    _zz_when_ArraySlice_l159_202_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_202_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_202_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_202_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_202_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_202_6;
  wire       [7:0]    _zz__zz_realValue_0_202;
  wire       [7:0]    _zz__zz_realValue_0_202_1;
  wire       [7:0]    _zz_realValue_0_202_1;
  wire       [7:0]    _zz_realValue_0_202_2;
  wire       [7:0]    _zz_realValue_0_202_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_202;
  wire       [6:0]    _zz_when_ArraySlice_l166_202_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_202_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_202_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_202_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_202_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_202_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_202_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_203;
  wire       [7:0]    _zz_when_ArraySlice_l158_203_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_203_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_203_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_203;
  wire       [6:0]    _zz_when_ArraySlice_l159_203_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_203_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_203_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_203_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_203_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_203_6;
  wire       [7:0]    _zz__zz_realValue_0_203;
  wire       [7:0]    _zz__zz_realValue_0_203_1;
  wire       [7:0]    _zz_realValue_0_203_1;
  wire       [7:0]    _zz_realValue_0_203_2;
  wire       [7:0]    _zz_realValue_0_203_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_203;
  wire       [6:0]    _zz_when_ArraySlice_l166_203_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_203_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_203_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_203_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_203_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_203_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_203_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_204;
  wire       [7:0]    _zz_when_ArraySlice_l158_204_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_204_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_204_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_204;
  wire       [6:0]    _zz_when_ArraySlice_l159_204_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_204_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_204_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_204_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_204_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_204_6;
  wire       [7:0]    _zz__zz_realValue_0_204;
  wire       [7:0]    _zz__zz_realValue_0_204_1;
  wire       [7:0]    _zz_realValue_0_204_1;
  wire       [7:0]    _zz_realValue_0_204_2;
  wire       [7:0]    _zz_realValue_0_204_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_204;
  wire       [6:0]    _zz_when_ArraySlice_l166_204_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_204_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_204_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_204_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_204_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_204_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_204_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_205;
  wire       [7:0]    _zz_when_ArraySlice_l158_205_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_205_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_205_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_205;
  wire       [5:0]    _zz_when_ArraySlice_l159_205_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_205_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_205_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_205_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_205_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_205_6;
  wire       [7:0]    _zz__zz_realValue_0_205;
  wire       [7:0]    _zz__zz_realValue_0_205_1;
  wire       [7:0]    _zz_realValue_0_205_1;
  wire       [7:0]    _zz_realValue_0_205_2;
  wire       [7:0]    _zz_realValue_0_205_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_205;
  wire       [5:0]    _zz_when_ArraySlice_l166_205_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_205_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_205_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_205_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_205_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_205_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_205_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_206;
  wire       [7:0]    _zz_when_ArraySlice_l158_206_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_206_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_206_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_206;
  wire       [5:0]    _zz_when_ArraySlice_l159_206_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_206_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_206_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_206_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_206_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_206_6;
  wire       [7:0]    _zz__zz_realValue_0_206;
  wire       [7:0]    _zz__zz_realValue_0_206_1;
  wire       [7:0]    _zz_realValue_0_206_1;
  wire       [7:0]    _zz_realValue_0_206_2;
  wire       [7:0]    _zz_realValue_0_206_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_206;
  wire       [5:0]    _zz_when_ArraySlice_l166_206_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_206_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_206_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_206_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_206_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_206_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_206_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_207;
  wire       [7:0]    _zz_when_ArraySlice_l158_207_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_207_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_207_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_207;
  wire       [4:0]    _zz_when_ArraySlice_l159_207_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_207_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_207_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_207_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_207_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_207_6;
  wire       [7:0]    _zz__zz_realValue_0_207;
  wire       [7:0]    _zz__zz_realValue_0_207_1;
  wire       [7:0]    _zz_realValue_0_207_1;
  wire       [7:0]    _zz_realValue_0_207_2;
  wire       [7:0]    _zz_realValue_0_207_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_207;
  wire       [4:0]    _zz_when_ArraySlice_l166_207_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_207_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_207_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_207_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_207_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_207_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_207_7;
  wire                _zz_when_ArraySlice_l478;
  wire                _zz_when_ArraySlice_l478_1;
  wire                _zz_when_ArraySlice_l478_2;
  wire                _zz_when_ArraySlice_l478_3;
  wire                _zz_when_ArraySlice_l478_4;
  wire                _zz_when_ArraySlice_l478_5;
  wire       [7:0]    _zz_when_ArraySlice_l233;
  wire       [7:0]    _zz_when_ArraySlice_l233_1;
  wire       [3:0]    _zz_when_ArraySlice_l233_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_3;
  reg        [6:0]    _zz_when_ArraySlice_l234;
  wire       [6:0]    _zz_when_ArraySlice_l234_1;
  wire       [7:0]    _zz_when_ArraySlice_l234_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_3;
  wire       [3:0]    _zz_when_ArraySlice_l234_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_0_valid_1_1;
  wire       [3:0]    _zz__zz_outputStreamArrayData_0_valid_1_2;
  wire       [6:0]    _zz__zz_11;
  reg                 _zz_outputStreamArrayData_0_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_0_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_0_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_0_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240;
  wire       [6:0]    _zz_when_ArraySlice_l240_1;
  wire       [7:0]    _zz_when_ArraySlice_l240_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_3;
  wire       [3:0]    _zz_when_ArraySlice_l240_4;
  wire       [12:0]   _zz_when_ArraySlice_l241;
  wire       [7:0]    _zz_when_ArraySlice_l241_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_2;
  wire       [7:0]    _zz_selectReadFifo_0_16;
  wire       [7:0]    _zz_selectReadFifo_0_17;
  wire       [12:0]   _zz_when_ArraySlice_l244;
  wire       [12:0]   _zz_when_ArraySlice_l244_1;
  reg        [6:0]    _zz_when_ArraySlice_l249;
  wire       [6:0]    _zz_when_ArraySlice_l249_1;
  wire       [7:0]    _zz_when_ArraySlice_l249_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_3;
  wire       [3:0]    _zz_when_ArraySlice_l249_4;
  wire       [12:0]   _zz_when_ArraySlice_l250;
  wire       [7:0]    _zz_when_ArraySlice_l250_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_2;
  wire       [7:0]    _zz__zz_realValue1_0_24;
  wire       [7:0]    _zz__zz_realValue1_0_24_1;
  wire       [7:0]    _zz_realValue1_0_24_1;
  wire       [7:0]    _zz_realValue1_0_24_2;
  wire       [7:0]    _zz_realValue1_0_24_3;
  wire       [7:0]    _zz_when_ArraySlice_l252;
  wire       [6:0]    _zz_when_ArraySlice_l252_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_2;
  wire       [7:0]    _zz_selectReadFifo_0_18;
  wire       [7:0]    _zz_selectReadFifo_0_19;
  wire       [7:0]    _zz_selectReadFifo_0_20;
  wire       [0:0]    _zz_selectReadFifo_0_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_208;
  wire       [7:0]    _zz_when_ArraySlice_l158_208_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_208_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_208_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_208;
  wire       [7:0]    _zz_when_ArraySlice_l159_208_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_208_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_208_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_208_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_208_5;
  wire       [7:0]    _zz__zz_realValue_0_208;
  wire       [7:0]    _zz__zz_realValue_0_208_1;
  wire       [7:0]    _zz_realValue_0_208_1;
  wire       [7:0]    _zz_realValue_0_208_2;
  wire       [7:0]    _zz_realValue_0_208_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_208;
  wire       [7:0]    _zz_when_ArraySlice_l166_208_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_208_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_208_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_208_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_208_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_208_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_209;
  wire       [7:0]    _zz_when_ArraySlice_l158_209_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_209_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_209_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_209;
  wire       [6:0]    _zz_when_ArraySlice_l159_209_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_209_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_209_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_209_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_209_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_209_6;
  wire       [7:0]    _zz__zz_realValue_0_209;
  wire       [7:0]    _zz__zz_realValue_0_209_1;
  wire       [7:0]    _zz_realValue_0_209_1;
  wire       [7:0]    _zz_realValue_0_209_2;
  wire       [7:0]    _zz_realValue_0_209_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_209;
  wire       [6:0]    _zz_when_ArraySlice_l166_209_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_209_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_209_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_209_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_209_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_209_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_209_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_210;
  wire       [7:0]    _zz_when_ArraySlice_l158_210_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_210_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_210_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_210;
  wire       [6:0]    _zz_when_ArraySlice_l159_210_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_210_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_210_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_210_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_210_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_210_6;
  wire       [7:0]    _zz__zz_realValue_0_210;
  wire       [7:0]    _zz__zz_realValue_0_210_1;
  wire       [7:0]    _zz_realValue_0_210_1;
  wire       [7:0]    _zz_realValue_0_210_2;
  wire       [7:0]    _zz_realValue_0_210_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_210;
  wire       [6:0]    _zz_when_ArraySlice_l166_210_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_210_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_210_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_210_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_210_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_210_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_210_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_211;
  wire       [7:0]    _zz_when_ArraySlice_l158_211_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_211_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_211_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_211;
  wire       [6:0]    _zz_when_ArraySlice_l159_211_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_211_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_211_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_211_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_211_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_211_6;
  wire       [7:0]    _zz__zz_realValue_0_211;
  wire       [7:0]    _zz__zz_realValue_0_211_1;
  wire       [7:0]    _zz_realValue_0_211_1;
  wire       [7:0]    _zz_realValue_0_211_2;
  wire       [7:0]    _zz_realValue_0_211_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_211;
  wire       [6:0]    _zz_when_ArraySlice_l166_211_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_211_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_211_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_211_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_211_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_211_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_211_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_212;
  wire       [7:0]    _zz_when_ArraySlice_l158_212_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_212_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_212_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_212;
  wire       [6:0]    _zz_when_ArraySlice_l159_212_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_212_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_212_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_212_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_212_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_212_6;
  wire       [7:0]    _zz__zz_realValue_0_212;
  wire       [7:0]    _zz__zz_realValue_0_212_1;
  wire       [7:0]    _zz_realValue_0_212_1;
  wire       [7:0]    _zz_realValue_0_212_2;
  wire       [7:0]    _zz_realValue_0_212_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_212;
  wire       [6:0]    _zz_when_ArraySlice_l166_212_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_212_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_212_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_212_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_212_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_212_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_212_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_213;
  wire       [7:0]    _zz_when_ArraySlice_l158_213_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_213_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_213_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_213;
  wire       [5:0]    _zz_when_ArraySlice_l159_213_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_213_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_213_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_213_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_213_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_213_6;
  wire       [7:0]    _zz__zz_realValue_0_213;
  wire       [7:0]    _zz__zz_realValue_0_213_1;
  wire       [7:0]    _zz_realValue_0_213_1;
  wire       [7:0]    _zz_realValue_0_213_2;
  wire       [7:0]    _zz_realValue_0_213_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_213;
  wire       [5:0]    _zz_when_ArraySlice_l166_213_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_213_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_213_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_213_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_213_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_213_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_213_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_214;
  wire       [7:0]    _zz_when_ArraySlice_l158_214_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_214_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_214_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_214;
  wire       [5:0]    _zz_when_ArraySlice_l159_214_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_214_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_214_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_214_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_214_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_214_6;
  wire       [7:0]    _zz__zz_realValue_0_214;
  wire       [7:0]    _zz__zz_realValue_0_214_1;
  wire       [7:0]    _zz_realValue_0_214_1;
  wire       [7:0]    _zz_realValue_0_214_2;
  wire       [7:0]    _zz_realValue_0_214_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_214;
  wire       [5:0]    _zz_when_ArraySlice_l166_214_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_214_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_214_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_214_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_214_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_214_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_214_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_215;
  wire       [7:0]    _zz_when_ArraySlice_l158_215_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_215_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_215_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_215;
  wire       [4:0]    _zz_when_ArraySlice_l159_215_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_215_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_215_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_215_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_215_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_215_6;
  wire       [7:0]    _zz__zz_realValue_0_215;
  wire       [7:0]    _zz__zz_realValue_0_215_1;
  wire       [7:0]    _zz_realValue_0_215_1;
  wire       [7:0]    _zz_realValue_0_215_2;
  wire       [7:0]    _zz_realValue_0_215_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_215;
  wire       [4:0]    _zz_when_ArraySlice_l166_215_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_215_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_215_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_215_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_215_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_215_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_215_7;
  wire                _zz_when_ArraySlice_l257;
  wire                _zz_when_ArraySlice_l257_1;
  wire                _zz_when_ArraySlice_l257_2;
  wire                _zz_when_ArraySlice_l257_3;
  wire                _zz_when_ArraySlice_l257_4;
  wire                _zz_when_ArraySlice_l257_5;
  wire       [7:0]    _zz_when_ArraySlice_l260;
  wire       [7:0]    _zz_when_ArraySlice_l260_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_4;
  wire       [6:0]    _zz_when_ArraySlice_l260_5;
  wire       [7:0]    _zz_when_ArraySlice_l260_6;
  wire       [3:0]    _zz_when_ArraySlice_l260_7;
  wire       [7:0]    _zz_when_ArraySlice_l263;
  wire       [7:0]    _zz_when_ArraySlice_l263_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_3;
  wire       [6:0]    _zz_when_ArraySlice_l263_4;
  wire       [7:0]    _zz_selectReadFifo_0_22;
  wire       [7:0]    _zz_selectReadFifo_0_23;
  wire       [6:0]    _zz_selectReadFifo_0_24;
  wire       [12:0]   _zz_when_ArraySlice_l270;
  wire       [12:0]   _zz_when_ArraySlice_l270_1;
  reg        [6:0]    _zz_when_ArraySlice_l274;
  wire       [6:0]    _zz_when_ArraySlice_l274_1;
  wire       [7:0]    _zz_when_ArraySlice_l274_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_3;
  wire       [3:0]    _zz_when_ArraySlice_l274_4;
  wire       [12:0]   _zz_when_ArraySlice_l275;
  wire       [7:0]    _zz_when_ArraySlice_l275_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_3;
  wire       [0:0]    _zz_when_ArraySlice_l275_4;
  wire       [7:0]    _zz__zz_realValue1_0_25;
  wire       [7:0]    _zz__zz_realValue1_0_25_1;
  wire       [7:0]    _zz_realValue1_0_25_1;
  wire       [7:0]    _zz_realValue1_0_25_2;
  wire       [7:0]    _zz_realValue1_0_25_3;
  wire       [7:0]    _zz_when_ArraySlice_l277;
  wire       [6:0]    _zz_when_ArraySlice_l277_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_2;
  wire       [7:0]    _zz_selectReadFifo_0_25;
  wire       [7:0]    _zz_selectReadFifo_0_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_216;
  wire       [7:0]    _zz_when_ArraySlice_l158_216_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_216_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_216_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_216;
  wire       [7:0]    _zz_when_ArraySlice_l159_216_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_216_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_216_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_216_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_216_5;
  wire       [7:0]    _zz__zz_realValue_0_216;
  wire       [7:0]    _zz__zz_realValue_0_216_1;
  wire       [7:0]    _zz_realValue_0_216_1;
  wire       [7:0]    _zz_realValue_0_216_2;
  wire       [7:0]    _zz_realValue_0_216_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_216;
  wire       [7:0]    _zz_when_ArraySlice_l166_216_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_216_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_216_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_216_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_216_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_216_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_217;
  wire       [7:0]    _zz_when_ArraySlice_l158_217_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_217_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_217_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_217;
  wire       [6:0]    _zz_when_ArraySlice_l159_217_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_217_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_217_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_217_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_217_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_217_6;
  wire       [7:0]    _zz__zz_realValue_0_217;
  wire       [7:0]    _zz__zz_realValue_0_217_1;
  wire       [7:0]    _zz_realValue_0_217_1;
  wire       [7:0]    _zz_realValue_0_217_2;
  wire       [7:0]    _zz_realValue_0_217_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_217;
  wire       [6:0]    _zz_when_ArraySlice_l166_217_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_217_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_217_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_217_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_217_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_217_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_217_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_218;
  wire       [7:0]    _zz_when_ArraySlice_l158_218_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_218_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_218_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_218;
  wire       [6:0]    _zz_when_ArraySlice_l159_218_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_218_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_218_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_218_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_218_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_218_6;
  wire       [7:0]    _zz__zz_realValue_0_218;
  wire       [7:0]    _zz__zz_realValue_0_218_1;
  wire       [7:0]    _zz_realValue_0_218_1;
  wire       [7:0]    _zz_realValue_0_218_2;
  wire       [7:0]    _zz_realValue_0_218_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_218;
  wire       [6:0]    _zz_when_ArraySlice_l166_218_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_218_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_218_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_218_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_218_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_218_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_218_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_219;
  wire       [7:0]    _zz_when_ArraySlice_l158_219_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_219_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_219_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_219;
  wire       [6:0]    _zz_when_ArraySlice_l159_219_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_219_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_219_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_219_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_219_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_219_6;
  wire       [7:0]    _zz__zz_realValue_0_219;
  wire       [7:0]    _zz__zz_realValue_0_219_1;
  wire       [7:0]    _zz_realValue_0_219_1;
  wire       [7:0]    _zz_realValue_0_219_2;
  wire       [7:0]    _zz_realValue_0_219_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_219;
  wire       [6:0]    _zz_when_ArraySlice_l166_219_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_219_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_219_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_219_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_219_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_219_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_219_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_220;
  wire       [7:0]    _zz_when_ArraySlice_l158_220_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_220_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_220_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_220;
  wire       [6:0]    _zz_when_ArraySlice_l159_220_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_220_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_220_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_220_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_220_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_220_6;
  wire       [7:0]    _zz__zz_realValue_0_220;
  wire       [7:0]    _zz__zz_realValue_0_220_1;
  wire       [7:0]    _zz_realValue_0_220_1;
  wire       [7:0]    _zz_realValue_0_220_2;
  wire       [7:0]    _zz_realValue_0_220_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_220;
  wire       [6:0]    _zz_when_ArraySlice_l166_220_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_220_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_220_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_220_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_220_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_220_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_220_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_221;
  wire       [7:0]    _zz_when_ArraySlice_l158_221_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_221_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_221_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_221;
  wire       [5:0]    _zz_when_ArraySlice_l159_221_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_221_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_221_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_221_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_221_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_221_6;
  wire       [7:0]    _zz__zz_realValue_0_221;
  wire       [7:0]    _zz__zz_realValue_0_221_1;
  wire       [7:0]    _zz_realValue_0_221_1;
  wire       [7:0]    _zz_realValue_0_221_2;
  wire       [7:0]    _zz_realValue_0_221_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_221;
  wire       [5:0]    _zz_when_ArraySlice_l166_221_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_221_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_221_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_221_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_221_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_221_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_221_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_222;
  wire       [7:0]    _zz_when_ArraySlice_l158_222_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_222_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_222_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_222;
  wire       [5:0]    _zz_when_ArraySlice_l159_222_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_222_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_222_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_222_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_222_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_222_6;
  wire       [7:0]    _zz__zz_realValue_0_222;
  wire       [7:0]    _zz__zz_realValue_0_222_1;
  wire       [7:0]    _zz_realValue_0_222_1;
  wire       [7:0]    _zz_realValue_0_222_2;
  wire       [7:0]    _zz_realValue_0_222_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_222;
  wire       [5:0]    _zz_when_ArraySlice_l166_222_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_222_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_222_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_222_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_222_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_222_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_222_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_223;
  wire       [7:0]    _zz_when_ArraySlice_l158_223_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_223_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_223_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_223;
  wire       [4:0]    _zz_when_ArraySlice_l159_223_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_223_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_223_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_223_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_223_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_223_6;
  wire       [7:0]    _zz__zz_realValue_0_223;
  wire       [7:0]    _zz__zz_realValue_0_223_1;
  wire       [7:0]    _zz_realValue_0_223_1;
  wire       [7:0]    _zz_realValue_0_223_2;
  wire       [7:0]    _zz_realValue_0_223_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_223;
  wire       [4:0]    _zz_when_ArraySlice_l166_223_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_223_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_223_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_223_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_223_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_223_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_223_7;
  wire                _zz_when_ArraySlice_l282;
  wire                _zz_when_ArraySlice_l282_1;
  wire                _zz_when_ArraySlice_l282_2;
  wire                _zz_when_ArraySlice_l282_3;
  wire                _zz_when_ArraySlice_l282_4;
  wire                _zz_when_ArraySlice_l282_5;
  wire       [7:0]    _zz_when_ArraySlice_l285;
  wire       [7:0]    _zz_when_ArraySlice_l285_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_4;
  wire       [6:0]    _zz_when_ArraySlice_l285_5;
  wire       [7:0]    _zz_when_ArraySlice_l285_6;
  wire       [3:0]    _zz_when_ArraySlice_l285_7;
  wire       [7:0]    _zz_when_ArraySlice_l288;
  wire       [7:0]    _zz_when_ArraySlice_l288_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_3;
  wire       [6:0]    _zz_when_ArraySlice_l288_4;
  wire       [7:0]    _zz_selectReadFifo_0_27;
  wire       [7:0]    _zz_selectReadFifo_0_28;
  wire       [6:0]    _zz_selectReadFifo_0_29;
  wire       [12:0]   _zz_when_ArraySlice_l295;
  wire       [12:0]   _zz_when_ArraySlice_l295_1;
  wire       [12:0]   _zz_when_ArraySlice_l306;
  wire       [7:0]    _zz_when_ArraySlice_l306_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_2;
  wire       [7:0]    _zz__zz_realValue1_0_26;
  wire       [7:0]    _zz__zz_realValue1_0_26_1;
  wire       [7:0]    _zz_realValue1_0_26_1;
  wire       [7:0]    _zz_realValue1_0_26_2;
  wire       [7:0]    _zz_realValue1_0_26_3;
  wire       [7:0]    _zz_when_ArraySlice_l307;
  wire       [6:0]    _zz_when_ArraySlice_l307_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_2;
  wire       [7:0]    _zz_selectReadFifo_0_30;
  wire       [7:0]    _zz_selectReadFifo_0_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_224;
  wire       [7:0]    _zz_when_ArraySlice_l158_224_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_224_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_224_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_224;
  wire       [7:0]    _zz_when_ArraySlice_l159_224_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_224_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_224_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_224_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_224_5;
  wire       [7:0]    _zz__zz_realValue_0_224;
  wire       [7:0]    _zz__zz_realValue_0_224_1;
  wire       [7:0]    _zz_realValue_0_224_1;
  wire       [7:0]    _zz_realValue_0_224_2;
  wire       [7:0]    _zz_realValue_0_224_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_224;
  wire       [7:0]    _zz_when_ArraySlice_l166_224_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_224_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_224_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_224_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_224_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_224_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_225;
  wire       [7:0]    _zz_when_ArraySlice_l158_225_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_225_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_225_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_225;
  wire       [6:0]    _zz_when_ArraySlice_l159_225_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_225_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_225_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_225_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_225_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_225_6;
  wire       [7:0]    _zz__zz_realValue_0_225;
  wire       [7:0]    _zz__zz_realValue_0_225_1;
  wire       [7:0]    _zz_realValue_0_225_1;
  wire       [7:0]    _zz_realValue_0_225_2;
  wire       [7:0]    _zz_realValue_0_225_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_225;
  wire       [6:0]    _zz_when_ArraySlice_l166_225_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_225_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_225_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_225_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_225_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_225_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_225_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_226;
  wire       [7:0]    _zz_when_ArraySlice_l158_226_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_226_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_226_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_226;
  wire       [6:0]    _zz_when_ArraySlice_l159_226_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_226_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_226_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_226_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_226_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_226_6;
  wire       [7:0]    _zz__zz_realValue_0_226;
  wire       [7:0]    _zz__zz_realValue_0_226_1;
  wire       [7:0]    _zz_realValue_0_226_1;
  wire       [7:0]    _zz_realValue_0_226_2;
  wire       [7:0]    _zz_realValue_0_226_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_226;
  wire       [6:0]    _zz_when_ArraySlice_l166_226_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_226_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_226_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_226_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_226_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_226_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_226_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_227;
  wire       [7:0]    _zz_when_ArraySlice_l158_227_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_227_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_227_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_227;
  wire       [6:0]    _zz_when_ArraySlice_l159_227_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_227_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_227_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_227_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_227_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_227_6;
  wire       [7:0]    _zz__zz_realValue_0_227;
  wire       [7:0]    _zz__zz_realValue_0_227_1;
  wire       [7:0]    _zz_realValue_0_227_1;
  wire       [7:0]    _zz_realValue_0_227_2;
  wire       [7:0]    _zz_realValue_0_227_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_227;
  wire       [6:0]    _zz_when_ArraySlice_l166_227_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_227_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_227_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_227_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_227_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_227_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_227_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_228;
  wire       [7:0]    _zz_when_ArraySlice_l158_228_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_228_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_228_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_228;
  wire       [6:0]    _zz_when_ArraySlice_l159_228_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_228_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_228_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_228_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_228_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_228_6;
  wire       [7:0]    _zz__zz_realValue_0_228;
  wire       [7:0]    _zz__zz_realValue_0_228_1;
  wire       [7:0]    _zz_realValue_0_228_1;
  wire       [7:0]    _zz_realValue_0_228_2;
  wire       [7:0]    _zz_realValue_0_228_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_228;
  wire       [6:0]    _zz_when_ArraySlice_l166_228_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_228_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_228_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_228_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_228_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_228_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_228_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_229;
  wire       [7:0]    _zz_when_ArraySlice_l158_229_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_229_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_229_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_229;
  wire       [5:0]    _zz_when_ArraySlice_l159_229_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_229_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_229_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_229_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_229_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_229_6;
  wire       [7:0]    _zz__zz_realValue_0_229;
  wire       [7:0]    _zz__zz_realValue_0_229_1;
  wire       [7:0]    _zz_realValue_0_229_1;
  wire       [7:0]    _zz_realValue_0_229_2;
  wire       [7:0]    _zz_realValue_0_229_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_229;
  wire       [5:0]    _zz_when_ArraySlice_l166_229_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_229_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_229_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_229_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_229_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_229_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_229_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_230;
  wire       [7:0]    _zz_when_ArraySlice_l158_230_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_230_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_230_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_230;
  wire       [5:0]    _zz_when_ArraySlice_l159_230_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_230_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_230_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_230_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_230_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_230_6;
  wire       [7:0]    _zz__zz_realValue_0_230;
  wire       [7:0]    _zz__zz_realValue_0_230_1;
  wire       [7:0]    _zz_realValue_0_230_1;
  wire       [7:0]    _zz_realValue_0_230_2;
  wire       [7:0]    _zz_realValue_0_230_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_230;
  wire       [5:0]    _zz_when_ArraySlice_l166_230_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_230_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_230_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_230_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_230_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_230_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_230_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_231;
  wire       [7:0]    _zz_when_ArraySlice_l158_231_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_231_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_231_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_231;
  wire       [4:0]    _zz_when_ArraySlice_l159_231_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_231_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_231_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_231_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_231_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_231_6;
  wire       [7:0]    _zz__zz_realValue_0_231;
  wire       [7:0]    _zz__zz_realValue_0_231_1;
  wire       [7:0]    _zz_realValue_0_231_1;
  wire       [7:0]    _zz_realValue_0_231_2;
  wire       [7:0]    _zz_realValue_0_231_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_231;
  wire       [4:0]    _zz_when_ArraySlice_l166_231_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_231_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_231_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_231_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_231_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_231_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_231_7;
  wire                _zz_when_ArraySlice_l314;
  wire                _zz_when_ArraySlice_l314_1;
  wire                _zz_when_ArraySlice_l314_2;
  wire                _zz_when_ArraySlice_l314_3;
  wire                _zz_when_ArraySlice_l314_4;
  wire                _zz_when_ArraySlice_l314_5;
  wire       [12:0]   _zz_when_ArraySlice_l318;
  wire       [12:0]   _zz_when_ArraySlice_l318_1;
  wire       [7:0]    _zz_when_ArraySlice_l304;
  wire       [7:0]    _zz_when_ArraySlice_l304_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_2;
  wire       [3:0]    _zz_when_ArraySlice_l304_3;
  wire       [12:0]   _zz_when_ArraySlice_l325;
  wire       [7:0]    _zz_when_ArraySlice_l325_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l233_1_2;
  wire       [4:0]    _zz_when_ArraySlice_l233_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l233_1_4;
  reg        [6:0]    _zz_when_ArraySlice_l234_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l234_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l234_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l234_1_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_1_valid_1_1;
  wire       [4:0]    _zz__zz_outputStreamArrayData_1_valid_1_2;
  wire       [6:0]    _zz__zz_12;
  reg                 _zz_outputStreamArrayData_1_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_1_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_1_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_1_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l240_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l240_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l240_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l241_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l241_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_16;
  wire       [7:0]    _zz_selectReadFifo_1_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l244_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l249_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l249_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l249_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l249_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l250_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l250_1_3;
  wire       [7:0]    _zz__zz_realValue1_0_27;
  wire       [7:0]    _zz__zz_realValue1_0_27_1;
  wire       [7:0]    _zz_realValue1_0_27_1;
  wire       [7:0]    _zz_realValue1_0_27_2;
  wire       [7:0]    _zz_realValue1_0_27_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l252_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l252_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_18;
  wire       [7:0]    _zz_selectReadFifo_1_19;
  wire       [7:0]    _zz_selectReadFifo_1_20;
  wire       [0:0]    _zz_selectReadFifo_1_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_232;
  wire       [7:0]    _zz_when_ArraySlice_l158_232_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_232_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_232_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_232;
  wire       [7:0]    _zz_when_ArraySlice_l159_232_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_232_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_232_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_232_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_232_5;
  wire       [7:0]    _zz__zz_realValue_0_232;
  wire       [7:0]    _zz__zz_realValue_0_232_1;
  wire       [7:0]    _zz_realValue_0_232_1;
  wire       [7:0]    _zz_realValue_0_232_2;
  wire       [7:0]    _zz_realValue_0_232_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_232;
  wire       [7:0]    _zz_when_ArraySlice_l166_232_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_232_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_232_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_232_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_232_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_232_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_233;
  wire       [7:0]    _zz_when_ArraySlice_l158_233_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_233_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_233_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_233;
  wire       [6:0]    _zz_when_ArraySlice_l159_233_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_233_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_233_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_233_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_233_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_233_6;
  wire       [7:0]    _zz__zz_realValue_0_233;
  wire       [7:0]    _zz__zz_realValue_0_233_1;
  wire       [7:0]    _zz_realValue_0_233_1;
  wire       [7:0]    _zz_realValue_0_233_2;
  wire       [7:0]    _zz_realValue_0_233_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_233;
  wire       [6:0]    _zz_when_ArraySlice_l166_233_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_233_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_233_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_233_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_233_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_233_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_233_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_234;
  wire       [7:0]    _zz_when_ArraySlice_l158_234_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_234_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_234_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_234;
  wire       [6:0]    _zz_when_ArraySlice_l159_234_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_234_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_234_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_234_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_234_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_234_6;
  wire       [7:0]    _zz__zz_realValue_0_234;
  wire       [7:0]    _zz__zz_realValue_0_234_1;
  wire       [7:0]    _zz_realValue_0_234_1;
  wire       [7:0]    _zz_realValue_0_234_2;
  wire       [7:0]    _zz_realValue_0_234_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_234;
  wire       [6:0]    _zz_when_ArraySlice_l166_234_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_234_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_234_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_234_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_234_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_234_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_234_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_235;
  wire       [7:0]    _zz_when_ArraySlice_l158_235_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_235_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_235_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_235;
  wire       [6:0]    _zz_when_ArraySlice_l159_235_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_235_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_235_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_235_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_235_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_235_6;
  wire       [7:0]    _zz__zz_realValue_0_235;
  wire       [7:0]    _zz__zz_realValue_0_235_1;
  wire       [7:0]    _zz_realValue_0_235_1;
  wire       [7:0]    _zz_realValue_0_235_2;
  wire       [7:0]    _zz_realValue_0_235_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_235;
  wire       [6:0]    _zz_when_ArraySlice_l166_235_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_235_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_235_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_235_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_235_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_235_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_235_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_236;
  wire       [7:0]    _zz_when_ArraySlice_l158_236_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_236_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_236_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_236;
  wire       [6:0]    _zz_when_ArraySlice_l159_236_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_236_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_236_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_236_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_236_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_236_6;
  wire       [7:0]    _zz__zz_realValue_0_236;
  wire       [7:0]    _zz__zz_realValue_0_236_1;
  wire       [7:0]    _zz_realValue_0_236_1;
  wire       [7:0]    _zz_realValue_0_236_2;
  wire       [7:0]    _zz_realValue_0_236_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_236;
  wire       [6:0]    _zz_when_ArraySlice_l166_236_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_236_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_236_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_236_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_236_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_236_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_236_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_237;
  wire       [7:0]    _zz_when_ArraySlice_l158_237_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_237_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_237_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_237;
  wire       [5:0]    _zz_when_ArraySlice_l159_237_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_237_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_237_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_237_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_237_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_237_6;
  wire       [7:0]    _zz__zz_realValue_0_237;
  wire       [7:0]    _zz__zz_realValue_0_237_1;
  wire       [7:0]    _zz_realValue_0_237_1;
  wire       [7:0]    _zz_realValue_0_237_2;
  wire       [7:0]    _zz_realValue_0_237_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_237;
  wire       [5:0]    _zz_when_ArraySlice_l166_237_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_237_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_237_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_237_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_237_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_237_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_237_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_238;
  wire       [7:0]    _zz_when_ArraySlice_l158_238_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_238_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_238_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_238;
  wire       [5:0]    _zz_when_ArraySlice_l159_238_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_238_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_238_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_238_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_238_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_238_6;
  wire       [7:0]    _zz__zz_realValue_0_238;
  wire       [7:0]    _zz__zz_realValue_0_238_1;
  wire       [7:0]    _zz_realValue_0_238_1;
  wire       [7:0]    _zz_realValue_0_238_2;
  wire       [7:0]    _zz_realValue_0_238_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_238;
  wire       [5:0]    _zz_when_ArraySlice_l166_238_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_238_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_238_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_238_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_238_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_238_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_238_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_239;
  wire       [7:0]    _zz_when_ArraySlice_l158_239_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_239_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_239_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_239;
  wire       [4:0]    _zz_when_ArraySlice_l159_239_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_239_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_239_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_239_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_239_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_239_6;
  wire       [7:0]    _zz__zz_realValue_0_239;
  wire       [7:0]    _zz__zz_realValue_0_239_1;
  wire       [7:0]    _zz_realValue_0_239_1;
  wire       [7:0]    _zz_realValue_0_239_2;
  wire       [7:0]    _zz_realValue_0_239_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_239;
  wire       [4:0]    _zz_when_ArraySlice_l166_239_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_239_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_239_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_239_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_239_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_239_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_239_7;
  wire                _zz_when_ArraySlice_l257_1_1;
  wire                _zz_when_ArraySlice_l257_1_2;
  wire                _zz_when_ArraySlice_l257_1_3;
  wire                _zz_when_ArraySlice_l257_1_4;
  wire                _zz_when_ArraySlice_l257_1_5;
  wire                _zz_when_ArraySlice_l257_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_1_7;
  wire       [4:0]    _zz_when_ArraySlice_l260_1_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l263_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l263_1_5;
  wire       [7:0]    _zz_selectReadFifo_1_22;
  wire       [7:0]    _zz_selectReadFifo_1_23;
  wire       [6:0]    _zz_selectReadFifo_1_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l270_1_2;
  reg        [6:0]    _zz_when_ArraySlice_l274_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l274_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l274_1_4;
  wire       [4:0]    _zz_when_ArraySlice_l274_1_5;
  wire       [12:0]   _zz_when_ArraySlice_l275_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l275_1_4;
  wire       [0:0]    _zz_when_ArraySlice_l275_1_5;
  wire       [7:0]    _zz__zz_realValue1_0_28;
  wire       [7:0]    _zz__zz_realValue1_0_28_1;
  wire       [7:0]    _zz_realValue1_0_28_1;
  wire       [7:0]    _zz_realValue1_0_28_2;
  wire       [7:0]    _zz_realValue1_0_28_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l277_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l277_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_25;
  wire       [7:0]    _zz_selectReadFifo_1_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_240;
  wire       [7:0]    _zz_when_ArraySlice_l158_240_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_240_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_240_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_240;
  wire       [7:0]    _zz_when_ArraySlice_l159_240_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_240_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_240_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_240_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_240_5;
  wire       [7:0]    _zz__zz_realValue_0_240;
  wire       [7:0]    _zz__zz_realValue_0_240_1;
  wire       [7:0]    _zz_realValue_0_240_1;
  wire       [7:0]    _zz_realValue_0_240_2;
  wire       [7:0]    _zz_realValue_0_240_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_240;
  wire       [7:0]    _zz_when_ArraySlice_l166_240_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_240_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_240_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_240_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_240_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_240_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_241;
  wire       [7:0]    _zz_when_ArraySlice_l158_241_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_241_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_241_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_241;
  wire       [6:0]    _zz_when_ArraySlice_l159_241_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_241_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_241_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_241_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_241_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_241_6;
  wire       [7:0]    _zz__zz_realValue_0_241;
  wire       [7:0]    _zz__zz_realValue_0_241_1;
  wire       [7:0]    _zz_realValue_0_241_1;
  wire       [7:0]    _zz_realValue_0_241_2;
  wire       [7:0]    _zz_realValue_0_241_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_241;
  wire       [6:0]    _zz_when_ArraySlice_l166_241_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_241_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_241_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_241_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_241_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_241_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_241_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_242;
  wire       [7:0]    _zz_when_ArraySlice_l158_242_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_242_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_242_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_242;
  wire       [6:0]    _zz_when_ArraySlice_l159_242_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_242_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_242_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_242_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_242_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_242_6;
  wire       [7:0]    _zz__zz_realValue_0_242;
  wire       [7:0]    _zz__zz_realValue_0_242_1;
  wire       [7:0]    _zz_realValue_0_242_1;
  wire       [7:0]    _zz_realValue_0_242_2;
  wire       [7:0]    _zz_realValue_0_242_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_242;
  wire       [6:0]    _zz_when_ArraySlice_l166_242_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_242_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_242_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_242_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_242_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_242_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_242_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_243;
  wire       [7:0]    _zz_when_ArraySlice_l158_243_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_243_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_243_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_243;
  wire       [6:0]    _zz_when_ArraySlice_l159_243_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_243_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_243_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_243_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_243_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_243_6;
  wire       [7:0]    _zz__zz_realValue_0_243;
  wire       [7:0]    _zz__zz_realValue_0_243_1;
  wire       [7:0]    _zz_realValue_0_243_1;
  wire       [7:0]    _zz_realValue_0_243_2;
  wire       [7:0]    _zz_realValue_0_243_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_243;
  wire       [6:0]    _zz_when_ArraySlice_l166_243_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_243_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_243_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_243_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_243_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_243_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_243_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_244;
  wire       [7:0]    _zz_when_ArraySlice_l158_244_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_244_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_244_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_244;
  wire       [6:0]    _zz_when_ArraySlice_l159_244_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_244_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_244_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_244_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_244_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_244_6;
  wire       [7:0]    _zz__zz_realValue_0_244;
  wire       [7:0]    _zz__zz_realValue_0_244_1;
  wire       [7:0]    _zz_realValue_0_244_1;
  wire       [7:0]    _zz_realValue_0_244_2;
  wire       [7:0]    _zz_realValue_0_244_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_244;
  wire       [6:0]    _zz_when_ArraySlice_l166_244_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_244_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_244_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_244_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_244_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_244_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_244_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_245;
  wire       [7:0]    _zz_when_ArraySlice_l158_245_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_245_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_245_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_245;
  wire       [5:0]    _zz_when_ArraySlice_l159_245_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_245_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_245_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_245_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_245_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_245_6;
  wire       [7:0]    _zz__zz_realValue_0_245;
  wire       [7:0]    _zz__zz_realValue_0_245_1;
  wire       [7:0]    _zz_realValue_0_245_1;
  wire       [7:0]    _zz_realValue_0_245_2;
  wire       [7:0]    _zz_realValue_0_245_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_245;
  wire       [5:0]    _zz_when_ArraySlice_l166_245_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_245_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_245_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_245_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_245_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_245_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_245_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_246;
  wire       [7:0]    _zz_when_ArraySlice_l158_246_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_246_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_246_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_246;
  wire       [5:0]    _zz_when_ArraySlice_l159_246_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_246_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_246_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_246_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_246_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_246_6;
  wire       [7:0]    _zz__zz_realValue_0_246;
  wire       [7:0]    _zz__zz_realValue_0_246_1;
  wire       [7:0]    _zz_realValue_0_246_1;
  wire       [7:0]    _zz_realValue_0_246_2;
  wire       [7:0]    _zz_realValue_0_246_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_246;
  wire       [5:0]    _zz_when_ArraySlice_l166_246_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_246_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_246_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_246_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_246_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_246_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_246_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_247;
  wire       [7:0]    _zz_when_ArraySlice_l158_247_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_247_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_247_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_247;
  wire       [4:0]    _zz_when_ArraySlice_l159_247_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_247_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_247_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_247_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_247_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_247_6;
  wire       [7:0]    _zz__zz_realValue_0_247;
  wire       [7:0]    _zz__zz_realValue_0_247_1;
  wire       [7:0]    _zz_realValue_0_247_1;
  wire       [7:0]    _zz_realValue_0_247_2;
  wire       [7:0]    _zz_realValue_0_247_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_247;
  wire       [4:0]    _zz_when_ArraySlice_l166_247_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_247_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_247_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_247_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_247_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_247_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_247_7;
  wire                _zz_when_ArraySlice_l282_1_1;
  wire                _zz_when_ArraySlice_l282_1_2;
  wire                _zz_when_ArraySlice_l282_1_3;
  wire                _zz_when_ArraySlice_l282_1_4;
  wire                _zz_when_ArraySlice_l282_1_5;
  wire                _zz_when_ArraySlice_l282_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_1_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_1_7;
  wire       [4:0]    _zz_when_ArraySlice_l285_1_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l288_1_4;
  wire       [6:0]    _zz_when_ArraySlice_l288_1_5;
  wire       [7:0]    _zz_selectReadFifo_1_27;
  wire       [7:0]    _zz_selectReadFifo_1_28;
  wire       [6:0]    _zz_selectReadFifo_1_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l295_1_2;
  wire       [12:0]   _zz_when_ArraySlice_l306_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l306_1_3;
  wire       [7:0]    _zz__zz_realValue1_0_29;
  wire       [7:0]    _zz__zz_realValue1_0_29_1;
  wire       [7:0]    _zz_realValue1_0_29_1;
  wire       [7:0]    _zz_realValue1_0_29_2;
  wire       [7:0]    _zz_realValue1_0_29_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_1_1;
  wire       [6:0]    _zz_when_ArraySlice_l307_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l307_1_3;
  wire       [7:0]    _zz_selectReadFifo_1_30;
  wire       [7:0]    _zz_selectReadFifo_1_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_248;
  wire       [7:0]    _zz_when_ArraySlice_l158_248_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_248_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_248_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_248;
  wire       [7:0]    _zz_when_ArraySlice_l159_248_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_248_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_248_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_248_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_248_5;
  wire       [7:0]    _zz__zz_realValue_0_248;
  wire       [7:0]    _zz__zz_realValue_0_248_1;
  wire       [7:0]    _zz_realValue_0_248_1;
  wire       [7:0]    _zz_realValue_0_248_2;
  wire       [7:0]    _zz_realValue_0_248_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_248;
  wire       [7:0]    _zz_when_ArraySlice_l166_248_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_248_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_248_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_248_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_248_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_248_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_249;
  wire       [7:0]    _zz_when_ArraySlice_l158_249_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_249_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_249_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_249;
  wire       [6:0]    _zz_when_ArraySlice_l159_249_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_249_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_249_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_249_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_249_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_249_6;
  wire       [7:0]    _zz__zz_realValue_0_249;
  wire       [7:0]    _zz__zz_realValue_0_249_1;
  wire       [7:0]    _zz_realValue_0_249_1;
  wire       [7:0]    _zz_realValue_0_249_2;
  wire       [7:0]    _zz_realValue_0_249_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_249;
  wire       [6:0]    _zz_when_ArraySlice_l166_249_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_249_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_249_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_249_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_249_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_249_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_249_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_250;
  wire       [7:0]    _zz_when_ArraySlice_l158_250_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_250_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_250_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_250;
  wire       [6:0]    _zz_when_ArraySlice_l159_250_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_250_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_250_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_250_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_250_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_250_6;
  wire       [7:0]    _zz__zz_realValue_0_250;
  wire       [7:0]    _zz__zz_realValue_0_250_1;
  wire       [7:0]    _zz_realValue_0_250_1;
  wire       [7:0]    _zz_realValue_0_250_2;
  wire       [7:0]    _zz_realValue_0_250_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_250;
  wire       [6:0]    _zz_when_ArraySlice_l166_250_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_250_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_250_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_250_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_250_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_250_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_250_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_251;
  wire       [7:0]    _zz_when_ArraySlice_l158_251_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_251_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_251_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_251;
  wire       [6:0]    _zz_when_ArraySlice_l159_251_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_251_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_251_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_251_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_251_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_251_6;
  wire       [7:0]    _zz__zz_realValue_0_251;
  wire       [7:0]    _zz__zz_realValue_0_251_1;
  wire       [7:0]    _zz_realValue_0_251_1;
  wire       [7:0]    _zz_realValue_0_251_2;
  wire       [7:0]    _zz_realValue_0_251_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_251;
  wire       [6:0]    _zz_when_ArraySlice_l166_251_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_251_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_251_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_251_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_251_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_251_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_251_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_252;
  wire       [7:0]    _zz_when_ArraySlice_l158_252_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_252_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_252_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_252;
  wire       [6:0]    _zz_when_ArraySlice_l159_252_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_252_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_252_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_252_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_252_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_252_6;
  wire       [7:0]    _zz__zz_realValue_0_252;
  wire       [7:0]    _zz__zz_realValue_0_252_1;
  wire       [7:0]    _zz_realValue_0_252_1;
  wire       [7:0]    _zz_realValue_0_252_2;
  wire       [7:0]    _zz_realValue_0_252_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_252;
  wire       [6:0]    _zz_when_ArraySlice_l166_252_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_252_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_252_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_252_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_252_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_252_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_252_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_253;
  wire       [7:0]    _zz_when_ArraySlice_l158_253_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_253_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_253_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_253;
  wire       [5:0]    _zz_when_ArraySlice_l159_253_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_253_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_253_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_253_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_253_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_253_6;
  wire       [7:0]    _zz__zz_realValue_0_253;
  wire       [7:0]    _zz__zz_realValue_0_253_1;
  wire       [7:0]    _zz_realValue_0_253_1;
  wire       [7:0]    _zz_realValue_0_253_2;
  wire       [7:0]    _zz_realValue_0_253_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_253;
  wire       [5:0]    _zz_when_ArraySlice_l166_253_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_253_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_253_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_253_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_253_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_253_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_253_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_254;
  wire       [7:0]    _zz_when_ArraySlice_l158_254_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_254_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_254_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_254;
  wire       [5:0]    _zz_when_ArraySlice_l159_254_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_254_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_254_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_254_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_254_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_254_6;
  wire       [7:0]    _zz__zz_realValue_0_254;
  wire       [7:0]    _zz__zz_realValue_0_254_1;
  wire       [7:0]    _zz_realValue_0_254_1;
  wire       [7:0]    _zz_realValue_0_254_2;
  wire       [7:0]    _zz_realValue_0_254_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_254;
  wire       [5:0]    _zz_when_ArraySlice_l166_254_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_254_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_254_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_254_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_254_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_254_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_254_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_255;
  wire       [7:0]    _zz_when_ArraySlice_l158_255_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_255_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_255_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_255;
  wire       [4:0]    _zz_when_ArraySlice_l159_255_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_255_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_255_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_255_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_255_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_255_6;
  wire       [7:0]    _zz__zz_realValue_0_255;
  wire       [7:0]    _zz__zz_realValue_0_255_1;
  wire       [7:0]    _zz_realValue_0_255_1;
  wire       [7:0]    _zz_realValue_0_255_2;
  wire       [7:0]    _zz_realValue_0_255_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_255;
  wire       [4:0]    _zz_when_ArraySlice_l166_255_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_255_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_255_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_255_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_255_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_255_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_255_7;
  wire                _zz_when_ArraySlice_l314_1_1;
  wire                _zz_when_ArraySlice_l314_1_2;
  wire                _zz_when_ArraySlice_l314_1_3;
  wire                _zz_when_ArraySlice_l314_1_4;
  wire                _zz_when_ArraySlice_l314_1_5;
  wire                _zz_when_ArraySlice_l314_1_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_1_1;
  wire       [12:0]   _zz_when_ArraySlice_l318_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l304_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l304_1_3;
  wire       [4:0]    _zz_when_ArraySlice_l304_1_4;
  wire       [12:0]   _zz_when_ArraySlice_l325_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l325_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l233_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l233_2_2;
  wire       [5:0]    _zz_when_ArraySlice_l233_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l233_2_4;
  reg        [6:0]    _zz_when_ArraySlice_l234_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l234_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l234_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l234_2_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_2_valid_1_1;
  wire       [5:0]    _zz__zz_outputStreamArrayData_2_valid_1_2;
  wire       [6:0]    _zz__zz_13;
  reg                 _zz_outputStreamArrayData_2_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_2_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_2_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_2_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l240_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l240_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l241_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l241_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_16;
  wire       [7:0]    _zz_selectReadFifo_2_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_2;
  wire       [12:0]   _zz_when_ArraySlice_l244_2_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l249_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l249_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l249_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l250_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l250_2_3;
  wire       [7:0]    _zz__zz_realValue1_0_30;
  wire       [7:0]    _zz__zz_realValue1_0_30_1;
  wire       [7:0]    _zz_realValue1_0_30_1;
  wire       [7:0]    _zz_realValue1_0_30_2;
  wire       [7:0]    _zz_realValue1_0_30_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l252_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l252_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_18;
  wire       [7:0]    _zz_selectReadFifo_2_19;
  wire       [7:0]    _zz_selectReadFifo_2_20;
  wire       [0:0]    _zz_selectReadFifo_2_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_256;
  wire       [7:0]    _zz_when_ArraySlice_l158_256_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_256_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_256_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_256;
  wire       [7:0]    _zz_when_ArraySlice_l159_256_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_256_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_256_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_256_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_256_5;
  wire       [7:0]    _zz__zz_realValue_0_256;
  wire       [7:0]    _zz__zz_realValue_0_256_1;
  wire       [7:0]    _zz_realValue_0_256_1;
  wire       [7:0]    _zz_realValue_0_256_2;
  wire       [7:0]    _zz_realValue_0_256_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_256;
  wire       [7:0]    _zz_when_ArraySlice_l166_256_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_256_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_256_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_256_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_256_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_256_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_257;
  wire       [7:0]    _zz_when_ArraySlice_l158_257_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_257_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_257_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_257;
  wire       [6:0]    _zz_when_ArraySlice_l159_257_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_257_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_257_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_257_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_257_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_257_6;
  wire       [7:0]    _zz__zz_realValue_0_257;
  wire       [7:0]    _zz__zz_realValue_0_257_1;
  wire       [7:0]    _zz_realValue_0_257_1;
  wire       [7:0]    _zz_realValue_0_257_2;
  wire       [7:0]    _zz_realValue_0_257_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_257;
  wire       [6:0]    _zz_when_ArraySlice_l166_257_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_257_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_257_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_257_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_257_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_257_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_257_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_258;
  wire       [7:0]    _zz_when_ArraySlice_l158_258_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_258_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_258_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_258;
  wire       [6:0]    _zz_when_ArraySlice_l159_258_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_258_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_258_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_258_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_258_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_258_6;
  wire       [7:0]    _zz__zz_realValue_0_258;
  wire       [7:0]    _zz__zz_realValue_0_258_1;
  wire       [7:0]    _zz_realValue_0_258_1;
  wire       [7:0]    _zz_realValue_0_258_2;
  wire       [7:0]    _zz_realValue_0_258_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_258;
  wire       [6:0]    _zz_when_ArraySlice_l166_258_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_258_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_258_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_258_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_258_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_258_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_258_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_259;
  wire       [7:0]    _zz_when_ArraySlice_l158_259_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_259_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_259_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_259;
  wire       [6:0]    _zz_when_ArraySlice_l159_259_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_259_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_259_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_259_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_259_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_259_6;
  wire       [7:0]    _zz__zz_realValue_0_259;
  wire       [7:0]    _zz__zz_realValue_0_259_1;
  wire       [7:0]    _zz_realValue_0_259_1;
  wire       [7:0]    _zz_realValue_0_259_2;
  wire       [7:0]    _zz_realValue_0_259_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_259;
  wire       [6:0]    _zz_when_ArraySlice_l166_259_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_259_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_259_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_259_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_259_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_259_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_259_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_260;
  wire       [7:0]    _zz_when_ArraySlice_l158_260_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_260_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_260_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_260;
  wire       [6:0]    _zz_when_ArraySlice_l159_260_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_260_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_260_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_260_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_260_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_260_6;
  wire       [7:0]    _zz__zz_realValue_0_260;
  wire       [7:0]    _zz__zz_realValue_0_260_1;
  wire       [7:0]    _zz_realValue_0_260_1;
  wire       [7:0]    _zz_realValue_0_260_2;
  wire       [7:0]    _zz_realValue_0_260_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_260;
  wire       [6:0]    _zz_when_ArraySlice_l166_260_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_260_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_260_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_260_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_260_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_260_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_260_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_261;
  wire       [7:0]    _zz_when_ArraySlice_l158_261_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_261_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_261_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_261;
  wire       [5:0]    _zz_when_ArraySlice_l159_261_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_261_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_261_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_261_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_261_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_261_6;
  wire       [7:0]    _zz__zz_realValue_0_261;
  wire       [7:0]    _zz__zz_realValue_0_261_1;
  wire       [7:0]    _zz_realValue_0_261_1;
  wire       [7:0]    _zz_realValue_0_261_2;
  wire       [7:0]    _zz_realValue_0_261_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_261;
  wire       [5:0]    _zz_when_ArraySlice_l166_261_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_261_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_261_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_261_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_261_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_261_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_261_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_262;
  wire       [7:0]    _zz_when_ArraySlice_l158_262_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_262_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_262_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_262;
  wire       [5:0]    _zz_when_ArraySlice_l159_262_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_262_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_262_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_262_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_262_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_262_6;
  wire       [7:0]    _zz__zz_realValue_0_262;
  wire       [7:0]    _zz__zz_realValue_0_262_1;
  wire       [7:0]    _zz_realValue_0_262_1;
  wire       [7:0]    _zz_realValue_0_262_2;
  wire       [7:0]    _zz_realValue_0_262_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_262;
  wire       [5:0]    _zz_when_ArraySlice_l166_262_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_262_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_262_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_262_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_262_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_262_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_262_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_263;
  wire       [7:0]    _zz_when_ArraySlice_l158_263_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_263_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_263_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_263;
  wire       [4:0]    _zz_when_ArraySlice_l159_263_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_263_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_263_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_263_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_263_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_263_6;
  wire       [7:0]    _zz__zz_realValue_0_263;
  wire       [7:0]    _zz__zz_realValue_0_263_1;
  wire       [7:0]    _zz_realValue_0_263_1;
  wire       [7:0]    _zz_realValue_0_263_2;
  wire       [7:0]    _zz_realValue_0_263_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_263;
  wire       [4:0]    _zz_when_ArraySlice_l166_263_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_263_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_263_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_263_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_263_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_263_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_263_7;
  wire                _zz_when_ArraySlice_l257_2_1;
  wire                _zz_when_ArraySlice_l257_2_2;
  wire                _zz_when_ArraySlice_l257_2_3;
  wire                _zz_when_ArraySlice_l257_2_4;
  wire                _zz_when_ArraySlice_l257_2_5;
  wire                _zz_when_ArraySlice_l257_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_2_7;
  wire       [5:0]    _zz_when_ArraySlice_l260_2_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l263_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l263_2_5;
  wire       [7:0]    _zz_selectReadFifo_2_22;
  wire       [7:0]    _zz_selectReadFifo_2_23;
  wire       [6:0]    _zz_selectReadFifo_2_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_2;
  wire       [12:0]   _zz_when_ArraySlice_l270_2_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l274_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l274_2_4;
  wire       [5:0]    _zz_when_ArraySlice_l274_2_5;
  wire       [12:0]   _zz_when_ArraySlice_l275_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l275_2_4;
  wire       [0:0]    _zz_when_ArraySlice_l275_2_5;
  wire       [7:0]    _zz__zz_realValue1_0_31;
  wire       [7:0]    _zz__zz_realValue1_0_31_1;
  wire       [7:0]    _zz_realValue1_0_31_1;
  wire       [7:0]    _zz_realValue1_0_31_2;
  wire       [7:0]    _zz_realValue1_0_31_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l277_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l277_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_25;
  wire       [7:0]    _zz_selectReadFifo_2_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_264;
  wire       [7:0]    _zz_when_ArraySlice_l158_264_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_264_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_264_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_264;
  wire       [7:0]    _zz_when_ArraySlice_l159_264_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_264_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_264_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_264_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_264_5;
  wire       [7:0]    _zz__zz_realValue_0_264;
  wire       [7:0]    _zz__zz_realValue_0_264_1;
  wire       [7:0]    _zz_realValue_0_264_1;
  wire       [7:0]    _zz_realValue_0_264_2;
  wire       [7:0]    _zz_realValue_0_264_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_264;
  wire       [7:0]    _zz_when_ArraySlice_l166_264_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_264_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_264_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_264_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_264_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_264_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_265;
  wire       [7:0]    _zz_when_ArraySlice_l158_265_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_265_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_265_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_265;
  wire       [6:0]    _zz_when_ArraySlice_l159_265_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_265_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_265_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_265_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_265_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_265_6;
  wire       [7:0]    _zz__zz_realValue_0_265;
  wire       [7:0]    _zz__zz_realValue_0_265_1;
  wire       [7:0]    _zz_realValue_0_265_1;
  wire       [7:0]    _zz_realValue_0_265_2;
  wire       [7:0]    _zz_realValue_0_265_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_265;
  wire       [6:0]    _zz_when_ArraySlice_l166_265_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_265_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_265_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_265_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_265_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_265_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_265_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_266;
  wire       [7:0]    _zz_when_ArraySlice_l158_266_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_266_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_266_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_266;
  wire       [6:0]    _zz_when_ArraySlice_l159_266_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_266_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_266_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_266_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_266_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_266_6;
  wire       [7:0]    _zz__zz_realValue_0_266;
  wire       [7:0]    _zz__zz_realValue_0_266_1;
  wire       [7:0]    _zz_realValue_0_266_1;
  wire       [7:0]    _zz_realValue_0_266_2;
  wire       [7:0]    _zz_realValue_0_266_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_266;
  wire       [6:0]    _zz_when_ArraySlice_l166_266_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_266_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_266_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_266_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_266_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_266_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_266_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_267;
  wire       [7:0]    _zz_when_ArraySlice_l158_267_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_267_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_267_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_267;
  wire       [6:0]    _zz_when_ArraySlice_l159_267_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_267_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_267_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_267_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_267_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_267_6;
  wire       [7:0]    _zz__zz_realValue_0_267;
  wire       [7:0]    _zz__zz_realValue_0_267_1;
  wire       [7:0]    _zz_realValue_0_267_1;
  wire       [7:0]    _zz_realValue_0_267_2;
  wire       [7:0]    _zz_realValue_0_267_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_267;
  wire       [6:0]    _zz_when_ArraySlice_l166_267_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_267_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_267_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_267_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_267_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_267_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_267_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_268;
  wire       [7:0]    _zz_when_ArraySlice_l158_268_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_268_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_268_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_268;
  wire       [6:0]    _zz_when_ArraySlice_l159_268_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_268_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_268_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_268_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_268_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_268_6;
  wire       [7:0]    _zz__zz_realValue_0_268;
  wire       [7:0]    _zz__zz_realValue_0_268_1;
  wire       [7:0]    _zz_realValue_0_268_1;
  wire       [7:0]    _zz_realValue_0_268_2;
  wire       [7:0]    _zz_realValue_0_268_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_268;
  wire       [6:0]    _zz_when_ArraySlice_l166_268_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_268_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_268_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_268_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_268_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_268_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_268_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_269;
  wire       [7:0]    _zz_when_ArraySlice_l158_269_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_269_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_269_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_269;
  wire       [5:0]    _zz_when_ArraySlice_l159_269_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_269_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_269_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_269_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_269_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_269_6;
  wire       [7:0]    _zz__zz_realValue_0_269;
  wire       [7:0]    _zz__zz_realValue_0_269_1;
  wire       [7:0]    _zz_realValue_0_269_1;
  wire       [7:0]    _zz_realValue_0_269_2;
  wire       [7:0]    _zz_realValue_0_269_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_269;
  wire       [5:0]    _zz_when_ArraySlice_l166_269_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_269_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_269_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_269_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_269_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_269_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_269_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_270;
  wire       [7:0]    _zz_when_ArraySlice_l158_270_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_270_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_270_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_270;
  wire       [5:0]    _zz_when_ArraySlice_l159_270_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_270_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_270_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_270_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_270_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_270_6;
  wire       [7:0]    _zz__zz_realValue_0_270;
  wire       [7:0]    _zz__zz_realValue_0_270_1;
  wire       [7:0]    _zz_realValue_0_270_1;
  wire       [7:0]    _zz_realValue_0_270_2;
  wire       [7:0]    _zz_realValue_0_270_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_270;
  wire       [5:0]    _zz_when_ArraySlice_l166_270_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_270_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_270_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_270_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_270_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_270_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_270_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_271;
  wire       [7:0]    _zz_when_ArraySlice_l158_271_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_271_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_271_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_271;
  wire       [4:0]    _zz_when_ArraySlice_l159_271_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_271_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_271_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_271_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_271_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_271_6;
  wire       [7:0]    _zz__zz_realValue_0_271;
  wire       [7:0]    _zz__zz_realValue_0_271_1;
  wire       [7:0]    _zz_realValue_0_271_1;
  wire       [7:0]    _zz_realValue_0_271_2;
  wire       [7:0]    _zz_realValue_0_271_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_271;
  wire       [4:0]    _zz_when_ArraySlice_l166_271_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_271_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_271_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_271_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_271_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_271_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_271_7;
  wire                _zz_when_ArraySlice_l282_2_1;
  wire                _zz_when_ArraySlice_l282_2_2;
  wire                _zz_when_ArraySlice_l282_2_3;
  wire                _zz_when_ArraySlice_l282_2_4;
  wire                _zz_when_ArraySlice_l282_2_5;
  wire                _zz_when_ArraySlice_l282_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_2_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_2_7;
  wire       [5:0]    _zz_when_ArraySlice_l285_2_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l288_2_4;
  wire       [6:0]    _zz_when_ArraySlice_l288_2_5;
  wire       [7:0]    _zz_selectReadFifo_2_27;
  wire       [7:0]    _zz_selectReadFifo_2_28;
  wire       [6:0]    _zz_selectReadFifo_2_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_2;
  wire       [12:0]   _zz_when_ArraySlice_l295_2_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l306_2_3;
  wire       [7:0]    _zz__zz_realValue1_0_32;
  wire       [7:0]    _zz__zz_realValue1_0_32_1;
  wire       [7:0]    _zz_realValue1_0_32_1;
  wire       [7:0]    _zz_realValue1_0_32_2;
  wire       [7:0]    _zz_realValue1_0_32_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_2_1;
  wire       [6:0]    _zz_when_ArraySlice_l307_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l307_2_3;
  wire       [7:0]    _zz_selectReadFifo_2_30;
  wire       [7:0]    _zz_selectReadFifo_2_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_272;
  wire       [7:0]    _zz_when_ArraySlice_l158_272_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_272_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_272_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_272;
  wire       [7:0]    _zz_when_ArraySlice_l159_272_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_272_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_272_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_272_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_272_5;
  wire       [7:0]    _zz__zz_realValue_0_272;
  wire       [7:0]    _zz__zz_realValue_0_272_1;
  wire       [7:0]    _zz_realValue_0_272_1;
  wire       [7:0]    _zz_realValue_0_272_2;
  wire       [7:0]    _zz_realValue_0_272_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_272;
  wire       [7:0]    _zz_when_ArraySlice_l166_272_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_272_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_272_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_272_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_272_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_272_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_273;
  wire       [7:0]    _zz_when_ArraySlice_l158_273_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_273_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_273_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_273;
  wire       [6:0]    _zz_when_ArraySlice_l159_273_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_273_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_273_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_273_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_273_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_273_6;
  wire       [7:0]    _zz__zz_realValue_0_273;
  wire       [7:0]    _zz__zz_realValue_0_273_1;
  wire       [7:0]    _zz_realValue_0_273_1;
  wire       [7:0]    _zz_realValue_0_273_2;
  wire       [7:0]    _zz_realValue_0_273_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_273;
  wire       [6:0]    _zz_when_ArraySlice_l166_273_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_273_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_273_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_273_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_273_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_273_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_273_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_274;
  wire       [7:0]    _zz_when_ArraySlice_l158_274_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_274_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_274_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_274;
  wire       [6:0]    _zz_when_ArraySlice_l159_274_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_274_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_274_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_274_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_274_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_274_6;
  wire       [7:0]    _zz__zz_realValue_0_274;
  wire       [7:0]    _zz__zz_realValue_0_274_1;
  wire       [7:0]    _zz_realValue_0_274_1;
  wire       [7:0]    _zz_realValue_0_274_2;
  wire       [7:0]    _zz_realValue_0_274_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_274;
  wire       [6:0]    _zz_when_ArraySlice_l166_274_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_274_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_274_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_274_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_274_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_274_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_274_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_275;
  wire       [7:0]    _zz_when_ArraySlice_l158_275_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_275_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_275_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_275;
  wire       [6:0]    _zz_when_ArraySlice_l159_275_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_275_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_275_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_275_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_275_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_275_6;
  wire       [7:0]    _zz__zz_realValue_0_275;
  wire       [7:0]    _zz__zz_realValue_0_275_1;
  wire       [7:0]    _zz_realValue_0_275_1;
  wire       [7:0]    _zz_realValue_0_275_2;
  wire       [7:0]    _zz_realValue_0_275_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_275;
  wire       [6:0]    _zz_when_ArraySlice_l166_275_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_275_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_275_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_275_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_275_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_275_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_275_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_276;
  wire       [7:0]    _zz_when_ArraySlice_l158_276_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_276_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_276_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_276;
  wire       [6:0]    _zz_when_ArraySlice_l159_276_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_276_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_276_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_276_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_276_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_276_6;
  wire       [7:0]    _zz__zz_realValue_0_276;
  wire       [7:0]    _zz__zz_realValue_0_276_1;
  wire       [7:0]    _zz_realValue_0_276_1;
  wire       [7:0]    _zz_realValue_0_276_2;
  wire       [7:0]    _zz_realValue_0_276_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_276;
  wire       [6:0]    _zz_when_ArraySlice_l166_276_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_276_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_276_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_276_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_276_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_276_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_276_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_277;
  wire       [7:0]    _zz_when_ArraySlice_l158_277_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_277_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_277_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_277;
  wire       [5:0]    _zz_when_ArraySlice_l159_277_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_277_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_277_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_277_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_277_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_277_6;
  wire       [7:0]    _zz__zz_realValue_0_277;
  wire       [7:0]    _zz__zz_realValue_0_277_1;
  wire       [7:0]    _zz_realValue_0_277_1;
  wire       [7:0]    _zz_realValue_0_277_2;
  wire       [7:0]    _zz_realValue_0_277_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_277;
  wire       [5:0]    _zz_when_ArraySlice_l166_277_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_277_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_277_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_277_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_277_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_277_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_277_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_278;
  wire       [7:0]    _zz_when_ArraySlice_l158_278_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_278_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_278_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_278;
  wire       [5:0]    _zz_when_ArraySlice_l159_278_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_278_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_278_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_278_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_278_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_278_6;
  wire       [7:0]    _zz__zz_realValue_0_278;
  wire       [7:0]    _zz__zz_realValue_0_278_1;
  wire       [7:0]    _zz_realValue_0_278_1;
  wire       [7:0]    _zz_realValue_0_278_2;
  wire       [7:0]    _zz_realValue_0_278_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_278;
  wire       [5:0]    _zz_when_ArraySlice_l166_278_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_278_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_278_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_278_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_278_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_278_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_278_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_279;
  wire       [7:0]    _zz_when_ArraySlice_l158_279_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_279_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_279_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_279;
  wire       [4:0]    _zz_when_ArraySlice_l159_279_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_279_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_279_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_279_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_279_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_279_6;
  wire       [7:0]    _zz__zz_realValue_0_279;
  wire       [7:0]    _zz__zz_realValue_0_279_1;
  wire       [7:0]    _zz_realValue_0_279_1;
  wire       [7:0]    _zz_realValue_0_279_2;
  wire       [7:0]    _zz_realValue_0_279_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_279;
  wire       [4:0]    _zz_when_ArraySlice_l166_279_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_279_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_279_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_279_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_279_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_279_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_279_7;
  wire                _zz_when_ArraySlice_l314_2_1;
  wire                _zz_when_ArraySlice_l314_2_2;
  wire                _zz_when_ArraySlice_l314_2_3;
  wire                _zz_when_ArraySlice_l314_2_4;
  wire                _zz_when_ArraySlice_l314_2_5;
  wire                _zz_when_ArraySlice_l314_2_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_2;
  wire       [12:0]   _zz_when_ArraySlice_l318_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l304_2_3;
  wire       [5:0]    _zz_when_ArraySlice_l304_2_4;
  wire       [12:0]   _zz_when_ArraySlice_l325_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l325_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l233_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l233_3_2;
  wire       [5:0]    _zz_when_ArraySlice_l233_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l233_3_4;
  reg        [6:0]    _zz_when_ArraySlice_l234_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l234_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l234_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l234_3_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_3_valid_1_1;
  wire       [5:0]    _zz__zz_outputStreamArrayData_3_valid_1_2;
  wire       [6:0]    _zz__zz_14;
  reg                 _zz_outputStreamArrayData_3_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_3_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_3_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_3_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l240_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l240_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l240_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l241_3;
  wire       [7:0]    _zz_when_ArraySlice_l241_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_16;
  wire       [7:0]    _zz_selectReadFifo_3_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_3;
  wire       [12:0]   _zz_when_ArraySlice_l244_3_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l249_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l249_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l249_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l250_3;
  wire       [7:0]    _zz_when_ArraySlice_l250_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_3_2;
  wire       [7:0]    _zz__zz_realValue1_0_33;
  wire       [7:0]    _zz__zz_realValue1_0_33_1;
  wire       [7:0]    _zz_realValue1_0_33_1;
  wire       [7:0]    _zz_realValue1_0_33_2;
  wire       [7:0]    _zz_realValue1_0_33_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_3;
  wire       [6:0]    _zz_when_ArraySlice_l252_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_18;
  wire       [7:0]    _zz_selectReadFifo_3_19;
  wire       [7:0]    _zz_selectReadFifo_3_20;
  wire       [0:0]    _zz_selectReadFifo_3_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_280;
  wire       [7:0]    _zz_when_ArraySlice_l158_280_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_280_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_280_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_280;
  wire       [7:0]    _zz_when_ArraySlice_l159_280_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_280_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_280_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_280_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_280_5;
  wire       [7:0]    _zz__zz_realValue_0_280;
  wire       [7:0]    _zz__zz_realValue_0_280_1;
  wire       [7:0]    _zz_realValue_0_280_1;
  wire       [7:0]    _zz_realValue_0_280_2;
  wire       [7:0]    _zz_realValue_0_280_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_280;
  wire       [7:0]    _zz_when_ArraySlice_l166_280_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_280_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_280_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_280_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_280_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_280_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_281;
  wire       [7:0]    _zz_when_ArraySlice_l158_281_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_281_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_281_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_281;
  wire       [6:0]    _zz_when_ArraySlice_l159_281_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_281_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_281_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_281_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_281_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_281_6;
  wire       [7:0]    _zz__zz_realValue_0_281;
  wire       [7:0]    _zz__zz_realValue_0_281_1;
  wire       [7:0]    _zz_realValue_0_281_1;
  wire       [7:0]    _zz_realValue_0_281_2;
  wire       [7:0]    _zz_realValue_0_281_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_281;
  wire       [6:0]    _zz_when_ArraySlice_l166_281_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_281_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_281_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_281_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_281_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_281_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_281_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_282;
  wire       [7:0]    _zz_when_ArraySlice_l158_282_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_282_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_282_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_282;
  wire       [6:0]    _zz_when_ArraySlice_l159_282_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_282_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_282_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_282_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_282_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_282_6;
  wire       [7:0]    _zz__zz_realValue_0_282;
  wire       [7:0]    _zz__zz_realValue_0_282_1;
  wire       [7:0]    _zz_realValue_0_282_1;
  wire       [7:0]    _zz_realValue_0_282_2;
  wire       [7:0]    _zz_realValue_0_282_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_282;
  wire       [6:0]    _zz_when_ArraySlice_l166_282_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_282_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_282_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_282_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_282_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_282_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_282_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_283;
  wire       [7:0]    _zz_when_ArraySlice_l158_283_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_283_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_283_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_283;
  wire       [6:0]    _zz_when_ArraySlice_l159_283_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_283_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_283_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_283_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_283_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_283_6;
  wire       [7:0]    _zz__zz_realValue_0_283;
  wire       [7:0]    _zz__zz_realValue_0_283_1;
  wire       [7:0]    _zz_realValue_0_283_1;
  wire       [7:0]    _zz_realValue_0_283_2;
  wire       [7:0]    _zz_realValue_0_283_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_283;
  wire       [6:0]    _zz_when_ArraySlice_l166_283_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_283_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_283_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_283_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_283_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_283_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_283_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_284;
  wire       [7:0]    _zz_when_ArraySlice_l158_284_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_284_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_284_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_284;
  wire       [6:0]    _zz_when_ArraySlice_l159_284_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_284_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_284_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_284_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_284_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_284_6;
  wire       [7:0]    _zz__zz_realValue_0_284;
  wire       [7:0]    _zz__zz_realValue_0_284_1;
  wire       [7:0]    _zz_realValue_0_284_1;
  wire       [7:0]    _zz_realValue_0_284_2;
  wire       [7:0]    _zz_realValue_0_284_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_284;
  wire       [6:0]    _zz_when_ArraySlice_l166_284_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_284_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_284_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_284_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_284_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_284_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_284_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_285;
  wire       [7:0]    _zz_when_ArraySlice_l158_285_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_285_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_285_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_285;
  wire       [5:0]    _zz_when_ArraySlice_l159_285_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_285_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_285_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_285_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_285_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_285_6;
  wire       [7:0]    _zz__zz_realValue_0_285;
  wire       [7:0]    _zz__zz_realValue_0_285_1;
  wire       [7:0]    _zz_realValue_0_285_1;
  wire       [7:0]    _zz_realValue_0_285_2;
  wire       [7:0]    _zz_realValue_0_285_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_285;
  wire       [5:0]    _zz_when_ArraySlice_l166_285_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_285_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_285_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_285_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_285_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_285_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_285_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_286;
  wire       [7:0]    _zz_when_ArraySlice_l158_286_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_286_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_286_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_286;
  wire       [5:0]    _zz_when_ArraySlice_l159_286_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_286_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_286_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_286_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_286_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_286_6;
  wire       [7:0]    _zz__zz_realValue_0_286;
  wire       [7:0]    _zz__zz_realValue_0_286_1;
  wire       [7:0]    _zz_realValue_0_286_1;
  wire       [7:0]    _zz_realValue_0_286_2;
  wire       [7:0]    _zz_realValue_0_286_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_286;
  wire       [5:0]    _zz_when_ArraySlice_l166_286_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_286_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_286_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_286_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_286_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_286_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_286_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_287;
  wire       [7:0]    _zz_when_ArraySlice_l158_287_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_287_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_287_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_287;
  wire       [4:0]    _zz_when_ArraySlice_l159_287_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_287_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_287_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_287_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_287_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_287_6;
  wire       [7:0]    _zz__zz_realValue_0_287;
  wire       [7:0]    _zz__zz_realValue_0_287_1;
  wire       [7:0]    _zz_realValue_0_287_1;
  wire       [7:0]    _zz_realValue_0_287_2;
  wire       [7:0]    _zz_realValue_0_287_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_287;
  wire       [4:0]    _zz_when_ArraySlice_l166_287_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_287_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_287_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_287_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_287_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_287_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_287_7;
  wire                _zz_when_ArraySlice_l257_3_1;
  wire                _zz_when_ArraySlice_l257_3_2;
  wire                _zz_when_ArraySlice_l257_3_3;
  wire                _zz_when_ArraySlice_l257_3_4;
  wire                _zz_when_ArraySlice_l257_3_5;
  wire                _zz_when_ArraySlice_l257_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_3_7;
  wire       [5:0]    _zz_when_ArraySlice_l260_3_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l263_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l263_3_5;
  wire       [7:0]    _zz_selectReadFifo_3_22;
  wire       [7:0]    _zz_selectReadFifo_3_23;
  wire       [6:0]    _zz_selectReadFifo_3_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_3;
  wire       [12:0]   _zz_when_ArraySlice_l270_3_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_3_1;
  wire       [6:0]    _zz_when_ArraySlice_l274_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l274_3_4;
  wire       [5:0]    _zz_when_ArraySlice_l274_3_5;
  wire       [12:0]   _zz_when_ArraySlice_l275_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l275_3_4;
  wire       [0:0]    _zz_when_ArraySlice_l275_3_5;
  wire       [7:0]    _zz__zz_realValue1_0_34;
  wire       [7:0]    _zz__zz_realValue1_0_34_1;
  wire       [7:0]    _zz_realValue1_0_34_1;
  wire       [7:0]    _zz_realValue1_0_34_2;
  wire       [7:0]    _zz_realValue1_0_34_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_3;
  wire       [6:0]    _zz_when_ArraySlice_l277_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_25;
  wire       [7:0]    _zz_selectReadFifo_3_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_288;
  wire       [7:0]    _zz_when_ArraySlice_l158_288_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_288_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_288_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_288;
  wire       [7:0]    _zz_when_ArraySlice_l159_288_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_288_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_288_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_288_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_288_5;
  wire       [7:0]    _zz__zz_realValue_0_288;
  wire       [7:0]    _zz__zz_realValue_0_288_1;
  wire       [7:0]    _zz_realValue_0_288_1;
  wire       [7:0]    _zz_realValue_0_288_2;
  wire       [7:0]    _zz_realValue_0_288_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_288;
  wire       [7:0]    _zz_when_ArraySlice_l166_288_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_288_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_288_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_288_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_288_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_288_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_289;
  wire       [7:0]    _zz_when_ArraySlice_l158_289_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_289_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_289_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_289;
  wire       [6:0]    _zz_when_ArraySlice_l159_289_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_289_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_289_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_289_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_289_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_289_6;
  wire       [7:0]    _zz__zz_realValue_0_289;
  wire       [7:0]    _zz__zz_realValue_0_289_1;
  wire       [7:0]    _zz_realValue_0_289_1;
  wire       [7:0]    _zz_realValue_0_289_2;
  wire       [7:0]    _zz_realValue_0_289_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_289;
  wire       [6:0]    _zz_when_ArraySlice_l166_289_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_289_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_289_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_289_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_289_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_289_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_289_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_290;
  wire       [7:0]    _zz_when_ArraySlice_l158_290_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_290_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_290_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_290;
  wire       [6:0]    _zz_when_ArraySlice_l159_290_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_290_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_290_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_290_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_290_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_290_6;
  wire       [7:0]    _zz__zz_realValue_0_290;
  wire       [7:0]    _zz__zz_realValue_0_290_1;
  wire       [7:0]    _zz_realValue_0_290_1;
  wire       [7:0]    _zz_realValue_0_290_2;
  wire       [7:0]    _zz_realValue_0_290_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_290;
  wire       [6:0]    _zz_when_ArraySlice_l166_290_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_290_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_290_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_290_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_290_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_290_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_290_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_291;
  wire       [7:0]    _zz_when_ArraySlice_l158_291_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_291_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_291_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_291;
  wire       [6:0]    _zz_when_ArraySlice_l159_291_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_291_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_291_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_291_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_291_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_291_6;
  wire       [7:0]    _zz__zz_realValue_0_291;
  wire       [7:0]    _zz__zz_realValue_0_291_1;
  wire       [7:0]    _zz_realValue_0_291_1;
  wire       [7:0]    _zz_realValue_0_291_2;
  wire       [7:0]    _zz_realValue_0_291_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_291;
  wire       [6:0]    _zz_when_ArraySlice_l166_291_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_291_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_291_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_291_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_291_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_291_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_291_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_292;
  wire       [7:0]    _zz_when_ArraySlice_l158_292_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_292_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_292_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_292;
  wire       [6:0]    _zz_when_ArraySlice_l159_292_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_292_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_292_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_292_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_292_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_292_6;
  wire       [7:0]    _zz__zz_realValue_0_292;
  wire       [7:0]    _zz__zz_realValue_0_292_1;
  wire       [7:0]    _zz_realValue_0_292_1;
  wire       [7:0]    _zz_realValue_0_292_2;
  wire       [7:0]    _zz_realValue_0_292_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_292;
  wire       [6:0]    _zz_when_ArraySlice_l166_292_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_292_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_292_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_292_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_292_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_292_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_292_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_293;
  wire       [7:0]    _zz_when_ArraySlice_l158_293_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_293_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_293_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_293;
  wire       [5:0]    _zz_when_ArraySlice_l159_293_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_293_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_293_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_293_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_293_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_293_6;
  wire       [7:0]    _zz__zz_realValue_0_293;
  wire       [7:0]    _zz__zz_realValue_0_293_1;
  wire       [7:0]    _zz_realValue_0_293_1;
  wire       [7:0]    _zz_realValue_0_293_2;
  wire       [7:0]    _zz_realValue_0_293_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_293;
  wire       [5:0]    _zz_when_ArraySlice_l166_293_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_293_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_293_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_293_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_293_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_293_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_293_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_294;
  wire       [7:0]    _zz_when_ArraySlice_l158_294_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_294_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_294_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_294;
  wire       [5:0]    _zz_when_ArraySlice_l159_294_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_294_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_294_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_294_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_294_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_294_6;
  wire       [7:0]    _zz__zz_realValue_0_294;
  wire       [7:0]    _zz__zz_realValue_0_294_1;
  wire       [7:0]    _zz_realValue_0_294_1;
  wire       [7:0]    _zz_realValue_0_294_2;
  wire       [7:0]    _zz_realValue_0_294_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_294;
  wire       [5:0]    _zz_when_ArraySlice_l166_294_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_294_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_294_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_294_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_294_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_294_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_294_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_295;
  wire       [7:0]    _zz_when_ArraySlice_l158_295_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_295_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_295_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_295;
  wire       [4:0]    _zz_when_ArraySlice_l159_295_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_295_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_295_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_295_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_295_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_295_6;
  wire       [7:0]    _zz__zz_realValue_0_295;
  wire       [7:0]    _zz__zz_realValue_0_295_1;
  wire       [7:0]    _zz_realValue_0_295_1;
  wire       [7:0]    _zz_realValue_0_295_2;
  wire       [7:0]    _zz_realValue_0_295_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_295;
  wire       [4:0]    _zz_when_ArraySlice_l166_295_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_295_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_295_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_295_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_295_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_295_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_295_7;
  wire                _zz_when_ArraySlice_l282_3_1;
  wire                _zz_when_ArraySlice_l282_3_2;
  wire                _zz_when_ArraySlice_l282_3_3;
  wire                _zz_when_ArraySlice_l282_3_4;
  wire                _zz_when_ArraySlice_l282_3_5;
  wire                _zz_when_ArraySlice_l282_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_3_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_3_7;
  wire       [5:0]    _zz_when_ArraySlice_l285_3_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_3_3;
  wire       [7:0]    _zz_when_ArraySlice_l288_3_4;
  wire       [6:0]    _zz_when_ArraySlice_l288_3_5;
  wire       [7:0]    _zz_selectReadFifo_3_27;
  wire       [7:0]    _zz_selectReadFifo_3_28;
  wire       [6:0]    _zz_selectReadFifo_3_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_3;
  wire       [12:0]   _zz_when_ArraySlice_l295_3_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_3;
  wire       [7:0]    _zz_when_ArraySlice_l306_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_3_2;
  wire       [7:0]    _zz__zz_realValue1_0_35;
  wire       [7:0]    _zz__zz_realValue1_0_35_1;
  wire       [7:0]    _zz_realValue1_0_35_1;
  wire       [7:0]    _zz_realValue1_0_35_2;
  wire       [7:0]    _zz_realValue1_0_35_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_3;
  wire       [6:0]    _zz_when_ArraySlice_l307_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_3_2;
  wire       [7:0]    _zz_selectReadFifo_3_30;
  wire       [7:0]    _zz_selectReadFifo_3_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_296;
  wire       [7:0]    _zz_when_ArraySlice_l158_296_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_296_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_296_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_296;
  wire       [7:0]    _zz_when_ArraySlice_l159_296_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_296_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_296_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_296_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_296_5;
  wire       [7:0]    _zz__zz_realValue_0_296;
  wire       [7:0]    _zz__zz_realValue_0_296_1;
  wire       [7:0]    _zz_realValue_0_296_1;
  wire       [7:0]    _zz_realValue_0_296_2;
  wire       [7:0]    _zz_realValue_0_296_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_296;
  wire       [7:0]    _zz_when_ArraySlice_l166_296_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_296_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_296_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_296_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_296_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_296_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_297;
  wire       [7:0]    _zz_when_ArraySlice_l158_297_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_297_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_297_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_297;
  wire       [6:0]    _zz_when_ArraySlice_l159_297_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_297_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_297_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_297_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_297_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_297_6;
  wire       [7:0]    _zz__zz_realValue_0_297;
  wire       [7:0]    _zz__zz_realValue_0_297_1;
  wire       [7:0]    _zz_realValue_0_297_1;
  wire       [7:0]    _zz_realValue_0_297_2;
  wire       [7:0]    _zz_realValue_0_297_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_297;
  wire       [6:0]    _zz_when_ArraySlice_l166_297_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_297_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_297_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_297_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_297_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_297_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_297_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_298;
  wire       [7:0]    _zz_when_ArraySlice_l158_298_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_298_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_298_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_298;
  wire       [6:0]    _zz_when_ArraySlice_l159_298_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_298_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_298_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_298_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_298_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_298_6;
  wire       [7:0]    _zz__zz_realValue_0_298;
  wire       [7:0]    _zz__zz_realValue_0_298_1;
  wire       [7:0]    _zz_realValue_0_298_1;
  wire       [7:0]    _zz_realValue_0_298_2;
  wire       [7:0]    _zz_realValue_0_298_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_298;
  wire       [6:0]    _zz_when_ArraySlice_l166_298_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_298_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_298_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_298_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_298_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_298_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_298_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_299;
  wire       [7:0]    _zz_when_ArraySlice_l158_299_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_299_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_299_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_299;
  wire       [6:0]    _zz_when_ArraySlice_l159_299_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_299_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_299_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_299_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_299_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_299_6;
  wire       [7:0]    _zz__zz_realValue_0_299;
  wire       [7:0]    _zz__zz_realValue_0_299_1;
  wire       [7:0]    _zz_realValue_0_299_1;
  wire       [7:0]    _zz_realValue_0_299_2;
  wire       [7:0]    _zz_realValue_0_299_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_299;
  wire       [6:0]    _zz_when_ArraySlice_l166_299_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_299_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_299_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_299_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_299_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_299_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_299_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_300;
  wire       [7:0]    _zz_when_ArraySlice_l158_300_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_300_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_300_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_300;
  wire       [6:0]    _zz_when_ArraySlice_l159_300_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_300_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_300_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_300_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_300_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_300_6;
  wire       [7:0]    _zz__zz_realValue_0_300;
  wire       [7:0]    _zz__zz_realValue_0_300_1;
  wire       [7:0]    _zz_realValue_0_300_1;
  wire       [7:0]    _zz_realValue_0_300_2;
  wire       [7:0]    _zz_realValue_0_300_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_300;
  wire       [6:0]    _zz_when_ArraySlice_l166_300_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_300_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_300_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_300_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_300_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_300_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_300_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_301;
  wire       [7:0]    _zz_when_ArraySlice_l158_301_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_301_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_301_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_301;
  wire       [5:0]    _zz_when_ArraySlice_l159_301_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_301_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_301_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_301_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_301_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_301_6;
  wire       [7:0]    _zz__zz_realValue_0_301;
  wire       [7:0]    _zz__zz_realValue_0_301_1;
  wire       [7:0]    _zz_realValue_0_301_1;
  wire       [7:0]    _zz_realValue_0_301_2;
  wire       [7:0]    _zz_realValue_0_301_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_301;
  wire       [5:0]    _zz_when_ArraySlice_l166_301_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_301_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_301_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_301_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_301_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_301_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_301_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_302;
  wire       [7:0]    _zz_when_ArraySlice_l158_302_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_302_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_302_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_302;
  wire       [5:0]    _zz_when_ArraySlice_l159_302_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_302_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_302_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_302_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_302_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_302_6;
  wire       [7:0]    _zz__zz_realValue_0_302;
  wire       [7:0]    _zz__zz_realValue_0_302_1;
  wire       [7:0]    _zz_realValue_0_302_1;
  wire       [7:0]    _zz_realValue_0_302_2;
  wire       [7:0]    _zz_realValue_0_302_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_302;
  wire       [5:0]    _zz_when_ArraySlice_l166_302_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_302_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_302_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_302_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_302_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_302_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_302_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_303;
  wire       [7:0]    _zz_when_ArraySlice_l158_303_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_303_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_303_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_303;
  wire       [4:0]    _zz_when_ArraySlice_l159_303_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_303_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_303_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_303_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_303_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_303_6;
  wire       [7:0]    _zz__zz_realValue_0_303;
  wire       [7:0]    _zz__zz_realValue_0_303_1;
  wire       [7:0]    _zz_realValue_0_303_1;
  wire       [7:0]    _zz_realValue_0_303_2;
  wire       [7:0]    _zz_realValue_0_303_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_303;
  wire       [4:0]    _zz_when_ArraySlice_l166_303_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_303_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_303_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_303_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_303_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_303_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_303_7;
  wire                _zz_when_ArraySlice_l314_3_1;
  wire                _zz_when_ArraySlice_l314_3_2;
  wire                _zz_when_ArraySlice_l314_3_3;
  wire                _zz_when_ArraySlice_l314_3_4;
  wire                _zz_when_ArraySlice_l314_3_5;
  wire                _zz_when_ArraySlice_l314_3_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_3;
  wire       [12:0]   _zz_when_ArraySlice_l318_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l304_3_3;
  wire       [5:0]    _zz_when_ArraySlice_l304_3_4;
  wire       [12:0]   _zz_when_ArraySlice_l325_3;
  wire       [7:0]    _zz_when_ArraySlice_l325_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_4;
  wire       [7:0]    _zz_when_ArraySlice_l233_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l233_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_4_3;
  reg        [6:0]    _zz_when_ArraySlice_l234_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l234_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l234_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l234_4_5;
  wire       [7:0]    _zz__zz_outputStreamArrayData_4_valid_1_1;
  wire       [6:0]    _zz__zz_outputStreamArrayData_4_valid_1_2;
  wire       [6:0]    _zz__zz_15;
  reg                 _zz_outputStreamArrayData_4_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_4_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_4_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_4_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l240_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l240_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l240_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l241_4;
  wire       [7:0]    _zz_when_ArraySlice_l241_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_16;
  wire       [7:0]    _zz_selectReadFifo_4_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_4;
  wire       [12:0]   _zz_when_ArraySlice_l244_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l249_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l249_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l249_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l250_4;
  wire       [7:0]    _zz_when_ArraySlice_l250_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_4_2;
  wire       [7:0]    _zz__zz_realValue1_0_36;
  wire       [7:0]    _zz__zz_realValue1_0_36_1;
  wire       [7:0]    _zz_realValue1_0_36_1;
  wire       [7:0]    _zz_realValue1_0_36_2;
  wire       [7:0]    _zz_realValue1_0_36_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_4;
  wire       [6:0]    _zz_when_ArraySlice_l252_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_18;
  wire       [7:0]    _zz_selectReadFifo_4_19;
  wire       [7:0]    _zz_selectReadFifo_4_20;
  wire       [0:0]    _zz_selectReadFifo_4_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_304;
  wire       [7:0]    _zz_when_ArraySlice_l158_304_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_304_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_304_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_304;
  wire       [7:0]    _zz_when_ArraySlice_l159_304_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_304_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_304_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_304_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_304_5;
  wire       [7:0]    _zz__zz_realValue_0_304;
  wire       [7:0]    _zz__zz_realValue_0_304_1;
  wire       [7:0]    _zz_realValue_0_304_1;
  wire       [7:0]    _zz_realValue_0_304_2;
  wire       [7:0]    _zz_realValue_0_304_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_304;
  wire       [7:0]    _zz_when_ArraySlice_l166_304_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_304_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_304_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_304_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_304_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_304_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_305;
  wire       [7:0]    _zz_when_ArraySlice_l158_305_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_305_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_305_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_305;
  wire       [6:0]    _zz_when_ArraySlice_l159_305_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_305_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_305_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_305_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_305_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_305_6;
  wire       [7:0]    _zz__zz_realValue_0_305;
  wire       [7:0]    _zz__zz_realValue_0_305_1;
  wire       [7:0]    _zz_realValue_0_305_1;
  wire       [7:0]    _zz_realValue_0_305_2;
  wire       [7:0]    _zz_realValue_0_305_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_305;
  wire       [6:0]    _zz_when_ArraySlice_l166_305_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_305_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_305_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_305_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_305_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_305_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_305_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_306;
  wire       [7:0]    _zz_when_ArraySlice_l158_306_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_306_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_306_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_306;
  wire       [6:0]    _zz_when_ArraySlice_l159_306_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_306_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_306_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_306_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_306_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_306_6;
  wire       [7:0]    _zz__zz_realValue_0_306;
  wire       [7:0]    _zz__zz_realValue_0_306_1;
  wire       [7:0]    _zz_realValue_0_306_1;
  wire       [7:0]    _zz_realValue_0_306_2;
  wire       [7:0]    _zz_realValue_0_306_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_306;
  wire       [6:0]    _zz_when_ArraySlice_l166_306_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_306_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_306_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_306_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_306_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_306_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_306_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_307;
  wire       [7:0]    _zz_when_ArraySlice_l158_307_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_307_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_307_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_307;
  wire       [6:0]    _zz_when_ArraySlice_l159_307_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_307_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_307_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_307_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_307_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_307_6;
  wire       [7:0]    _zz__zz_realValue_0_307;
  wire       [7:0]    _zz__zz_realValue_0_307_1;
  wire       [7:0]    _zz_realValue_0_307_1;
  wire       [7:0]    _zz_realValue_0_307_2;
  wire       [7:0]    _zz_realValue_0_307_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_307;
  wire       [6:0]    _zz_when_ArraySlice_l166_307_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_307_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_307_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_307_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_307_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_307_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_307_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_308;
  wire       [7:0]    _zz_when_ArraySlice_l158_308_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_308_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_308_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_308;
  wire       [6:0]    _zz_when_ArraySlice_l159_308_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_308_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_308_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_308_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_308_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_308_6;
  wire       [7:0]    _zz__zz_realValue_0_308;
  wire       [7:0]    _zz__zz_realValue_0_308_1;
  wire       [7:0]    _zz_realValue_0_308_1;
  wire       [7:0]    _zz_realValue_0_308_2;
  wire       [7:0]    _zz_realValue_0_308_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_308;
  wire       [6:0]    _zz_when_ArraySlice_l166_308_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_308_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_308_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_308_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_308_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_308_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_308_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_309;
  wire       [7:0]    _zz_when_ArraySlice_l158_309_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_309_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_309_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_309;
  wire       [5:0]    _zz_when_ArraySlice_l159_309_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_309_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_309_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_309_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_309_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_309_6;
  wire       [7:0]    _zz__zz_realValue_0_309;
  wire       [7:0]    _zz__zz_realValue_0_309_1;
  wire       [7:0]    _zz_realValue_0_309_1;
  wire       [7:0]    _zz_realValue_0_309_2;
  wire       [7:0]    _zz_realValue_0_309_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_309;
  wire       [5:0]    _zz_when_ArraySlice_l166_309_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_309_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_309_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_309_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_309_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_309_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_309_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_310;
  wire       [7:0]    _zz_when_ArraySlice_l158_310_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_310_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_310_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_310;
  wire       [5:0]    _zz_when_ArraySlice_l159_310_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_310_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_310_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_310_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_310_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_310_6;
  wire       [7:0]    _zz__zz_realValue_0_310;
  wire       [7:0]    _zz__zz_realValue_0_310_1;
  wire       [7:0]    _zz_realValue_0_310_1;
  wire       [7:0]    _zz_realValue_0_310_2;
  wire       [7:0]    _zz_realValue_0_310_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_310;
  wire       [5:0]    _zz_when_ArraySlice_l166_310_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_310_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_310_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_310_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_310_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_310_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_310_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_311;
  wire       [7:0]    _zz_when_ArraySlice_l158_311_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_311_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_311_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_311;
  wire       [4:0]    _zz_when_ArraySlice_l159_311_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_311_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_311_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_311_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_311_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_311_6;
  wire       [7:0]    _zz__zz_realValue_0_311;
  wire       [7:0]    _zz__zz_realValue_0_311_1;
  wire       [7:0]    _zz_realValue_0_311_1;
  wire       [7:0]    _zz_realValue_0_311_2;
  wire       [7:0]    _zz_realValue_0_311_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_311;
  wire       [4:0]    _zz_when_ArraySlice_l166_311_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_311_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_311_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_311_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_311_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_311_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_311_7;
  wire                _zz_when_ArraySlice_l257_4_1;
  wire                _zz_when_ArraySlice_l257_4_2;
  wire                _zz_when_ArraySlice_l257_4_3;
  wire                _zz_when_ArraySlice_l257_4_4;
  wire                _zz_when_ArraySlice_l257_4_5;
  wire                _zz_when_ArraySlice_l257_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_4_7;
  wire       [6:0]    _zz_when_ArraySlice_l260_4_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l263_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l263_4_5;
  wire       [7:0]    _zz_selectReadFifo_4_22;
  wire       [7:0]    _zz_selectReadFifo_4_23;
  wire       [6:0]    _zz_selectReadFifo_4_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_4;
  wire       [12:0]   _zz_when_ArraySlice_l270_4_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_4_1;
  wire       [6:0]    _zz_when_ArraySlice_l274_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l274_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l274_4_5;
  wire       [12:0]   _zz_when_ArraySlice_l275_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l275_4_4;
  wire       [0:0]    _zz_when_ArraySlice_l275_4_5;
  wire       [7:0]    _zz__zz_realValue1_0_37;
  wire       [7:0]    _zz__zz_realValue1_0_37_1;
  wire       [7:0]    _zz_realValue1_0_37_1;
  wire       [7:0]    _zz_realValue1_0_37_2;
  wire       [7:0]    _zz_realValue1_0_37_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_4;
  wire       [6:0]    _zz_when_ArraySlice_l277_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_25;
  wire       [7:0]    _zz_selectReadFifo_4_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_312;
  wire       [7:0]    _zz_when_ArraySlice_l158_312_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_312_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_312_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_312;
  wire       [7:0]    _zz_when_ArraySlice_l159_312_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_312_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_312_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_312_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_312_5;
  wire       [7:0]    _zz__zz_realValue_0_312;
  wire       [7:0]    _zz__zz_realValue_0_312_1;
  wire       [7:0]    _zz_realValue_0_312_1;
  wire       [7:0]    _zz_realValue_0_312_2;
  wire       [7:0]    _zz_realValue_0_312_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_312;
  wire       [7:0]    _zz_when_ArraySlice_l166_312_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_312_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_312_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_312_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_312_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_312_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_313;
  wire       [7:0]    _zz_when_ArraySlice_l158_313_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_313_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_313_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_313;
  wire       [6:0]    _zz_when_ArraySlice_l159_313_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_313_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_313_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_313_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_313_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_313_6;
  wire       [7:0]    _zz__zz_realValue_0_313;
  wire       [7:0]    _zz__zz_realValue_0_313_1;
  wire       [7:0]    _zz_realValue_0_313_1;
  wire       [7:0]    _zz_realValue_0_313_2;
  wire       [7:0]    _zz_realValue_0_313_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_313;
  wire       [6:0]    _zz_when_ArraySlice_l166_313_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_313_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_313_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_313_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_313_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_313_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_313_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_314;
  wire       [7:0]    _zz_when_ArraySlice_l158_314_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_314_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_314_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_314;
  wire       [6:0]    _zz_when_ArraySlice_l159_314_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_314_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_314_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_314_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_314_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_314_6;
  wire       [7:0]    _zz__zz_realValue_0_314;
  wire       [7:0]    _zz__zz_realValue_0_314_1;
  wire       [7:0]    _zz_realValue_0_314_1;
  wire       [7:0]    _zz_realValue_0_314_2;
  wire       [7:0]    _zz_realValue_0_314_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_314;
  wire       [6:0]    _zz_when_ArraySlice_l166_314_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_314_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_314_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_314_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_314_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_314_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_314_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_315;
  wire       [7:0]    _zz_when_ArraySlice_l158_315_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_315_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_315_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_315;
  wire       [6:0]    _zz_when_ArraySlice_l159_315_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_315_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_315_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_315_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_315_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_315_6;
  wire       [7:0]    _zz__zz_realValue_0_315;
  wire       [7:0]    _zz__zz_realValue_0_315_1;
  wire       [7:0]    _zz_realValue_0_315_1;
  wire       [7:0]    _zz_realValue_0_315_2;
  wire       [7:0]    _zz_realValue_0_315_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_315;
  wire       [6:0]    _zz_when_ArraySlice_l166_315_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_315_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_315_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_315_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_315_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_315_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_315_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_316;
  wire       [7:0]    _zz_when_ArraySlice_l158_316_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_316_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_316_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_316;
  wire       [6:0]    _zz_when_ArraySlice_l159_316_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_316_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_316_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_316_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_316_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_316_6;
  wire       [7:0]    _zz__zz_realValue_0_316;
  wire       [7:0]    _zz__zz_realValue_0_316_1;
  wire       [7:0]    _zz_realValue_0_316_1;
  wire       [7:0]    _zz_realValue_0_316_2;
  wire       [7:0]    _zz_realValue_0_316_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_316;
  wire       [6:0]    _zz_when_ArraySlice_l166_316_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_316_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_316_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_316_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_316_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_316_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_316_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_317;
  wire       [7:0]    _zz_when_ArraySlice_l158_317_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_317_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_317_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_317;
  wire       [5:0]    _zz_when_ArraySlice_l159_317_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_317_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_317_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_317_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_317_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_317_6;
  wire       [7:0]    _zz__zz_realValue_0_317;
  wire       [7:0]    _zz__zz_realValue_0_317_1;
  wire       [7:0]    _zz_realValue_0_317_1;
  wire       [7:0]    _zz_realValue_0_317_2;
  wire       [7:0]    _zz_realValue_0_317_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_317;
  wire       [5:0]    _zz_when_ArraySlice_l166_317_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_317_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_317_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_317_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_317_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_317_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_317_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_318;
  wire       [7:0]    _zz_when_ArraySlice_l158_318_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_318_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_318_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_318;
  wire       [5:0]    _zz_when_ArraySlice_l159_318_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_318_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_318_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_318_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_318_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_318_6;
  wire       [7:0]    _zz__zz_realValue_0_318;
  wire       [7:0]    _zz__zz_realValue_0_318_1;
  wire       [7:0]    _zz_realValue_0_318_1;
  wire       [7:0]    _zz_realValue_0_318_2;
  wire       [7:0]    _zz_realValue_0_318_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_318;
  wire       [5:0]    _zz_when_ArraySlice_l166_318_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_318_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_318_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_318_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_318_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_318_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_318_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_319;
  wire       [7:0]    _zz_when_ArraySlice_l158_319_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_319_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_319_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_319;
  wire       [4:0]    _zz_when_ArraySlice_l159_319_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_319_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_319_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_319_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_319_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_319_6;
  wire       [7:0]    _zz__zz_realValue_0_319;
  wire       [7:0]    _zz__zz_realValue_0_319_1;
  wire       [7:0]    _zz_realValue_0_319_1;
  wire       [7:0]    _zz_realValue_0_319_2;
  wire       [7:0]    _zz_realValue_0_319_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_319;
  wire       [4:0]    _zz_when_ArraySlice_l166_319_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_319_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_319_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_319_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_319_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_319_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_319_7;
  wire                _zz_when_ArraySlice_l282_4_1;
  wire                _zz_when_ArraySlice_l282_4_2;
  wire                _zz_when_ArraySlice_l282_4_3;
  wire                _zz_when_ArraySlice_l282_4_4;
  wire                _zz_when_ArraySlice_l282_4_5;
  wire                _zz_when_ArraySlice_l282_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_4_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_4_7;
  wire       [6:0]    _zz_when_ArraySlice_l285_4_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_4_3;
  wire       [7:0]    _zz_when_ArraySlice_l288_4_4;
  wire       [6:0]    _zz_when_ArraySlice_l288_4_5;
  wire       [7:0]    _zz_selectReadFifo_4_27;
  wire       [7:0]    _zz_selectReadFifo_4_28;
  wire       [6:0]    _zz_selectReadFifo_4_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_4;
  wire       [12:0]   _zz_when_ArraySlice_l295_4_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_4;
  wire       [7:0]    _zz_when_ArraySlice_l306_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_4_2;
  wire       [7:0]    _zz__zz_realValue1_0_38;
  wire       [7:0]    _zz__zz_realValue1_0_38_1;
  wire       [7:0]    _zz_realValue1_0_38_1;
  wire       [7:0]    _zz_realValue1_0_38_2;
  wire       [7:0]    _zz_realValue1_0_38_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_4;
  wire       [6:0]    _zz_when_ArraySlice_l307_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_4_2;
  wire       [7:0]    _zz_selectReadFifo_4_30;
  wire       [7:0]    _zz_selectReadFifo_4_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_320;
  wire       [7:0]    _zz_when_ArraySlice_l158_320_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_320_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_320_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_320;
  wire       [7:0]    _zz_when_ArraySlice_l159_320_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_320_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_320_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_320_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_320_5;
  wire       [7:0]    _zz__zz_realValue_0_320;
  wire       [7:0]    _zz__zz_realValue_0_320_1;
  wire       [7:0]    _zz_realValue_0_320_1;
  wire       [7:0]    _zz_realValue_0_320_2;
  wire       [7:0]    _zz_realValue_0_320_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_320;
  wire       [7:0]    _zz_when_ArraySlice_l166_320_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_320_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_320_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_320_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_320_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_320_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_321;
  wire       [7:0]    _zz_when_ArraySlice_l158_321_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_321_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_321_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_321;
  wire       [6:0]    _zz_when_ArraySlice_l159_321_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_321_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_321_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_321_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_321_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_321_6;
  wire       [7:0]    _zz__zz_realValue_0_321;
  wire       [7:0]    _zz__zz_realValue_0_321_1;
  wire       [7:0]    _zz_realValue_0_321_1;
  wire       [7:0]    _zz_realValue_0_321_2;
  wire       [7:0]    _zz_realValue_0_321_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_321;
  wire       [6:0]    _zz_when_ArraySlice_l166_321_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_321_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_321_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_321_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_321_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_321_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_321_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_322;
  wire       [7:0]    _zz_when_ArraySlice_l158_322_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_322_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_322_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_322;
  wire       [6:0]    _zz_when_ArraySlice_l159_322_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_322_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_322_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_322_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_322_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_322_6;
  wire       [7:0]    _zz__zz_realValue_0_322;
  wire       [7:0]    _zz__zz_realValue_0_322_1;
  wire       [7:0]    _zz_realValue_0_322_1;
  wire       [7:0]    _zz_realValue_0_322_2;
  wire       [7:0]    _zz_realValue_0_322_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_322;
  wire       [6:0]    _zz_when_ArraySlice_l166_322_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_322_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_322_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_322_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_322_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_322_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_322_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_323;
  wire       [7:0]    _zz_when_ArraySlice_l158_323_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_323_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_323_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_323;
  wire       [6:0]    _zz_when_ArraySlice_l159_323_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_323_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_323_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_323_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_323_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_323_6;
  wire       [7:0]    _zz__zz_realValue_0_323;
  wire       [7:0]    _zz__zz_realValue_0_323_1;
  wire       [7:0]    _zz_realValue_0_323_1;
  wire       [7:0]    _zz_realValue_0_323_2;
  wire       [7:0]    _zz_realValue_0_323_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_323;
  wire       [6:0]    _zz_when_ArraySlice_l166_323_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_323_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_323_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_323_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_323_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_323_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_323_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_324;
  wire       [7:0]    _zz_when_ArraySlice_l158_324_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_324_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_324_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_324;
  wire       [6:0]    _zz_when_ArraySlice_l159_324_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_324_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_324_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_324_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_324_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_324_6;
  wire       [7:0]    _zz__zz_realValue_0_324;
  wire       [7:0]    _zz__zz_realValue_0_324_1;
  wire       [7:0]    _zz_realValue_0_324_1;
  wire       [7:0]    _zz_realValue_0_324_2;
  wire       [7:0]    _zz_realValue_0_324_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_324;
  wire       [6:0]    _zz_when_ArraySlice_l166_324_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_324_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_324_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_324_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_324_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_324_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_324_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_325;
  wire       [7:0]    _zz_when_ArraySlice_l158_325_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_325_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_325_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_325;
  wire       [5:0]    _zz_when_ArraySlice_l159_325_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_325_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_325_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_325_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_325_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_325_6;
  wire       [7:0]    _zz__zz_realValue_0_325;
  wire       [7:0]    _zz__zz_realValue_0_325_1;
  wire       [7:0]    _zz_realValue_0_325_1;
  wire       [7:0]    _zz_realValue_0_325_2;
  wire       [7:0]    _zz_realValue_0_325_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_325;
  wire       [5:0]    _zz_when_ArraySlice_l166_325_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_325_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_325_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_325_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_325_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_325_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_325_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_326;
  wire       [7:0]    _zz_when_ArraySlice_l158_326_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_326_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_326_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_326;
  wire       [5:0]    _zz_when_ArraySlice_l159_326_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_326_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_326_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_326_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_326_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_326_6;
  wire       [7:0]    _zz__zz_realValue_0_326;
  wire       [7:0]    _zz__zz_realValue_0_326_1;
  wire       [7:0]    _zz_realValue_0_326_1;
  wire       [7:0]    _zz_realValue_0_326_2;
  wire       [7:0]    _zz_realValue_0_326_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_326;
  wire       [5:0]    _zz_when_ArraySlice_l166_326_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_326_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_326_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_326_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_326_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_326_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_326_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_327;
  wire       [7:0]    _zz_when_ArraySlice_l158_327_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_327_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_327_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_327;
  wire       [4:0]    _zz_when_ArraySlice_l159_327_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_327_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_327_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_327_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_327_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_327_6;
  wire       [7:0]    _zz__zz_realValue_0_327;
  wire       [7:0]    _zz__zz_realValue_0_327_1;
  wire       [7:0]    _zz_realValue_0_327_1;
  wire       [7:0]    _zz_realValue_0_327_2;
  wire       [7:0]    _zz_realValue_0_327_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_327;
  wire       [4:0]    _zz_when_ArraySlice_l166_327_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_327_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_327_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_327_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_327_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_327_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_327_7;
  wire                _zz_when_ArraySlice_l314_4_1;
  wire                _zz_when_ArraySlice_l314_4_2;
  wire                _zz_when_ArraySlice_l314_4_3;
  wire                _zz_when_ArraySlice_l314_4_4;
  wire                _zz_when_ArraySlice_l314_4_5;
  wire                _zz_when_ArraySlice_l314_4_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_4;
  wire       [12:0]   _zz_when_ArraySlice_l318_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_4;
  wire       [7:0]    _zz_when_ArraySlice_l304_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_4_2;
  wire       [6:0]    _zz_when_ArraySlice_l304_4_3;
  wire       [12:0]   _zz_when_ArraySlice_l325_4;
  wire       [7:0]    _zz_when_ArraySlice_l325_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_5;
  wire       [7:0]    _zz_when_ArraySlice_l233_5_1;
  wire       [6:0]    _zz_when_ArraySlice_l233_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_5_3;
  reg        [6:0]    _zz_when_ArraySlice_l234_5;
  wire       [6:0]    _zz_when_ArraySlice_l234_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l234_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l234_5_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_5_valid_1_1;
  wire       [6:0]    _zz__zz_outputStreamArrayData_5_valid_1_2;
  wire       [6:0]    _zz__zz_16;
  reg                 _zz_outputStreamArrayData_5_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_5_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_5_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_5_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_5;
  wire       [6:0]    _zz_when_ArraySlice_l240_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l240_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l240_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l241_5;
  wire       [7:0]    _zz_when_ArraySlice_l241_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_16;
  wire       [7:0]    _zz_selectReadFifo_5_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_5;
  wire       [12:0]   _zz_when_ArraySlice_l244_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_5;
  wire       [6:0]    _zz_when_ArraySlice_l249_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l249_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l249_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l250_5;
  wire       [7:0]    _zz_when_ArraySlice_l250_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_5_2;
  wire       [7:0]    _zz__zz_realValue1_0_39;
  wire       [7:0]    _zz__zz_realValue1_0_39_1;
  wire       [7:0]    _zz_realValue1_0_39_1;
  wire       [7:0]    _zz_realValue1_0_39_2;
  wire       [7:0]    _zz_realValue1_0_39_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_5;
  wire       [6:0]    _zz_when_ArraySlice_l252_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_18;
  wire       [7:0]    _zz_selectReadFifo_5_19;
  wire       [7:0]    _zz_selectReadFifo_5_20;
  wire       [0:0]    _zz_selectReadFifo_5_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_328;
  wire       [7:0]    _zz_when_ArraySlice_l158_328_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_328_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_328_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_328;
  wire       [7:0]    _zz_when_ArraySlice_l159_328_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_328_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_328_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_328_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_328_5;
  wire       [7:0]    _zz__zz_realValue_0_328;
  wire       [7:0]    _zz__zz_realValue_0_328_1;
  wire       [7:0]    _zz_realValue_0_328_1;
  wire       [7:0]    _zz_realValue_0_328_2;
  wire       [7:0]    _zz_realValue_0_328_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_328;
  wire       [7:0]    _zz_when_ArraySlice_l166_328_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_328_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_328_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_328_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_328_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_328_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_329;
  wire       [7:0]    _zz_when_ArraySlice_l158_329_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_329_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_329_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_329;
  wire       [6:0]    _zz_when_ArraySlice_l159_329_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_329_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_329_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_329_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_329_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_329_6;
  wire       [7:0]    _zz__zz_realValue_0_329;
  wire       [7:0]    _zz__zz_realValue_0_329_1;
  wire       [7:0]    _zz_realValue_0_329_1;
  wire       [7:0]    _zz_realValue_0_329_2;
  wire       [7:0]    _zz_realValue_0_329_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_329;
  wire       [6:0]    _zz_when_ArraySlice_l166_329_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_329_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_329_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_329_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_329_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_329_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_329_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_330;
  wire       [7:0]    _zz_when_ArraySlice_l158_330_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_330_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_330_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_330;
  wire       [6:0]    _zz_when_ArraySlice_l159_330_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_330_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_330_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_330_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_330_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_330_6;
  wire       [7:0]    _zz__zz_realValue_0_330;
  wire       [7:0]    _zz__zz_realValue_0_330_1;
  wire       [7:0]    _zz_realValue_0_330_1;
  wire       [7:0]    _zz_realValue_0_330_2;
  wire       [7:0]    _zz_realValue_0_330_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_330;
  wire       [6:0]    _zz_when_ArraySlice_l166_330_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_330_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_330_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_330_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_330_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_330_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_330_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_331;
  wire       [7:0]    _zz_when_ArraySlice_l158_331_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_331_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_331_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_331;
  wire       [6:0]    _zz_when_ArraySlice_l159_331_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_331_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_331_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_331_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_331_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_331_6;
  wire       [7:0]    _zz__zz_realValue_0_331;
  wire       [7:0]    _zz__zz_realValue_0_331_1;
  wire       [7:0]    _zz_realValue_0_331_1;
  wire       [7:0]    _zz_realValue_0_331_2;
  wire       [7:0]    _zz_realValue_0_331_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_331;
  wire       [6:0]    _zz_when_ArraySlice_l166_331_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_331_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_331_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_331_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_331_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_331_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_331_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_332;
  wire       [7:0]    _zz_when_ArraySlice_l158_332_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_332_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_332_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_332;
  wire       [6:0]    _zz_when_ArraySlice_l159_332_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_332_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_332_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_332_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_332_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_332_6;
  wire       [7:0]    _zz__zz_realValue_0_332;
  wire       [7:0]    _zz__zz_realValue_0_332_1;
  wire       [7:0]    _zz_realValue_0_332_1;
  wire       [7:0]    _zz_realValue_0_332_2;
  wire       [7:0]    _zz_realValue_0_332_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_332;
  wire       [6:0]    _zz_when_ArraySlice_l166_332_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_332_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_332_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_332_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_332_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_332_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_332_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_333;
  wire       [7:0]    _zz_when_ArraySlice_l158_333_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_333_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_333_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_333;
  wire       [5:0]    _zz_when_ArraySlice_l159_333_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_333_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_333_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_333_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_333_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_333_6;
  wire       [7:0]    _zz__zz_realValue_0_333;
  wire       [7:0]    _zz__zz_realValue_0_333_1;
  wire       [7:0]    _zz_realValue_0_333_1;
  wire       [7:0]    _zz_realValue_0_333_2;
  wire       [7:0]    _zz_realValue_0_333_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_333;
  wire       [5:0]    _zz_when_ArraySlice_l166_333_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_333_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_333_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_333_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_333_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_333_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_333_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_334;
  wire       [7:0]    _zz_when_ArraySlice_l158_334_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_334_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_334_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_334;
  wire       [5:0]    _zz_when_ArraySlice_l159_334_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_334_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_334_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_334_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_334_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_334_6;
  wire       [7:0]    _zz__zz_realValue_0_334;
  wire       [7:0]    _zz__zz_realValue_0_334_1;
  wire       [7:0]    _zz_realValue_0_334_1;
  wire       [7:0]    _zz_realValue_0_334_2;
  wire       [7:0]    _zz_realValue_0_334_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_334;
  wire       [5:0]    _zz_when_ArraySlice_l166_334_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_334_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_334_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_334_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_334_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_334_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_334_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_335;
  wire       [7:0]    _zz_when_ArraySlice_l158_335_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_335_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_335_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_335;
  wire       [4:0]    _zz_when_ArraySlice_l159_335_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_335_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_335_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_335_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_335_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_335_6;
  wire       [7:0]    _zz__zz_realValue_0_335;
  wire       [7:0]    _zz__zz_realValue_0_335_1;
  wire       [7:0]    _zz_realValue_0_335_1;
  wire       [7:0]    _zz_realValue_0_335_2;
  wire       [7:0]    _zz_realValue_0_335_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_335;
  wire       [4:0]    _zz_when_ArraySlice_l166_335_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_335_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_335_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_335_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_335_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_335_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_335_7;
  wire                _zz_when_ArraySlice_l257_5_1;
  wire                _zz_when_ArraySlice_l257_5_2;
  wire                _zz_when_ArraySlice_l257_5_3;
  wire                _zz_when_ArraySlice_l257_5_4;
  wire                _zz_when_ArraySlice_l257_5_5;
  wire                _zz_when_ArraySlice_l257_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_5_7;
  wire       [6:0]    _zz_when_ArraySlice_l260_5_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_5;
  wire       [7:0]    _zz_when_ArraySlice_l263_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l263_5_4;
  wire       [7:0]    _zz_selectReadFifo_5_22;
  wire       [7:0]    _zz_selectReadFifo_5_23;
  wire       [6:0]    _zz_selectReadFifo_5_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_5;
  wire       [12:0]   _zz_when_ArraySlice_l270_5_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_5;
  wire       [6:0]    _zz_when_ArraySlice_l274_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l274_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l274_5_4;
  wire       [12:0]   _zz_when_ArraySlice_l275_5;
  wire       [7:0]    _zz_when_ArraySlice_l275_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_5_3;
  wire       [0:0]    _zz_when_ArraySlice_l275_5_4;
  wire       [7:0]    _zz__zz_realValue1_0_40;
  wire       [7:0]    _zz__zz_realValue1_0_40_1;
  wire       [7:0]    _zz_realValue1_0_40_1;
  wire       [7:0]    _zz_realValue1_0_40_2;
  wire       [7:0]    _zz_realValue1_0_40_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_5;
  wire       [6:0]    _zz_when_ArraySlice_l277_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_25;
  wire       [7:0]    _zz_selectReadFifo_5_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_336;
  wire       [7:0]    _zz_when_ArraySlice_l158_336_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_336_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_336_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_336;
  wire       [7:0]    _zz_when_ArraySlice_l159_336_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_336_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_336_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_336_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_336_5;
  wire       [7:0]    _zz__zz_realValue_0_336;
  wire       [7:0]    _zz__zz_realValue_0_336_1;
  wire       [7:0]    _zz_realValue_0_336_1;
  wire       [7:0]    _zz_realValue_0_336_2;
  wire       [7:0]    _zz_realValue_0_336_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_336;
  wire       [7:0]    _zz_when_ArraySlice_l166_336_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_336_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_336_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_336_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_336_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_336_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_337;
  wire       [7:0]    _zz_when_ArraySlice_l158_337_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_337_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_337_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_337;
  wire       [6:0]    _zz_when_ArraySlice_l159_337_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_337_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_337_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_337_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_337_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_337_6;
  wire       [7:0]    _zz__zz_realValue_0_337;
  wire       [7:0]    _zz__zz_realValue_0_337_1;
  wire       [7:0]    _zz_realValue_0_337_1;
  wire       [7:0]    _zz_realValue_0_337_2;
  wire       [7:0]    _zz_realValue_0_337_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_337;
  wire       [6:0]    _zz_when_ArraySlice_l166_337_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_337_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_337_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_337_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_337_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_337_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_337_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_338;
  wire       [7:0]    _zz_when_ArraySlice_l158_338_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_338_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_338_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_338;
  wire       [6:0]    _zz_when_ArraySlice_l159_338_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_338_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_338_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_338_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_338_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_338_6;
  wire       [7:0]    _zz__zz_realValue_0_338;
  wire       [7:0]    _zz__zz_realValue_0_338_1;
  wire       [7:0]    _zz_realValue_0_338_1;
  wire       [7:0]    _zz_realValue_0_338_2;
  wire       [7:0]    _zz_realValue_0_338_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_338;
  wire       [6:0]    _zz_when_ArraySlice_l166_338_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_338_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_338_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_338_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_338_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_338_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_338_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_339;
  wire       [7:0]    _zz_when_ArraySlice_l158_339_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_339_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_339_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_339;
  wire       [6:0]    _zz_when_ArraySlice_l159_339_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_339_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_339_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_339_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_339_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_339_6;
  wire       [7:0]    _zz__zz_realValue_0_339;
  wire       [7:0]    _zz__zz_realValue_0_339_1;
  wire       [7:0]    _zz_realValue_0_339_1;
  wire       [7:0]    _zz_realValue_0_339_2;
  wire       [7:0]    _zz_realValue_0_339_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_339;
  wire       [6:0]    _zz_when_ArraySlice_l166_339_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_339_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_339_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_339_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_339_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_339_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_339_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_340;
  wire       [7:0]    _zz_when_ArraySlice_l158_340_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_340_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_340_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_340;
  wire       [6:0]    _zz_when_ArraySlice_l159_340_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_340_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_340_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_340_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_340_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_340_6;
  wire       [7:0]    _zz__zz_realValue_0_340;
  wire       [7:0]    _zz__zz_realValue_0_340_1;
  wire       [7:0]    _zz_realValue_0_340_1;
  wire       [7:0]    _zz_realValue_0_340_2;
  wire       [7:0]    _zz_realValue_0_340_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_340;
  wire       [6:0]    _zz_when_ArraySlice_l166_340_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_340_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_340_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_340_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_340_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_340_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_340_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_341;
  wire       [7:0]    _zz_when_ArraySlice_l158_341_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_341_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_341_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_341;
  wire       [5:0]    _zz_when_ArraySlice_l159_341_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_341_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_341_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_341_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_341_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_341_6;
  wire       [7:0]    _zz__zz_realValue_0_341;
  wire       [7:0]    _zz__zz_realValue_0_341_1;
  wire       [7:0]    _zz_realValue_0_341_1;
  wire       [7:0]    _zz_realValue_0_341_2;
  wire       [7:0]    _zz_realValue_0_341_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_341;
  wire       [5:0]    _zz_when_ArraySlice_l166_341_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_341_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_341_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_341_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_341_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_341_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_341_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_342;
  wire       [7:0]    _zz_when_ArraySlice_l158_342_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_342_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_342_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_342;
  wire       [5:0]    _zz_when_ArraySlice_l159_342_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_342_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_342_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_342_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_342_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_342_6;
  wire       [7:0]    _zz__zz_realValue_0_342;
  wire       [7:0]    _zz__zz_realValue_0_342_1;
  wire       [7:0]    _zz_realValue_0_342_1;
  wire       [7:0]    _zz_realValue_0_342_2;
  wire       [7:0]    _zz_realValue_0_342_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_342;
  wire       [5:0]    _zz_when_ArraySlice_l166_342_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_342_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_342_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_342_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_342_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_342_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_342_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_343;
  wire       [7:0]    _zz_when_ArraySlice_l158_343_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_343_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_343_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_343;
  wire       [4:0]    _zz_when_ArraySlice_l159_343_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_343_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_343_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_343_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_343_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_343_6;
  wire       [7:0]    _zz__zz_realValue_0_343;
  wire       [7:0]    _zz__zz_realValue_0_343_1;
  wire       [7:0]    _zz_realValue_0_343_1;
  wire       [7:0]    _zz_realValue_0_343_2;
  wire       [7:0]    _zz_realValue_0_343_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_343;
  wire       [4:0]    _zz_when_ArraySlice_l166_343_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_343_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_343_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_343_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_343_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_343_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_343_7;
  wire                _zz_when_ArraySlice_l282_5_1;
  wire                _zz_when_ArraySlice_l282_5_2;
  wire                _zz_when_ArraySlice_l282_5_3;
  wire                _zz_when_ArraySlice_l282_5_4;
  wire                _zz_when_ArraySlice_l282_5_5;
  wire                _zz_when_ArraySlice_l282_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_5_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_5_7;
  wire       [6:0]    _zz_when_ArraySlice_l285_5_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_5;
  wire       [7:0]    _zz_when_ArraySlice_l288_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_5_3;
  wire       [6:0]    _zz_when_ArraySlice_l288_5_4;
  wire       [7:0]    _zz_selectReadFifo_5_27;
  wire       [7:0]    _zz_selectReadFifo_5_28;
  wire       [6:0]    _zz_selectReadFifo_5_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_5;
  wire       [12:0]   _zz_when_ArraySlice_l295_5_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_5;
  wire       [7:0]    _zz_when_ArraySlice_l306_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_5_2;
  wire       [7:0]    _zz__zz_realValue1_0_41;
  wire       [7:0]    _zz__zz_realValue1_0_41_1;
  wire       [7:0]    _zz_realValue1_0_41_1;
  wire       [7:0]    _zz_realValue1_0_41_2;
  wire       [7:0]    _zz_realValue1_0_41_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_5;
  wire       [6:0]    _zz_when_ArraySlice_l307_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_5_2;
  wire       [7:0]    _zz_selectReadFifo_5_30;
  wire       [7:0]    _zz_selectReadFifo_5_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_344;
  wire       [7:0]    _zz_when_ArraySlice_l158_344_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_344_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_344_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_344;
  wire       [7:0]    _zz_when_ArraySlice_l159_344_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_344_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_344_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_344_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_344_5;
  wire       [7:0]    _zz__zz_realValue_0_344;
  wire       [7:0]    _zz__zz_realValue_0_344_1;
  wire       [7:0]    _zz_realValue_0_344_1;
  wire       [7:0]    _zz_realValue_0_344_2;
  wire       [7:0]    _zz_realValue_0_344_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_344;
  wire       [7:0]    _zz_when_ArraySlice_l166_344_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_344_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_344_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_344_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_344_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_344_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_345;
  wire       [7:0]    _zz_when_ArraySlice_l158_345_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_345_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_345_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_345;
  wire       [6:0]    _zz_when_ArraySlice_l159_345_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_345_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_345_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_345_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_345_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_345_6;
  wire       [7:0]    _zz__zz_realValue_0_345;
  wire       [7:0]    _zz__zz_realValue_0_345_1;
  wire       [7:0]    _zz_realValue_0_345_1;
  wire       [7:0]    _zz_realValue_0_345_2;
  wire       [7:0]    _zz_realValue_0_345_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_345;
  wire       [6:0]    _zz_when_ArraySlice_l166_345_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_345_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_345_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_345_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_345_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_345_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_345_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_346;
  wire       [7:0]    _zz_when_ArraySlice_l158_346_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_346_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_346_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_346;
  wire       [6:0]    _zz_when_ArraySlice_l159_346_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_346_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_346_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_346_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_346_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_346_6;
  wire       [7:0]    _zz__zz_realValue_0_346;
  wire       [7:0]    _zz__zz_realValue_0_346_1;
  wire       [7:0]    _zz_realValue_0_346_1;
  wire       [7:0]    _zz_realValue_0_346_2;
  wire       [7:0]    _zz_realValue_0_346_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_346;
  wire       [6:0]    _zz_when_ArraySlice_l166_346_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_346_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_346_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_346_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_346_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_346_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_346_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_347;
  wire       [7:0]    _zz_when_ArraySlice_l158_347_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_347_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_347_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_347;
  wire       [6:0]    _zz_when_ArraySlice_l159_347_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_347_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_347_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_347_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_347_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_347_6;
  wire       [7:0]    _zz__zz_realValue_0_347;
  wire       [7:0]    _zz__zz_realValue_0_347_1;
  wire       [7:0]    _zz_realValue_0_347_1;
  wire       [7:0]    _zz_realValue_0_347_2;
  wire       [7:0]    _zz_realValue_0_347_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_347;
  wire       [6:0]    _zz_when_ArraySlice_l166_347_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_347_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_347_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_347_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_347_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_347_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_347_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_348;
  wire       [7:0]    _zz_when_ArraySlice_l158_348_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_348_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_348_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_348;
  wire       [6:0]    _zz_when_ArraySlice_l159_348_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_348_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_348_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_348_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_348_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_348_6;
  wire       [7:0]    _zz__zz_realValue_0_348;
  wire       [7:0]    _zz__zz_realValue_0_348_1;
  wire       [7:0]    _zz_realValue_0_348_1;
  wire       [7:0]    _zz_realValue_0_348_2;
  wire       [7:0]    _zz_realValue_0_348_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_348;
  wire       [6:0]    _zz_when_ArraySlice_l166_348_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_348_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_348_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_348_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_348_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_348_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_348_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_349;
  wire       [7:0]    _zz_when_ArraySlice_l158_349_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_349_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_349_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_349;
  wire       [5:0]    _zz_when_ArraySlice_l159_349_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_349_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_349_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_349_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_349_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_349_6;
  wire       [7:0]    _zz__zz_realValue_0_349;
  wire       [7:0]    _zz__zz_realValue_0_349_1;
  wire       [7:0]    _zz_realValue_0_349_1;
  wire       [7:0]    _zz_realValue_0_349_2;
  wire       [7:0]    _zz_realValue_0_349_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_349;
  wire       [5:0]    _zz_when_ArraySlice_l166_349_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_349_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_349_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_349_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_349_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_349_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_349_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_350;
  wire       [7:0]    _zz_when_ArraySlice_l158_350_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_350_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_350_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_350;
  wire       [5:0]    _zz_when_ArraySlice_l159_350_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_350_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_350_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_350_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_350_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_350_6;
  wire       [7:0]    _zz__zz_realValue_0_350;
  wire       [7:0]    _zz__zz_realValue_0_350_1;
  wire       [7:0]    _zz_realValue_0_350_1;
  wire       [7:0]    _zz_realValue_0_350_2;
  wire       [7:0]    _zz_realValue_0_350_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_350;
  wire       [5:0]    _zz_when_ArraySlice_l166_350_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_350_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_350_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_350_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_350_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_350_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_350_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_351;
  wire       [7:0]    _zz_when_ArraySlice_l158_351_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_351_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_351_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_351;
  wire       [4:0]    _zz_when_ArraySlice_l159_351_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_351_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_351_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_351_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_351_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_351_6;
  wire       [7:0]    _zz__zz_realValue_0_351;
  wire       [7:0]    _zz__zz_realValue_0_351_1;
  wire       [7:0]    _zz_realValue_0_351_1;
  wire       [7:0]    _zz_realValue_0_351_2;
  wire       [7:0]    _zz_realValue_0_351_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_351;
  wire       [4:0]    _zz_when_ArraySlice_l166_351_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_351_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_351_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_351_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_351_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_351_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_351_7;
  wire                _zz_when_ArraySlice_l314_5_1;
  wire                _zz_when_ArraySlice_l314_5_2;
  wire                _zz_when_ArraySlice_l314_5_3;
  wire                _zz_when_ArraySlice_l314_5_4;
  wire                _zz_when_ArraySlice_l314_5_5;
  wire                _zz_when_ArraySlice_l314_5_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_5;
  wire       [12:0]   _zz_when_ArraySlice_l318_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_5;
  wire       [7:0]    _zz_when_ArraySlice_l304_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_5_2;
  wire       [6:0]    _zz_when_ArraySlice_l304_5_3;
  wire       [12:0]   _zz_when_ArraySlice_l325_5;
  wire       [7:0]    _zz_when_ArraySlice_l325_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_6;
  wire       [7:0]    _zz_when_ArraySlice_l233_6_1;
  wire       [6:0]    _zz_when_ArraySlice_l233_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_6_3;
  reg        [6:0]    _zz_when_ArraySlice_l234_6;
  wire       [6:0]    _zz_when_ArraySlice_l234_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l234_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l234_6_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_6_valid_1_1;
  wire       [6:0]    _zz__zz_outputStreamArrayData_6_valid_1_2;
  wire       [6:0]    _zz__zz_17;
  reg                 _zz_outputStreamArrayData_6_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_6_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_6_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_6_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_6;
  wire       [6:0]    _zz_when_ArraySlice_l240_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l240_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l240_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l241_6;
  wire       [7:0]    _zz_when_ArraySlice_l241_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_16;
  wire       [7:0]    _zz_selectReadFifo_6_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_6;
  wire       [12:0]   _zz_when_ArraySlice_l244_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_6;
  wire       [6:0]    _zz_when_ArraySlice_l249_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l249_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l249_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l250_6;
  wire       [7:0]    _zz_when_ArraySlice_l250_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_6_2;
  wire       [7:0]    _zz__zz_realValue1_0_42;
  wire       [7:0]    _zz__zz_realValue1_0_42_1;
  wire       [7:0]    _zz_realValue1_0_42_1;
  wire       [7:0]    _zz_realValue1_0_42_2;
  wire       [7:0]    _zz_realValue1_0_42_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_6;
  wire       [6:0]    _zz_when_ArraySlice_l252_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_18;
  wire       [7:0]    _zz_selectReadFifo_6_19;
  wire       [7:0]    _zz_selectReadFifo_6_20;
  wire       [0:0]    _zz_selectReadFifo_6_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_352;
  wire       [7:0]    _zz_when_ArraySlice_l158_352_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_352_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_352_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_352;
  wire       [7:0]    _zz_when_ArraySlice_l159_352_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_352_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_352_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_352_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_352_5;
  wire       [7:0]    _zz__zz_realValue_0_352;
  wire       [7:0]    _zz__zz_realValue_0_352_1;
  wire       [7:0]    _zz_realValue_0_352_1;
  wire       [7:0]    _zz_realValue_0_352_2;
  wire       [7:0]    _zz_realValue_0_352_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_352;
  wire       [7:0]    _zz_when_ArraySlice_l166_352_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_352_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_352_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_352_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_352_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_352_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_353;
  wire       [7:0]    _zz_when_ArraySlice_l158_353_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_353_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_353_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_353;
  wire       [6:0]    _zz_when_ArraySlice_l159_353_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_353_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_353_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_353_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_353_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_353_6;
  wire       [7:0]    _zz__zz_realValue_0_353;
  wire       [7:0]    _zz__zz_realValue_0_353_1;
  wire       [7:0]    _zz_realValue_0_353_1;
  wire       [7:0]    _zz_realValue_0_353_2;
  wire       [7:0]    _zz_realValue_0_353_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_353;
  wire       [6:0]    _zz_when_ArraySlice_l166_353_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_353_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_353_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_353_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_353_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_353_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_353_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_354;
  wire       [7:0]    _zz_when_ArraySlice_l158_354_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_354_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_354_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_354;
  wire       [6:0]    _zz_when_ArraySlice_l159_354_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_354_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_354_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_354_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_354_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_354_6;
  wire       [7:0]    _zz__zz_realValue_0_354;
  wire       [7:0]    _zz__zz_realValue_0_354_1;
  wire       [7:0]    _zz_realValue_0_354_1;
  wire       [7:0]    _zz_realValue_0_354_2;
  wire       [7:0]    _zz_realValue_0_354_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_354;
  wire       [6:0]    _zz_when_ArraySlice_l166_354_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_354_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_354_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_354_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_354_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_354_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_354_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_355;
  wire       [7:0]    _zz_when_ArraySlice_l158_355_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_355_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_355_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_355;
  wire       [6:0]    _zz_when_ArraySlice_l159_355_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_355_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_355_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_355_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_355_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_355_6;
  wire       [7:0]    _zz__zz_realValue_0_355;
  wire       [7:0]    _zz__zz_realValue_0_355_1;
  wire       [7:0]    _zz_realValue_0_355_1;
  wire       [7:0]    _zz_realValue_0_355_2;
  wire       [7:0]    _zz_realValue_0_355_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_355;
  wire       [6:0]    _zz_when_ArraySlice_l166_355_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_355_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_355_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_355_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_355_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_355_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_355_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_356;
  wire       [7:0]    _zz_when_ArraySlice_l158_356_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_356_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_356_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_356;
  wire       [6:0]    _zz_when_ArraySlice_l159_356_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_356_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_356_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_356_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_356_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_356_6;
  wire       [7:0]    _zz__zz_realValue_0_356;
  wire       [7:0]    _zz__zz_realValue_0_356_1;
  wire       [7:0]    _zz_realValue_0_356_1;
  wire       [7:0]    _zz_realValue_0_356_2;
  wire       [7:0]    _zz_realValue_0_356_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_356;
  wire       [6:0]    _zz_when_ArraySlice_l166_356_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_356_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_356_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_356_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_356_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_356_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_356_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_357;
  wire       [7:0]    _zz_when_ArraySlice_l158_357_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_357_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_357_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_357;
  wire       [5:0]    _zz_when_ArraySlice_l159_357_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_357_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_357_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_357_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_357_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_357_6;
  wire       [7:0]    _zz__zz_realValue_0_357;
  wire       [7:0]    _zz__zz_realValue_0_357_1;
  wire       [7:0]    _zz_realValue_0_357_1;
  wire       [7:0]    _zz_realValue_0_357_2;
  wire       [7:0]    _zz_realValue_0_357_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_357;
  wire       [5:0]    _zz_when_ArraySlice_l166_357_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_357_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_357_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_357_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_357_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_357_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_357_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_358;
  wire       [7:0]    _zz_when_ArraySlice_l158_358_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_358_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_358_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_358;
  wire       [5:0]    _zz_when_ArraySlice_l159_358_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_358_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_358_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_358_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_358_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_358_6;
  wire       [7:0]    _zz__zz_realValue_0_358;
  wire       [7:0]    _zz__zz_realValue_0_358_1;
  wire       [7:0]    _zz_realValue_0_358_1;
  wire       [7:0]    _zz_realValue_0_358_2;
  wire       [7:0]    _zz_realValue_0_358_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_358;
  wire       [5:0]    _zz_when_ArraySlice_l166_358_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_358_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_358_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_358_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_358_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_358_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_358_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_359;
  wire       [7:0]    _zz_when_ArraySlice_l158_359_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_359_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_359_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_359;
  wire       [4:0]    _zz_when_ArraySlice_l159_359_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_359_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_359_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_359_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_359_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_359_6;
  wire       [7:0]    _zz__zz_realValue_0_359;
  wire       [7:0]    _zz__zz_realValue_0_359_1;
  wire       [7:0]    _zz_realValue_0_359_1;
  wire       [7:0]    _zz_realValue_0_359_2;
  wire       [7:0]    _zz_realValue_0_359_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_359;
  wire       [4:0]    _zz_when_ArraySlice_l166_359_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_359_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_359_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_359_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_359_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_359_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_359_7;
  wire                _zz_when_ArraySlice_l257_6;
  wire                _zz_when_ArraySlice_l257_6_1;
  wire                _zz_when_ArraySlice_l257_6_2;
  wire                _zz_when_ArraySlice_l257_6_3;
  wire                _zz_when_ArraySlice_l257_6_4;
  wire                _zz_when_ArraySlice_l257_6_5;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_6_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_6_7;
  wire       [6:0]    _zz_when_ArraySlice_l260_6_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_6;
  wire       [7:0]    _zz_when_ArraySlice_l263_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l263_6_4;
  wire       [7:0]    _zz_selectReadFifo_6_22;
  wire       [7:0]    _zz_selectReadFifo_6_23;
  wire       [6:0]    _zz_selectReadFifo_6_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_6;
  wire       [12:0]   _zz_when_ArraySlice_l270_6_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_6;
  wire       [6:0]    _zz_when_ArraySlice_l274_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l274_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l274_6_4;
  wire       [12:0]   _zz_when_ArraySlice_l275_6;
  wire       [7:0]    _zz_when_ArraySlice_l275_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_6_3;
  wire       [0:0]    _zz_when_ArraySlice_l275_6_4;
  wire       [7:0]    _zz__zz_realValue1_0_43;
  wire       [7:0]    _zz__zz_realValue1_0_43_1;
  wire       [7:0]    _zz_realValue1_0_43_1;
  wire       [7:0]    _zz_realValue1_0_43_2;
  wire       [7:0]    _zz_realValue1_0_43_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_6;
  wire       [6:0]    _zz_when_ArraySlice_l277_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_25;
  wire       [7:0]    _zz_selectReadFifo_6_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_360;
  wire       [7:0]    _zz_when_ArraySlice_l158_360_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_360_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_360_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_360;
  wire       [7:0]    _zz_when_ArraySlice_l159_360_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_360_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_360_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_360_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_360_5;
  wire       [7:0]    _zz__zz_realValue_0_360;
  wire       [7:0]    _zz__zz_realValue_0_360_1;
  wire       [7:0]    _zz_realValue_0_360_1;
  wire       [7:0]    _zz_realValue_0_360_2;
  wire       [7:0]    _zz_realValue_0_360_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_360;
  wire       [7:0]    _zz_when_ArraySlice_l166_360_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_360_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_360_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_360_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_360_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_360_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_361;
  wire       [7:0]    _zz_when_ArraySlice_l158_361_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_361_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_361_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_361;
  wire       [6:0]    _zz_when_ArraySlice_l159_361_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_361_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_361_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_361_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_361_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_361_6;
  wire       [7:0]    _zz__zz_realValue_0_361;
  wire       [7:0]    _zz__zz_realValue_0_361_1;
  wire       [7:0]    _zz_realValue_0_361_1;
  wire       [7:0]    _zz_realValue_0_361_2;
  wire       [7:0]    _zz_realValue_0_361_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_361;
  wire       [6:0]    _zz_when_ArraySlice_l166_361_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_361_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_361_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_361_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_361_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_361_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_361_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_362;
  wire       [7:0]    _zz_when_ArraySlice_l158_362_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_362_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_362_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_362;
  wire       [6:0]    _zz_when_ArraySlice_l159_362_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_362_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_362_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_362_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_362_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_362_6;
  wire       [7:0]    _zz__zz_realValue_0_362;
  wire       [7:0]    _zz__zz_realValue_0_362_1;
  wire       [7:0]    _zz_realValue_0_362_1;
  wire       [7:0]    _zz_realValue_0_362_2;
  wire       [7:0]    _zz_realValue_0_362_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_362;
  wire       [6:0]    _zz_when_ArraySlice_l166_362_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_362_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_362_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_362_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_362_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_362_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_362_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_363;
  wire       [7:0]    _zz_when_ArraySlice_l158_363_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_363_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_363_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_363;
  wire       [6:0]    _zz_when_ArraySlice_l159_363_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_363_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_363_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_363_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_363_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_363_6;
  wire       [7:0]    _zz__zz_realValue_0_363;
  wire       [7:0]    _zz__zz_realValue_0_363_1;
  wire       [7:0]    _zz_realValue_0_363_1;
  wire       [7:0]    _zz_realValue_0_363_2;
  wire       [7:0]    _zz_realValue_0_363_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_363;
  wire       [6:0]    _zz_when_ArraySlice_l166_363_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_363_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_363_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_363_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_363_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_363_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_363_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_364;
  wire       [7:0]    _zz_when_ArraySlice_l158_364_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_364_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_364_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_364;
  wire       [6:0]    _zz_when_ArraySlice_l159_364_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_364_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_364_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_364_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_364_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_364_6;
  wire       [7:0]    _zz__zz_realValue_0_364;
  wire       [7:0]    _zz__zz_realValue_0_364_1;
  wire       [7:0]    _zz_realValue_0_364_1;
  wire       [7:0]    _zz_realValue_0_364_2;
  wire       [7:0]    _zz_realValue_0_364_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_364;
  wire       [6:0]    _zz_when_ArraySlice_l166_364_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_364_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_364_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_364_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_364_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_364_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_364_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_365;
  wire       [7:0]    _zz_when_ArraySlice_l158_365_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_365_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_365_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_365;
  wire       [5:0]    _zz_when_ArraySlice_l159_365_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_365_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_365_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_365_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_365_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_365_6;
  wire       [7:0]    _zz__zz_realValue_0_365;
  wire       [7:0]    _zz__zz_realValue_0_365_1;
  wire       [7:0]    _zz_realValue_0_365_1;
  wire       [7:0]    _zz_realValue_0_365_2;
  wire       [7:0]    _zz_realValue_0_365_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_365;
  wire       [5:0]    _zz_when_ArraySlice_l166_365_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_365_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_365_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_365_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_365_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_365_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_365_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_366;
  wire       [7:0]    _zz_when_ArraySlice_l158_366_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_366_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_366_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_366;
  wire       [5:0]    _zz_when_ArraySlice_l159_366_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_366_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_366_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_366_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_366_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_366_6;
  wire       [7:0]    _zz__zz_realValue_0_366;
  wire       [7:0]    _zz__zz_realValue_0_366_1;
  wire       [7:0]    _zz_realValue_0_366_1;
  wire       [7:0]    _zz_realValue_0_366_2;
  wire       [7:0]    _zz_realValue_0_366_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_366;
  wire       [5:0]    _zz_when_ArraySlice_l166_366_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_366_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_366_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_366_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_366_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_366_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_366_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_367;
  wire       [7:0]    _zz_when_ArraySlice_l158_367_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_367_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_367_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_367;
  wire       [4:0]    _zz_when_ArraySlice_l159_367_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_367_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_367_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_367_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_367_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_367_6;
  wire       [7:0]    _zz__zz_realValue_0_367;
  wire       [7:0]    _zz__zz_realValue_0_367_1;
  wire       [7:0]    _zz_realValue_0_367_1;
  wire       [7:0]    _zz_realValue_0_367_2;
  wire       [7:0]    _zz_realValue_0_367_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_367;
  wire       [4:0]    _zz_when_ArraySlice_l166_367_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_367_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_367_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_367_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_367_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_367_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_367_7;
  wire                _zz_when_ArraySlice_l282_6;
  wire                _zz_when_ArraySlice_l282_6_1;
  wire                _zz_when_ArraySlice_l282_6_2;
  wire                _zz_when_ArraySlice_l282_6_3;
  wire                _zz_when_ArraySlice_l282_6_4;
  wire                _zz_when_ArraySlice_l282_6_5;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_6_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_6_7;
  wire       [6:0]    _zz_when_ArraySlice_l285_6_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_6;
  wire       [7:0]    _zz_when_ArraySlice_l288_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_6_3;
  wire       [6:0]    _zz_when_ArraySlice_l288_6_4;
  wire       [7:0]    _zz_selectReadFifo_6_27;
  wire       [7:0]    _zz_selectReadFifo_6_28;
  wire       [6:0]    _zz_selectReadFifo_6_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_6;
  wire       [12:0]   _zz_when_ArraySlice_l295_6_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_6;
  wire       [7:0]    _zz_when_ArraySlice_l306_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_6_2;
  wire       [7:0]    _zz__zz_realValue1_0_44;
  wire       [7:0]    _zz__zz_realValue1_0_44_1;
  wire       [7:0]    _zz_realValue1_0_44_1;
  wire       [7:0]    _zz_realValue1_0_44_2;
  wire       [7:0]    _zz_realValue1_0_44_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_6;
  wire       [6:0]    _zz_when_ArraySlice_l307_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_6_2;
  wire       [7:0]    _zz_selectReadFifo_6_30;
  wire       [7:0]    _zz_selectReadFifo_6_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_368;
  wire       [7:0]    _zz_when_ArraySlice_l158_368_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_368_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_368_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_368;
  wire       [7:0]    _zz_when_ArraySlice_l159_368_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_368_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_368_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_368_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_368_5;
  wire       [7:0]    _zz__zz_realValue_0_368;
  wire       [7:0]    _zz__zz_realValue_0_368_1;
  wire       [7:0]    _zz_realValue_0_368_1;
  wire       [7:0]    _zz_realValue_0_368_2;
  wire       [7:0]    _zz_realValue_0_368_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_368;
  wire       [7:0]    _zz_when_ArraySlice_l166_368_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_368_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_368_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_368_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_368_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_368_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_369;
  wire       [7:0]    _zz_when_ArraySlice_l158_369_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_369_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_369_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_369;
  wire       [6:0]    _zz_when_ArraySlice_l159_369_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_369_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_369_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_369_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_369_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_369_6;
  wire       [7:0]    _zz__zz_realValue_0_369;
  wire       [7:0]    _zz__zz_realValue_0_369_1;
  wire       [7:0]    _zz_realValue_0_369_1;
  wire       [7:0]    _zz_realValue_0_369_2;
  wire       [7:0]    _zz_realValue_0_369_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_369;
  wire       [6:0]    _zz_when_ArraySlice_l166_369_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_369_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_369_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_369_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_369_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_369_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_369_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_370;
  wire       [7:0]    _zz_when_ArraySlice_l158_370_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_370_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_370_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_370;
  wire       [6:0]    _zz_when_ArraySlice_l159_370_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_370_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_370_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_370_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_370_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_370_6;
  wire       [7:0]    _zz__zz_realValue_0_370;
  wire       [7:0]    _zz__zz_realValue_0_370_1;
  wire       [7:0]    _zz_realValue_0_370_1;
  wire       [7:0]    _zz_realValue_0_370_2;
  wire       [7:0]    _zz_realValue_0_370_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_370;
  wire       [6:0]    _zz_when_ArraySlice_l166_370_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_370_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_370_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_370_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_370_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_370_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_370_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_371;
  wire       [7:0]    _zz_when_ArraySlice_l158_371_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_371_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_371_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_371;
  wire       [6:0]    _zz_when_ArraySlice_l159_371_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_371_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_371_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_371_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_371_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_371_6;
  wire       [7:0]    _zz__zz_realValue_0_371;
  wire       [7:0]    _zz__zz_realValue_0_371_1;
  wire       [7:0]    _zz_realValue_0_371_1;
  wire       [7:0]    _zz_realValue_0_371_2;
  wire       [7:0]    _zz_realValue_0_371_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_371;
  wire       [6:0]    _zz_when_ArraySlice_l166_371_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_371_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_371_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_371_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_371_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_371_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_371_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_372;
  wire       [7:0]    _zz_when_ArraySlice_l158_372_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_372_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_372_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_372;
  wire       [6:0]    _zz_when_ArraySlice_l159_372_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_372_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_372_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_372_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_372_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_372_6;
  wire       [7:0]    _zz__zz_realValue_0_372;
  wire       [7:0]    _zz__zz_realValue_0_372_1;
  wire       [7:0]    _zz_realValue_0_372_1;
  wire       [7:0]    _zz_realValue_0_372_2;
  wire       [7:0]    _zz_realValue_0_372_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_372;
  wire       [6:0]    _zz_when_ArraySlice_l166_372_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_372_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_372_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_372_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_372_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_372_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_372_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_373;
  wire       [7:0]    _zz_when_ArraySlice_l158_373_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_373_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_373_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_373;
  wire       [5:0]    _zz_when_ArraySlice_l159_373_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_373_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_373_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_373_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_373_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_373_6;
  wire       [7:0]    _zz__zz_realValue_0_373;
  wire       [7:0]    _zz__zz_realValue_0_373_1;
  wire       [7:0]    _zz_realValue_0_373_1;
  wire       [7:0]    _zz_realValue_0_373_2;
  wire       [7:0]    _zz_realValue_0_373_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_373;
  wire       [5:0]    _zz_when_ArraySlice_l166_373_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_373_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_373_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_373_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_373_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_373_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_373_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_374;
  wire       [7:0]    _zz_when_ArraySlice_l158_374_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_374_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_374_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_374;
  wire       [5:0]    _zz_when_ArraySlice_l159_374_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_374_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_374_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_374_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_374_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_374_6;
  wire       [7:0]    _zz__zz_realValue_0_374;
  wire       [7:0]    _zz__zz_realValue_0_374_1;
  wire       [7:0]    _zz_realValue_0_374_1;
  wire       [7:0]    _zz_realValue_0_374_2;
  wire       [7:0]    _zz_realValue_0_374_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_374;
  wire       [5:0]    _zz_when_ArraySlice_l166_374_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_374_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_374_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_374_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_374_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_374_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_374_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_375;
  wire       [7:0]    _zz_when_ArraySlice_l158_375_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_375_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_375_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_375;
  wire       [4:0]    _zz_when_ArraySlice_l159_375_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_375_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_375_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_375_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_375_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_375_6;
  wire       [7:0]    _zz__zz_realValue_0_375;
  wire       [7:0]    _zz__zz_realValue_0_375_1;
  wire       [7:0]    _zz_realValue_0_375_1;
  wire       [7:0]    _zz_realValue_0_375_2;
  wire       [7:0]    _zz_realValue_0_375_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_375;
  wire       [4:0]    _zz_when_ArraySlice_l166_375_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_375_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_375_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_375_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_375_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_375_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_375_7;
  wire                _zz_when_ArraySlice_l314_6;
  wire                _zz_when_ArraySlice_l314_6_1;
  wire                _zz_when_ArraySlice_l314_6_2;
  wire                _zz_when_ArraySlice_l314_6_3;
  wire                _zz_when_ArraySlice_l314_6_4;
  wire                _zz_when_ArraySlice_l314_6_5;
  wire       [12:0]   _zz_when_ArraySlice_l318_6;
  wire       [12:0]   _zz_when_ArraySlice_l318_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_6;
  wire       [7:0]    _zz_when_ArraySlice_l304_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_6_2;
  wire       [6:0]    _zz_when_ArraySlice_l304_6_3;
  wire       [12:0]   _zz_when_ArraySlice_l325_6;
  wire       [7:0]    _zz_when_ArraySlice_l325_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_7;
  wire       [7:0]    _zz_when_ArraySlice_l233_7_1;
  wire       [6:0]    _zz_when_ArraySlice_l233_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l233_7_3;
  reg        [6:0]    _zz_when_ArraySlice_l234_7;
  wire       [6:0]    _zz_when_ArraySlice_l234_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l234_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l234_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l234_7_4;
  wire       [7:0]    _zz__zz_outputStreamArrayData_7_valid_1_1;
  wire       [6:0]    _zz__zz_outputStreamArrayData_7_valid_1_2;
  wire       [6:0]    _zz__zz_18;
  reg                 _zz_outputStreamArrayData_7_valid_4;
  wire       [6:0]    _zz_outputStreamArrayData_7_valid_5;
  reg        [31:0]   _zz_outputStreamArrayData_7_payload_2;
  wire       [6:0]    _zz_outputStreamArrayData_7_payload_3;
  reg        [6:0]    _zz_when_ArraySlice_l240_7;
  wire       [6:0]    _zz_when_ArraySlice_l240_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l240_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l240_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l240_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l241_7;
  wire       [7:0]    _zz_when_ArraySlice_l241_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l241_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_16;
  wire       [7:0]    _zz_selectReadFifo_7_17;
  wire       [12:0]   _zz_when_ArraySlice_l244_7;
  wire       [12:0]   _zz_when_ArraySlice_l244_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l249_7;
  wire       [6:0]    _zz_when_ArraySlice_l249_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l249_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l249_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l249_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l250_7;
  wire       [7:0]    _zz_when_ArraySlice_l250_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l250_7_2;
  wire       [7:0]    _zz__zz_realValue1_0_45;
  wire       [7:0]    _zz__zz_realValue1_0_45_1;
  wire       [7:0]    _zz_realValue1_0_45_1;
  wire       [7:0]    _zz_realValue1_0_45_2;
  wire       [7:0]    _zz_realValue1_0_45_3;
  wire       [7:0]    _zz_when_ArraySlice_l252_7;
  wire       [6:0]    _zz_when_ArraySlice_l252_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l252_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_18;
  wire       [7:0]    _zz_selectReadFifo_7_19;
  wire       [7:0]    _zz_selectReadFifo_7_20;
  wire       [0:0]    _zz_selectReadFifo_7_21;
  wire       [7:0]    _zz_when_ArraySlice_l158_376;
  wire       [7:0]    _zz_when_ArraySlice_l158_376_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_376_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_376_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_376;
  wire       [7:0]    _zz_when_ArraySlice_l159_376_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_376_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_376_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_376_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_376_5;
  wire       [7:0]    _zz__zz_realValue_0_376;
  wire       [7:0]    _zz__zz_realValue_0_376_1;
  wire       [7:0]    _zz_realValue_0_376_1;
  wire       [7:0]    _zz_realValue_0_376_2;
  wire       [7:0]    _zz_realValue_0_376_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_376;
  wire       [7:0]    _zz_when_ArraySlice_l166_376_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_376_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_376_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_376_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_376_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_376_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_377;
  wire       [7:0]    _zz_when_ArraySlice_l158_377_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_377_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_377_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_377;
  wire       [6:0]    _zz_when_ArraySlice_l159_377_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_377_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_377_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_377_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_377_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_377_6;
  wire       [7:0]    _zz__zz_realValue_0_377;
  wire       [7:0]    _zz__zz_realValue_0_377_1;
  wire       [7:0]    _zz_realValue_0_377_1;
  wire       [7:0]    _zz_realValue_0_377_2;
  wire       [7:0]    _zz_realValue_0_377_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_377;
  wire       [6:0]    _zz_when_ArraySlice_l166_377_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_377_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_377_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_377_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_377_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_377_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_377_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_378;
  wire       [7:0]    _zz_when_ArraySlice_l158_378_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_378_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_378_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_378;
  wire       [6:0]    _zz_when_ArraySlice_l159_378_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_378_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_378_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_378_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_378_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_378_6;
  wire       [7:0]    _zz__zz_realValue_0_378;
  wire       [7:0]    _zz__zz_realValue_0_378_1;
  wire       [7:0]    _zz_realValue_0_378_1;
  wire       [7:0]    _zz_realValue_0_378_2;
  wire       [7:0]    _zz_realValue_0_378_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_378;
  wire       [6:0]    _zz_when_ArraySlice_l166_378_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_378_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_378_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_378_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_378_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_378_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_378_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_379;
  wire       [7:0]    _zz_when_ArraySlice_l158_379_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_379_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_379_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_379;
  wire       [6:0]    _zz_when_ArraySlice_l159_379_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_379_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_379_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_379_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_379_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_379_6;
  wire       [7:0]    _zz__zz_realValue_0_379;
  wire       [7:0]    _zz__zz_realValue_0_379_1;
  wire       [7:0]    _zz_realValue_0_379_1;
  wire       [7:0]    _zz_realValue_0_379_2;
  wire       [7:0]    _zz_realValue_0_379_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_379;
  wire       [6:0]    _zz_when_ArraySlice_l166_379_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_379_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_379_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_379_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_379_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_379_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_379_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_380;
  wire       [7:0]    _zz_when_ArraySlice_l158_380_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_380_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_380_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_380;
  wire       [6:0]    _zz_when_ArraySlice_l159_380_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_380_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_380_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_380_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_380_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_380_6;
  wire       [7:0]    _zz__zz_realValue_0_380;
  wire       [7:0]    _zz__zz_realValue_0_380_1;
  wire       [7:0]    _zz_realValue_0_380_1;
  wire       [7:0]    _zz_realValue_0_380_2;
  wire       [7:0]    _zz_realValue_0_380_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_380;
  wire       [6:0]    _zz_when_ArraySlice_l166_380_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_380_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_380_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_380_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_380_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_380_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_380_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_381;
  wire       [7:0]    _zz_when_ArraySlice_l158_381_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_381_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_381_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_381;
  wire       [5:0]    _zz_when_ArraySlice_l159_381_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_381_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_381_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_381_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_381_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_381_6;
  wire       [7:0]    _zz__zz_realValue_0_381;
  wire       [7:0]    _zz__zz_realValue_0_381_1;
  wire       [7:0]    _zz_realValue_0_381_1;
  wire       [7:0]    _zz_realValue_0_381_2;
  wire       [7:0]    _zz_realValue_0_381_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_381;
  wire       [5:0]    _zz_when_ArraySlice_l166_381_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_381_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_381_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_381_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_381_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_381_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_381_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_382;
  wire       [7:0]    _zz_when_ArraySlice_l158_382_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_382_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_382_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_382;
  wire       [5:0]    _zz_when_ArraySlice_l159_382_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_382_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_382_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_382_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_382_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_382_6;
  wire       [7:0]    _zz__zz_realValue_0_382;
  wire       [7:0]    _zz__zz_realValue_0_382_1;
  wire       [7:0]    _zz_realValue_0_382_1;
  wire       [7:0]    _zz_realValue_0_382_2;
  wire       [7:0]    _zz_realValue_0_382_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_382;
  wire       [5:0]    _zz_when_ArraySlice_l166_382_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_382_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_382_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_382_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_382_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_382_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_382_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_383;
  wire       [7:0]    _zz_when_ArraySlice_l158_383_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_383_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_383_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_383;
  wire       [4:0]    _zz_when_ArraySlice_l159_383_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_383_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_383_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_383_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_383_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_383_6;
  wire       [7:0]    _zz__zz_realValue_0_383;
  wire       [7:0]    _zz__zz_realValue_0_383_1;
  wire       [7:0]    _zz_realValue_0_383_1;
  wire       [7:0]    _zz_realValue_0_383_2;
  wire       [7:0]    _zz_realValue_0_383_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_383;
  wire       [4:0]    _zz_when_ArraySlice_l166_383_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_383_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_383_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_383_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_383_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_383_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_383_7;
  wire                _zz_when_ArraySlice_l257_7;
  wire                _zz_when_ArraySlice_l257_7_1;
  wire                _zz_when_ArraySlice_l257_7_2;
  wire                _zz_when_ArraySlice_l257_7_3;
  wire                _zz_when_ArraySlice_l257_7_4;
  wire                _zz_when_ArraySlice_l257_7_5;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l260_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l260_7_7;
  wire       [6:0]    _zz_when_ArraySlice_l260_7_8;
  wire       [7:0]    _zz_when_ArraySlice_l263_7;
  wire       [7:0]    _zz_when_ArraySlice_l263_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l263_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l263_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l263_7_4;
  wire       [7:0]    _zz_selectReadFifo_7_22;
  wire       [7:0]    _zz_selectReadFifo_7_23;
  wire       [6:0]    _zz_selectReadFifo_7_24;
  wire       [12:0]   _zz_when_ArraySlice_l270_7;
  wire       [12:0]   _zz_when_ArraySlice_l270_7_1;
  reg        [6:0]    _zz_when_ArraySlice_l274_7;
  wire       [6:0]    _zz_when_ArraySlice_l274_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l274_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l274_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l274_7_4;
  wire       [12:0]   _zz_when_ArraySlice_l275_7;
  wire       [7:0]    _zz_when_ArraySlice_l275_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l275_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l275_7_3;
  wire       [0:0]    _zz_when_ArraySlice_l275_7_4;
  wire       [7:0]    _zz__zz_realValue1_0_46;
  wire       [7:0]    _zz__zz_realValue1_0_46_1;
  wire       [7:0]    _zz_realValue1_0_46_1;
  wire       [7:0]    _zz_realValue1_0_46_2;
  wire       [7:0]    _zz_realValue1_0_46_3;
  wire       [7:0]    _zz_when_ArraySlice_l277_7;
  wire       [6:0]    _zz_when_ArraySlice_l277_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l277_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_25;
  wire       [7:0]    _zz_selectReadFifo_7_26;
  wire       [7:0]    _zz_when_ArraySlice_l158_384;
  wire       [7:0]    _zz_when_ArraySlice_l158_384_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_384_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_384_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_384;
  wire       [7:0]    _zz_when_ArraySlice_l159_384_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_384_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_384_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_384_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_384_5;
  wire       [7:0]    _zz__zz_realValue_0_384;
  wire       [7:0]    _zz__zz_realValue_0_384_1;
  wire       [7:0]    _zz_realValue_0_384_1;
  wire       [7:0]    _zz_realValue_0_384_2;
  wire       [7:0]    _zz_realValue_0_384_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_384;
  wire       [7:0]    _zz_when_ArraySlice_l166_384_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_384_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_384_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_384_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_384_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_384_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_385;
  wire       [7:0]    _zz_when_ArraySlice_l158_385_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_385_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_385_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_385;
  wire       [6:0]    _zz_when_ArraySlice_l159_385_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_385_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_385_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_385_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_385_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_385_6;
  wire       [7:0]    _zz__zz_realValue_0_385;
  wire       [7:0]    _zz__zz_realValue_0_385_1;
  wire       [7:0]    _zz_realValue_0_385_1;
  wire       [7:0]    _zz_realValue_0_385_2;
  wire       [7:0]    _zz_realValue_0_385_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_385;
  wire       [6:0]    _zz_when_ArraySlice_l166_385_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_385_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_385_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_385_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_385_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_385_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_385_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_386;
  wire       [7:0]    _zz_when_ArraySlice_l158_386_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_386_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_386_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_386;
  wire       [6:0]    _zz_when_ArraySlice_l159_386_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_386_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_386_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_386_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_386_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_386_6;
  wire       [7:0]    _zz__zz_realValue_0_386;
  wire       [7:0]    _zz__zz_realValue_0_386_1;
  wire       [7:0]    _zz_realValue_0_386_1;
  wire       [7:0]    _zz_realValue_0_386_2;
  wire       [7:0]    _zz_realValue_0_386_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_386;
  wire       [6:0]    _zz_when_ArraySlice_l166_386_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_386_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_386_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_386_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_386_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_386_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_386_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_387;
  wire       [7:0]    _zz_when_ArraySlice_l158_387_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_387_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_387_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_387;
  wire       [6:0]    _zz_when_ArraySlice_l159_387_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_387_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_387_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_387_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_387_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_387_6;
  wire       [7:0]    _zz__zz_realValue_0_387;
  wire       [7:0]    _zz__zz_realValue_0_387_1;
  wire       [7:0]    _zz_realValue_0_387_1;
  wire       [7:0]    _zz_realValue_0_387_2;
  wire       [7:0]    _zz_realValue_0_387_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_387;
  wire       [6:0]    _zz_when_ArraySlice_l166_387_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_387_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_387_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_387_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_387_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_387_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_387_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_388;
  wire       [7:0]    _zz_when_ArraySlice_l158_388_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_388_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_388_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_388;
  wire       [6:0]    _zz_when_ArraySlice_l159_388_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_388_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_388_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_388_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_388_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_388_6;
  wire       [7:0]    _zz__zz_realValue_0_388;
  wire       [7:0]    _zz__zz_realValue_0_388_1;
  wire       [7:0]    _zz_realValue_0_388_1;
  wire       [7:0]    _zz_realValue_0_388_2;
  wire       [7:0]    _zz_realValue_0_388_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_388;
  wire       [6:0]    _zz_when_ArraySlice_l166_388_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_388_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_388_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_388_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_388_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_388_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_388_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_389;
  wire       [7:0]    _zz_when_ArraySlice_l158_389_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_389_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_389_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_389;
  wire       [5:0]    _zz_when_ArraySlice_l159_389_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_389_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_389_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_389_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_389_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_389_6;
  wire       [7:0]    _zz__zz_realValue_0_389;
  wire       [7:0]    _zz__zz_realValue_0_389_1;
  wire       [7:0]    _zz_realValue_0_389_1;
  wire       [7:0]    _zz_realValue_0_389_2;
  wire       [7:0]    _zz_realValue_0_389_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_389;
  wire       [5:0]    _zz_when_ArraySlice_l166_389_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_389_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_389_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_389_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_389_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_389_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_389_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_390;
  wire       [7:0]    _zz_when_ArraySlice_l158_390_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_390_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_390_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_390;
  wire       [5:0]    _zz_when_ArraySlice_l159_390_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_390_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_390_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_390_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_390_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_390_6;
  wire       [7:0]    _zz__zz_realValue_0_390;
  wire       [7:0]    _zz__zz_realValue_0_390_1;
  wire       [7:0]    _zz_realValue_0_390_1;
  wire       [7:0]    _zz_realValue_0_390_2;
  wire       [7:0]    _zz_realValue_0_390_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_390;
  wire       [5:0]    _zz_when_ArraySlice_l166_390_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_390_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_390_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_390_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_390_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_390_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_390_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_391;
  wire       [7:0]    _zz_when_ArraySlice_l158_391_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_391_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_391_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_391;
  wire       [4:0]    _zz_when_ArraySlice_l159_391_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_391_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_391_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_391_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_391_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_391_6;
  wire       [7:0]    _zz__zz_realValue_0_391;
  wire       [7:0]    _zz__zz_realValue_0_391_1;
  wire       [7:0]    _zz_realValue_0_391_1;
  wire       [7:0]    _zz_realValue_0_391_2;
  wire       [7:0]    _zz_realValue_0_391_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_391;
  wire       [4:0]    _zz_when_ArraySlice_l166_391_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_391_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_391_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_391_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_391_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_391_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_391_7;
  wire                _zz_when_ArraySlice_l282_7;
  wire                _zz_when_ArraySlice_l282_7_1;
  wire                _zz_when_ArraySlice_l282_7_2;
  wire                _zz_when_ArraySlice_l282_7_3;
  wire                _zz_when_ArraySlice_l282_7_4;
  wire                _zz_when_ArraySlice_l282_7_5;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_3;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_4;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_5;
  wire       [6:0]    _zz_when_ArraySlice_l285_7_6;
  wire       [7:0]    _zz_when_ArraySlice_l285_7_7;
  wire       [6:0]    _zz_when_ArraySlice_l285_7_8;
  wire       [7:0]    _zz_when_ArraySlice_l288_7;
  wire       [7:0]    _zz_when_ArraySlice_l288_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l288_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l288_7_3;
  wire       [6:0]    _zz_when_ArraySlice_l288_7_4;
  wire       [7:0]    _zz_selectReadFifo_7_27;
  wire       [7:0]    _zz_selectReadFifo_7_28;
  wire       [6:0]    _zz_selectReadFifo_7_29;
  wire       [12:0]   _zz_when_ArraySlice_l295_7;
  wire       [12:0]   _zz_when_ArraySlice_l295_7_1;
  wire       [12:0]   _zz_when_ArraySlice_l306_7;
  wire       [7:0]    _zz_when_ArraySlice_l306_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l306_7_2;
  wire       [7:0]    _zz__zz_realValue1_0_47;
  wire       [7:0]    _zz__zz_realValue1_0_47_1;
  wire       [7:0]    _zz_realValue1_0_47_1;
  wire       [7:0]    _zz_realValue1_0_47_2;
  wire       [7:0]    _zz_realValue1_0_47_3;
  wire       [7:0]    _zz_when_ArraySlice_l307_7;
  wire       [6:0]    _zz_when_ArraySlice_l307_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l307_7_2;
  wire       [7:0]    _zz_selectReadFifo_7_30;
  wire       [7:0]    _zz_selectReadFifo_7_31;
  wire       [7:0]    _zz_when_ArraySlice_l158_392;
  wire       [7:0]    _zz_when_ArraySlice_l158_392_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_392_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_392_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_392;
  wire       [7:0]    _zz_when_ArraySlice_l159_392_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_392_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_392_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_392_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_392_5;
  wire       [7:0]    _zz__zz_realValue_0_392;
  wire       [7:0]    _zz__zz_realValue_0_392_1;
  wire       [7:0]    _zz_realValue_0_392_1;
  wire       [7:0]    _zz_realValue_0_392_2;
  wire       [7:0]    _zz_realValue_0_392_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_392;
  wire       [7:0]    _zz_when_ArraySlice_l166_392_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_392_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_392_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_392_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_392_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_392_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_393;
  wire       [7:0]    _zz_when_ArraySlice_l158_393_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_393_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_393_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_393;
  wire       [6:0]    _zz_when_ArraySlice_l159_393_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_393_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_393_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_393_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_393_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_393_6;
  wire       [7:0]    _zz__zz_realValue_0_393;
  wire       [7:0]    _zz__zz_realValue_0_393_1;
  wire       [7:0]    _zz_realValue_0_393_1;
  wire       [7:0]    _zz_realValue_0_393_2;
  wire       [7:0]    _zz_realValue_0_393_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_393;
  wire       [6:0]    _zz_when_ArraySlice_l166_393_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_393_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_393_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_393_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_393_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_393_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_393_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_394;
  wire       [7:0]    _zz_when_ArraySlice_l158_394_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_394_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_394_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_394;
  wire       [6:0]    _zz_when_ArraySlice_l159_394_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_394_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_394_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_394_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_394_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_394_6;
  wire       [7:0]    _zz__zz_realValue_0_394;
  wire       [7:0]    _zz__zz_realValue_0_394_1;
  wire       [7:0]    _zz_realValue_0_394_1;
  wire       [7:0]    _zz_realValue_0_394_2;
  wire       [7:0]    _zz_realValue_0_394_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_394;
  wire       [6:0]    _zz_when_ArraySlice_l166_394_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_394_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_394_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_394_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_394_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_394_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_394_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_395;
  wire       [7:0]    _zz_when_ArraySlice_l158_395_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_395_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_395_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_395;
  wire       [6:0]    _zz_when_ArraySlice_l159_395_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_395_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_395_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_395_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_395_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_395_6;
  wire       [7:0]    _zz__zz_realValue_0_395;
  wire       [7:0]    _zz__zz_realValue_0_395_1;
  wire       [7:0]    _zz_realValue_0_395_1;
  wire       [7:0]    _zz_realValue_0_395_2;
  wire       [7:0]    _zz_realValue_0_395_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_395;
  wire       [6:0]    _zz_when_ArraySlice_l166_395_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_395_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_395_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_395_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_395_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_395_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_395_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_396;
  wire       [7:0]    _zz_when_ArraySlice_l158_396_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_396_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_396_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_396;
  wire       [6:0]    _zz_when_ArraySlice_l159_396_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_396_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_396_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_396_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_396_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_396_6;
  wire       [7:0]    _zz__zz_realValue_0_396;
  wire       [7:0]    _zz__zz_realValue_0_396_1;
  wire       [7:0]    _zz_realValue_0_396_1;
  wire       [7:0]    _zz_realValue_0_396_2;
  wire       [7:0]    _zz_realValue_0_396_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_396;
  wire       [6:0]    _zz_when_ArraySlice_l166_396_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_396_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_396_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_396_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_396_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_396_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_396_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_397;
  wire       [7:0]    _zz_when_ArraySlice_l158_397_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_397_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_397_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_397;
  wire       [5:0]    _zz_when_ArraySlice_l159_397_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_397_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_397_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_397_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_397_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_397_6;
  wire       [7:0]    _zz__zz_realValue_0_397;
  wire       [7:0]    _zz__zz_realValue_0_397_1;
  wire       [7:0]    _zz_realValue_0_397_1;
  wire       [7:0]    _zz_realValue_0_397_2;
  wire       [7:0]    _zz_realValue_0_397_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_397;
  wire       [5:0]    _zz_when_ArraySlice_l166_397_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_397_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_397_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_397_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_397_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_397_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_397_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_398;
  wire       [7:0]    _zz_when_ArraySlice_l158_398_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_398_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_398_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_398;
  wire       [5:0]    _zz_when_ArraySlice_l159_398_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_398_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_398_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_398_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_398_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_398_6;
  wire       [7:0]    _zz__zz_realValue_0_398;
  wire       [7:0]    _zz__zz_realValue_0_398_1;
  wire       [7:0]    _zz_realValue_0_398_1;
  wire       [7:0]    _zz_realValue_0_398_2;
  wire       [7:0]    _zz_realValue_0_398_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_398;
  wire       [5:0]    _zz_when_ArraySlice_l166_398_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_398_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_398_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_398_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_398_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_398_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_398_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_399;
  wire       [7:0]    _zz_when_ArraySlice_l158_399_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_399_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_399_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_399;
  wire       [4:0]    _zz_when_ArraySlice_l159_399_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_399_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_399_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_399_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_399_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_399_6;
  wire       [7:0]    _zz__zz_realValue_0_399;
  wire       [7:0]    _zz__zz_realValue_0_399_1;
  wire       [7:0]    _zz_realValue_0_399_1;
  wire       [7:0]    _zz_realValue_0_399_2;
  wire       [7:0]    _zz_realValue_0_399_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_399;
  wire       [4:0]    _zz_when_ArraySlice_l166_399_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_399_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_399_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_399_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_399_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_399_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_399_7;
  wire                _zz_when_ArraySlice_l314_7;
  wire                _zz_when_ArraySlice_l314_7_1;
  wire                _zz_when_ArraySlice_l314_7_2;
  wire                _zz_when_ArraySlice_l314_7_3;
  wire                _zz_when_ArraySlice_l314_7_4;
  wire                _zz_when_ArraySlice_l314_7_5;
  wire       [12:0]   _zz_when_ArraySlice_l318_7;
  wire       [12:0]   _zz_when_ArraySlice_l318_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_7;
  wire       [7:0]    _zz_when_ArraySlice_l304_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l304_7_2;
  wire       [6:0]    _zz_when_ArraySlice_l304_7_3;
  wire       [12:0]   _zz_when_ArraySlice_l325_7;
  wire       [7:0]    _zz_when_ArraySlice_l325_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l325_7_2;
  wire       [7:0]    _zz_when_ArraySlice_l182;
  wire       [7:0]    _zz_when_ArraySlice_l182_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_1_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_1_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_1_3;
  wire       [7:0]    _zz_when_ArraySlice_l182_2_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_2_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_2_3;
  wire       [7:0]    _zz_when_ArraySlice_l182_3;
  wire       [7:0]    _zz_when_ArraySlice_l182_3_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_3_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_4;
  wire       [7:0]    _zz_when_ArraySlice_l182_4_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_4_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_5;
  wire       [7:0]    _zz_when_ArraySlice_l182_5_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_5_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_6;
  wire       [7:0]    _zz_when_ArraySlice_l182_6_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_6_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_7;
  wire       [7:0]    _zz_when_ArraySlice_l182_7_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_7_2;
  wire                _zz_when_ArraySlice_l336_8;
  wire                _zz_when_ArraySlice_l336_9;
  reg        [6:0]    _zz_when_ArraySlice_l337;
  reg                 _zz_inputStreamArrayData_ready_1;
  reg        [6:0]    _zz_when_ArraySlice_l341;
  wire       [6:0]    _zz_when_ArraySlice_l341_1;
  wire       [6:0]    _zz_when_ArraySlice_l342;
  wire       [7:0]    _zz_when_ArraySlice_l158_400;
  wire       [7:0]    _zz_when_ArraySlice_l158_400_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_400_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_400_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_400;
  wire       [7:0]    _zz_when_ArraySlice_l159_400_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_400_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_400_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_400_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_400_5;
  wire       [7:0]    _zz__zz_realValue_0_400;
  wire       [7:0]    _zz__zz_realValue_0_400_1;
  wire       [7:0]    _zz_realValue_0_400_1;
  wire       [7:0]    _zz_realValue_0_400_2;
  wire       [7:0]    _zz_realValue_0_400_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_400;
  wire       [7:0]    _zz_when_ArraySlice_l166_400_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_400_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_400_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_400_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_400_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_400_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_401;
  wire       [7:0]    _zz_when_ArraySlice_l158_401_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_401_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_401_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_401;
  wire       [6:0]    _zz_when_ArraySlice_l159_401_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_401_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_401_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_401_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_401_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_401_6;
  wire       [7:0]    _zz__zz_realValue_0_401;
  wire       [7:0]    _zz__zz_realValue_0_401_1;
  wire       [7:0]    _zz_realValue_0_401_1;
  wire       [7:0]    _zz_realValue_0_401_2;
  wire       [7:0]    _zz_realValue_0_401_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_401;
  wire       [6:0]    _zz_when_ArraySlice_l166_401_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_401_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_401_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_401_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_401_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_401_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_401_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_402;
  wire       [7:0]    _zz_when_ArraySlice_l158_402_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_402_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_402_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_402;
  wire       [6:0]    _zz_when_ArraySlice_l159_402_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_402_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_402_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_402_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_402_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_402_6;
  wire       [7:0]    _zz__zz_realValue_0_402;
  wire       [7:0]    _zz__zz_realValue_0_402_1;
  wire       [7:0]    _zz_realValue_0_402_1;
  wire       [7:0]    _zz_realValue_0_402_2;
  wire       [7:0]    _zz_realValue_0_402_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_402;
  wire       [6:0]    _zz_when_ArraySlice_l166_402_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_402_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_402_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_402_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_402_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_402_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_402_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_403;
  wire       [7:0]    _zz_when_ArraySlice_l158_403_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_403_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_403_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_403;
  wire       [6:0]    _zz_when_ArraySlice_l159_403_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_403_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_403_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_403_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_403_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_403_6;
  wire       [7:0]    _zz__zz_realValue_0_403;
  wire       [7:0]    _zz__zz_realValue_0_403_1;
  wire       [7:0]    _zz_realValue_0_403_1;
  wire       [7:0]    _zz_realValue_0_403_2;
  wire       [7:0]    _zz_realValue_0_403_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_403;
  wire       [6:0]    _zz_when_ArraySlice_l166_403_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_403_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_403_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_403_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_403_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_403_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_403_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_404;
  wire       [7:0]    _zz_when_ArraySlice_l158_404_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_404_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_404_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_404;
  wire       [6:0]    _zz_when_ArraySlice_l159_404_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_404_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_404_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_404_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_404_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_404_6;
  wire       [7:0]    _zz__zz_realValue_0_404;
  wire       [7:0]    _zz__zz_realValue_0_404_1;
  wire       [7:0]    _zz_realValue_0_404_1;
  wire       [7:0]    _zz_realValue_0_404_2;
  wire       [7:0]    _zz_realValue_0_404_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_404;
  wire       [6:0]    _zz_when_ArraySlice_l166_404_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_404_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_404_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_404_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_404_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_404_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_404_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_405;
  wire       [7:0]    _zz_when_ArraySlice_l158_405_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_405_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_405_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_405;
  wire       [5:0]    _zz_when_ArraySlice_l159_405_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_405_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_405_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_405_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_405_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_405_6;
  wire       [7:0]    _zz__zz_realValue_0_405;
  wire       [7:0]    _zz__zz_realValue_0_405_1;
  wire       [7:0]    _zz_realValue_0_405_1;
  wire       [7:0]    _zz_realValue_0_405_2;
  wire       [7:0]    _zz_realValue_0_405_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_405;
  wire       [5:0]    _zz_when_ArraySlice_l166_405_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_405_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_405_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_405_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_405_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_405_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_405_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_406;
  wire       [7:0]    _zz_when_ArraySlice_l158_406_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_406_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_406_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_406;
  wire       [5:0]    _zz_when_ArraySlice_l159_406_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_406_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_406_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_406_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_406_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_406_6;
  wire       [7:0]    _zz__zz_realValue_0_406;
  wire       [7:0]    _zz__zz_realValue_0_406_1;
  wire       [7:0]    _zz_realValue_0_406_1;
  wire       [7:0]    _zz_realValue_0_406_2;
  wire       [7:0]    _zz_realValue_0_406_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_406;
  wire       [5:0]    _zz_when_ArraySlice_l166_406_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_406_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_406_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_406_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_406_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_406_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_406_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_407;
  wire       [7:0]    _zz_when_ArraySlice_l158_407_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_407_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_407_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_407;
  wire       [4:0]    _zz_when_ArraySlice_l159_407_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_407_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_407_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_407_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_407_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_407_6;
  wire       [7:0]    _zz__zz_realValue_0_407;
  wire       [7:0]    _zz__zz_realValue_0_407_1;
  wire       [7:0]    _zz_realValue_0_407_1;
  wire       [7:0]    _zz_realValue_0_407_2;
  wire       [7:0]    _zz_realValue_0_407_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_407;
  wire       [4:0]    _zz_when_ArraySlice_l166_407_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_407_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_407_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_407_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_407_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_407_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_407_7;
  wire                _zz_when_ArraySlice_l353;
  wire                _zz_when_ArraySlice_l353_1;
  wire                _zz_when_ArraySlice_l353_2;
  wire                _zz_when_ArraySlice_l353_3;
  wire                _zz_when_ArraySlice_l353_4;
  wire                _zz_when_ArraySlice_l353_5;
  wire       [7:0]    _zz_when_ArraySlice_l158_408;
  wire       [7:0]    _zz_when_ArraySlice_l158_408_1;
  wire       [3:0]    _zz_when_ArraySlice_l158_408_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_408_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_408;
  wire       [7:0]    _zz_when_ArraySlice_l159_408_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_408_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_408_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_408_4;
  wire       [3:0]    _zz_when_ArraySlice_l159_408_5;
  wire       [7:0]    _zz__zz_realValue_0_408;
  wire       [7:0]    _zz__zz_realValue_0_408_1;
  wire       [7:0]    _zz_realValue_0_408_1;
  wire       [7:0]    _zz_realValue_0_408_2;
  wire       [7:0]    _zz_realValue_0_408_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_408;
  wire       [7:0]    _zz_when_ArraySlice_l166_408_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_408_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_408_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_408_4;
  wire       [3:0]    _zz_when_ArraySlice_l166_408_5;
  wire       [7:0]    _zz_when_ArraySlice_l166_408_6;
  wire       [7:0]    _zz_when_ArraySlice_l158_409;
  wire       [7:0]    _zz_when_ArraySlice_l158_409_1;
  wire       [4:0]    _zz_when_ArraySlice_l158_409_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_409_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_409;
  wire       [6:0]    _zz_when_ArraySlice_l159_409_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_409_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_409_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_409_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_409_5;
  wire       [4:0]    _zz_when_ArraySlice_l159_409_6;
  wire       [7:0]    _zz__zz_realValue_0_409;
  wire       [7:0]    _zz__zz_realValue_0_409_1;
  wire       [7:0]    _zz_realValue_0_409_1;
  wire       [7:0]    _zz_realValue_0_409_2;
  wire       [7:0]    _zz_realValue_0_409_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_409;
  wire       [6:0]    _zz_when_ArraySlice_l166_409_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_409_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_409_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_409_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_409_5;
  wire       [4:0]    _zz_when_ArraySlice_l166_409_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_409_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_410;
  wire       [7:0]    _zz_when_ArraySlice_l158_410_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_410_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_410_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_410;
  wire       [6:0]    _zz_when_ArraySlice_l159_410_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_410_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_410_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_410_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_410_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_410_6;
  wire       [7:0]    _zz__zz_realValue_0_410;
  wire       [7:0]    _zz__zz_realValue_0_410_1;
  wire       [7:0]    _zz_realValue_0_410_1;
  wire       [7:0]    _zz_realValue_0_410_2;
  wire       [7:0]    _zz_realValue_0_410_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_410;
  wire       [6:0]    _zz_when_ArraySlice_l166_410_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_410_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_410_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_410_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_410_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_410_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_410_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_411;
  wire       [7:0]    _zz_when_ArraySlice_l158_411_1;
  wire       [5:0]    _zz_when_ArraySlice_l158_411_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_411_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_411;
  wire       [6:0]    _zz_when_ArraySlice_l159_411_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_411_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_411_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_411_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_411_5;
  wire       [5:0]    _zz_when_ArraySlice_l159_411_6;
  wire       [7:0]    _zz__zz_realValue_0_411;
  wire       [7:0]    _zz__zz_realValue_0_411_1;
  wire       [7:0]    _zz_realValue_0_411_1;
  wire       [7:0]    _zz_realValue_0_411_2;
  wire       [7:0]    _zz_realValue_0_411_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_411;
  wire       [6:0]    _zz_when_ArraySlice_l166_411_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_411_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_411_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_411_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_411_5;
  wire       [5:0]    _zz_when_ArraySlice_l166_411_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_411_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_412;
  wire       [7:0]    _zz_when_ArraySlice_l158_412_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_412_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_412_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_412;
  wire       [6:0]    _zz_when_ArraySlice_l159_412_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_412_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_412_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_412_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_412_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_412_6;
  wire       [7:0]    _zz__zz_realValue_0_412;
  wire       [7:0]    _zz__zz_realValue_0_412_1;
  wire       [7:0]    _zz_realValue_0_412_1;
  wire       [7:0]    _zz_realValue_0_412_2;
  wire       [7:0]    _zz_realValue_0_412_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_412;
  wire       [6:0]    _zz_when_ArraySlice_l166_412_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_412_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_412_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_412_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_412_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_412_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_412_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_413;
  wire       [7:0]    _zz_when_ArraySlice_l158_413_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_413_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_413_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_413;
  wire       [5:0]    _zz_when_ArraySlice_l159_413_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_413_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_413_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_413_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_413_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_413_6;
  wire       [7:0]    _zz__zz_realValue_0_413;
  wire       [7:0]    _zz__zz_realValue_0_413_1;
  wire       [7:0]    _zz_realValue_0_413_1;
  wire       [7:0]    _zz_realValue_0_413_2;
  wire       [7:0]    _zz_realValue_0_413_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_413;
  wire       [5:0]    _zz_when_ArraySlice_l166_413_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_413_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_413_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_413_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_413_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_413_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_413_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_414;
  wire       [7:0]    _zz_when_ArraySlice_l158_414_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_414_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_414_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_414;
  wire       [5:0]    _zz_when_ArraySlice_l159_414_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_414_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_414_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_414_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_414_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_414_6;
  wire       [7:0]    _zz__zz_realValue_0_414;
  wire       [7:0]    _zz__zz_realValue_0_414_1;
  wire       [7:0]    _zz_realValue_0_414_1;
  wire       [7:0]    _zz_realValue_0_414_2;
  wire       [7:0]    _zz_realValue_0_414_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_414;
  wire       [5:0]    _zz_when_ArraySlice_l166_414_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_414_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_414_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_414_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_414_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_414_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_414_7;
  wire       [7:0]    _zz_when_ArraySlice_l158_415;
  wire       [7:0]    _zz_when_ArraySlice_l158_415_1;
  wire       [6:0]    _zz_when_ArraySlice_l158_415_2;
  wire       [7:0]    _zz_when_ArraySlice_l158_415_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_415;
  wire       [4:0]    _zz_when_ArraySlice_l159_415_1;
  wire       [7:0]    _zz_when_ArraySlice_l159_415_2;
  wire       [7:0]    _zz_when_ArraySlice_l159_415_3;
  wire       [7:0]    _zz_when_ArraySlice_l159_415_4;
  wire       [7:0]    _zz_when_ArraySlice_l159_415_5;
  wire       [6:0]    _zz_when_ArraySlice_l159_415_6;
  wire       [7:0]    _zz__zz_realValue_0_415;
  wire       [7:0]    _zz__zz_realValue_0_415_1;
  wire       [7:0]    _zz_realValue_0_415_1;
  wire       [7:0]    _zz_realValue_0_415_2;
  wire       [7:0]    _zz_realValue_0_415_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_415;
  wire       [4:0]    _zz_when_ArraySlice_l166_415_1;
  wire       [7:0]    _zz_when_ArraySlice_l166_415_2;
  wire       [7:0]    _zz_when_ArraySlice_l166_415_3;
  wire       [7:0]    _zz_when_ArraySlice_l166_415_4;
  wire       [7:0]    _zz_when_ArraySlice_l166_415_5;
  wire       [6:0]    _zz_when_ArraySlice_l166_415_6;
  wire       [7:0]    _zz_when_ArraySlice_l166_415_7;
  wire       [7:0]    _zz_when_ArraySlice_l182_8;
  wire       [7:0]    _zz_when_ArraySlice_l182_8_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_8_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_9;
  wire       [7:0]    _zz_when_ArraySlice_l182_9_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_9_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_10;
  wire       [7:0]    _zz_when_ArraySlice_l182_10_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_10_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_11;
  wire       [7:0]    _zz_when_ArraySlice_l182_11_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_11_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_12;
  wire       [7:0]    _zz_when_ArraySlice_l182_12_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_12_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_13;
  wire       [7:0]    _zz_when_ArraySlice_l182_13_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_13_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_14;
  wire       [7:0]    _zz_when_ArraySlice_l182_14_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_14_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_15;
  wire       [7:0]    _zz_when_ArraySlice_l182_15_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_15_2;
  wire                _zz_when_ArraySlice_l357_8;
  wire                _zz_when_ArraySlice_l357_9;
  wire                _zz_when_ArraySlice_l357_10;
  wire                _zz_when_ArraySlice_l357_11;
  wire                _zz_when_ArraySlice_l357_12;
  wire                _zz_when_ArraySlice_l357_13;
  wire                _zz_when_ArraySlice_l357_14;
  wire                _zz_when_ArraySlice_l357_15;
  wire                _zz_when_ArraySlice_l357_16;
  wire                _zz_when_ArraySlice_l357_17;
  wire                _zz_when_ArraySlice_l357_18;
  wire                _zz_when_ArraySlice_l357_19;
  wire                _zz_when_ArraySlice_l357_20;
  wire                _zz_when_ArraySlice_l357_21;
  wire                _zz_when_ArraySlice_l357_22;
  wire                _zz_when_ArraySlice_l357_23;
  wire                _zz_when_ArraySlice_l357_24;
  wire                _zz_when_ArraySlice_l357_25;
  wire       [7:0]    _zz_when_ArraySlice_l182_16;
  wire       [7:0]    _zz_when_ArraySlice_l182_16_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_16_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_17;
  wire       [7:0]    _zz_when_ArraySlice_l182_17_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_17_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_18;
  wire       [7:0]    _zz_when_ArraySlice_l182_18_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_18_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_19;
  wire       [7:0]    _zz_when_ArraySlice_l182_19_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_19_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_20;
  wire       [7:0]    _zz_when_ArraySlice_l182_20_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_20_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_21;
  wire       [7:0]    _zz_when_ArraySlice_l182_21_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_21_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_22;
  wire       [7:0]    _zz_when_ArraySlice_l182_22_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_22_2;
  wire       [7:0]    _zz_when_ArraySlice_l182_23;
  wire       [7:0]    _zz_when_ArraySlice_l182_23_1;
  wire       [7:0]    _zz_when_ArraySlice_l182_23_2;
  wire       [31:0]   arrayDataType;
  reg        [6:0]    wReg;
  reg        [6:0]    hReg;
  reg        [3:0]    aReg;
  reg        [3:0]    bReg;
  reg                 handshakeTimes_0_willIncrement;
  reg                 handshakeTimes_0_willClear;
  reg        [12:0]   handshakeTimes_0_valueNext;
  reg        [12:0]   handshakeTimes_0_value;
  wire                handshakeTimes_0_willOverflowIfInc;
  wire                handshakeTimes_0_willOverflow;
  reg                 handshakeTimes_1_willIncrement;
  reg                 handshakeTimes_1_willClear;
  reg        [12:0]   handshakeTimes_1_valueNext;
  reg        [12:0]   handshakeTimes_1_value;
  wire                handshakeTimes_1_willOverflowIfInc;
  wire                handshakeTimes_1_willOverflow;
  reg                 handshakeTimes_2_willIncrement;
  reg                 handshakeTimes_2_willClear;
  reg        [12:0]   handshakeTimes_2_valueNext;
  reg        [12:0]   handshakeTimes_2_value;
  wire                handshakeTimes_2_willOverflowIfInc;
  wire                handshakeTimes_2_willOverflow;
  reg                 handshakeTimes_3_willIncrement;
  reg                 handshakeTimes_3_willClear;
  reg        [12:0]   handshakeTimes_3_valueNext;
  reg        [12:0]   handshakeTimes_3_value;
  wire                handshakeTimes_3_willOverflowIfInc;
  wire                handshakeTimes_3_willOverflow;
  reg                 handshakeTimes_4_willIncrement;
  reg                 handshakeTimes_4_willClear;
  reg        [12:0]   handshakeTimes_4_valueNext;
  reg        [12:0]   handshakeTimes_4_value;
  wire                handshakeTimes_4_willOverflowIfInc;
  wire                handshakeTimes_4_willOverflow;
  reg                 handshakeTimes_5_willIncrement;
  reg                 handshakeTimes_5_willClear;
  reg        [12:0]   handshakeTimes_5_valueNext;
  reg        [12:0]   handshakeTimes_5_value;
  wire                handshakeTimes_5_willOverflowIfInc;
  wire                handshakeTimes_5_willOverflow;
  reg                 handshakeTimes_6_willIncrement;
  reg                 handshakeTimes_6_willClear;
  reg        [12:0]   handshakeTimes_6_valueNext;
  reg        [12:0]   handshakeTimes_6_value;
  wire                handshakeTimes_6_willOverflowIfInc;
  wire                handshakeTimes_6_willOverflow;
  reg                 handshakeTimes_7_willIncrement;
  reg                 handshakeTimes_7_willClear;
  reg        [12:0]   handshakeTimes_7_valueNext;
  reg        [12:0]   handshakeTimes_7_value;
  wire                handshakeTimes_7_willOverflowIfInc;
  wire                handshakeTimes_7_willOverflow;
  reg        [6:0]    selectWriteFifo;
  reg        [7:0]    selectReadFifo_0;
  reg        [7:0]    selectReadFifo_1;
  reg        [7:0]    selectReadFifo_2;
  reg        [7:0]    selectReadFifo_3;
  reg        [7:0]    selectReadFifo_4;
  reg        [7:0]    selectReadFifo_5;
  reg        [7:0]    selectReadFifo_6;
  reg        [7:0]    selectReadFifo_7;
  reg                 holdReadOp_0;
  reg                 holdReadOp_1;
  reg                 holdReadOp_2;
  reg                 holdReadOp_3;
  reg                 holdReadOp_4;
  reg                 holdReadOp_5;
  reg                 holdReadOp_6;
  reg                 holdReadOp_7;
  reg                 allowPadding_0;
  reg                 allowPadding_1;
  reg                 allowPadding_2;
  reg                 allowPadding_3;
  reg                 allowPadding_4;
  reg                 allowPadding_5;
  reg                 allowPadding_6;
  reg                 allowPadding_7;
  reg                 outSliceNumb_0_willIncrement;
  reg                 outSliceNumb_0_willClear;
  reg        [6:0]    outSliceNumb_0_valueNext;
  reg        [6:0]    outSliceNumb_0_value;
  wire                outSliceNumb_0_willOverflowIfInc;
  wire                outSliceNumb_0_willOverflow;
  reg                 outSliceNumb_1_willIncrement;
  reg                 outSliceNumb_1_willClear;
  reg        [6:0]    outSliceNumb_1_valueNext;
  reg        [6:0]    outSliceNumb_1_value;
  wire                outSliceNumb_1_willOverflowIfInc;
  wire                outSliceNumb_1_willOverflow;
  reg                 outSliceNumb_2_willIncrement;
  reg                 outSliceNumb_2_willClear;
  reg        [6:0]    outSliceNumb_2_valueNext;
  reg        [6:0]    outSliceNumb_2_value;
  wire                outSliceNumb_2_willOverflowIfInc;
  wire                outSliceNumb_2_willOverflow;
  reg                 outSliceNumb_3_willIncrement;
  reg                 outSliceNumb_3_willClear;
  reg        [6:0]    outSliceNumb_3_valueNext;
  reg        [6:0]    outSliceNumb_3_value;
  wire                outSliceNumb_3_willOverflowIfInc;
  wire                outSliceNumb_3_willOverflow;
  reg                 outSliceNumb_4_willIncrement;
  reg                 outSliceNumb_4_willClear;
  reg        [6:0]    outSliceNumb_4_valueNext;
  reg        [6:0]    outSliceNumb_4_value;
  wire                outSliceNumb_4_willOverflowIfInc;
  wire                outSliceNumb_4_willOverflow;
  reg                 outSliceNumb_5_willIncrement;
  reg                 outSliceNumb_5_willClear;
  reg        [6:0]    outSliceNumb_5_valueNext;
  reg        [6:0]    outSliceNumb_5_value;
  wire                outSliceNumb_5_willOverflowIfInc;
  wire                outSliceNumb_5_willOverflow;
  reg                 outSliceNumb_6_willIncrement;
  reg                 outSliceNumb_6_willClear;
  reg        [6:0]    outSliceNumb_6_valueNext;
  reg        [6:0]    outSliceNumb_6_value;
  wire                outSliceNumb_6_willOverflowIfInc;
  wire                outSliceNumb_6_willOverflow;
  reg                 outSliceNumb_7_willIncrement;
  reg                 outSliceNumb_7_willClear;
  reg        [6:0]    outSliceNumb_7_valueNext;
  reg        [6:0]    outSliceNumb_7_value;
  wire                outSliceNumb_7_willOverflowIfInc;
  wire                outSliceNumb_7_willOverflow;
  reg                 writeAround;
  reg                 readAround_0;
  reg                 readAround_1;
  reg                 readAround_2;
  reg                 readAround_3;
  reg                 readAround_4;
  reg                 readAround_5;
  reg                 readAround_6;
  reg                 readAround_7;
  wire                arraySliceStateMachine_wantExit;
  reg                 arraySliceStateMachine_wantStart;
  wire                arraySliceStateMachine_wantKill;
  wire       [1:0]    stateIndicate;
  reg        [1:0]    arraySliceStateMachine_stateReg;
  reg        [1:0]    arraySliceStateMachine_stateNext;
  wire                when_ArraySlice_l204;
  wire                _zz_io_push_valid;
  wire       [31:0]   _zz_io_push_payload;
  wire       [127:0]  _zz_1;
  wire       [127:0]  _zz_2;
  wire                inputStreamArrayData_fire;
  wire                when_ArraySlice_l208;
  wire                when_ArraySlice_l209;
  reg                 debug_0 /* verilator public */ ;
  reg                 debug_1 /* verilator public */ ;
  reg                 debug_2 /* verilator public */ ;
  reg                 debug_3 /* verilator public */ ;
  reg                 debug_4 /* verilator public */ ;
  reg                 debug_5 /* verilator public */ ;
  reg                 debug_6 /* verilator public */ ;
  reg                 debug_7 /* verilator public */ ;
  wire                when_ArraySlice_l158;
  wire                when_ArraySlice_l159;
  reg        [7:0]    realValue_0 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0;
  wire                when_ArraySlice_l110;
  wire                when_ArraySlice_l166;
  wire                when_ArraySlice_l158_1;
  wire                when_ArraySlice_l159_1;
  reg        [7:0]    realValue_0_1 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_1;
  wire                when_ArraySlice_l110_1;
  wire                when_ArraySlice_l166_1;
  wire                when_ArraySlice_l158_2;
  wire                when_ArraySlice_l159_2;
  reg        [7:0]    realValue_0_2 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_2;
  wire                when_ArraySlice_l110_2;
  wire                when_ArraySlice_l166_2;
  wire                when_ArraySlice_l158_3;
  wire                when_ArraySlice_l159_3;
  reg        [7:0]    realValue_0_3 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_3;
  wire                when_ArraySlice_l110_3;
  wire                when_ArraySlice_l166_3;
  wire                when_ArraySlice_l158_4;
  wire                when_ArraySlice_l159_4;
  reg        [7:0]    realValue_0_4 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_4;
  wire                when_ArraySlice_l110_4;
  wire                when_ArraySlice_l166_4;
  wire                when_ArraySlice_l158_5;
  wire                when_ArraySlice_l159_5;
  reg        [7:0]    realValue_0_5 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_5;
  wire                when_ArraySlice_l110_5;
  wire                when_ArraySlice_l166_5;
  wire                when_ArraySlice_l158_6;
  wire                when_ArraySlice_l159_6;
  reg        [7:0]    realValue_0_6 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_6;
  wire                when_ArraySlice_l110_6;
  wire                when_ArraySlice_l166_6;
  wire                when_ArraySlice_l158_7;
  wire                when_ArraySlice_l159_7;
  reg        [7:0]    realValue_0_7 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_7;
  wire                when_ArraySlice_l110_7;
  wire                when_ArraySlice_l166_7;
  wire                when_ArraySlice_l216;
  wire                when_ArraySlice_l222;
  wire                when_ArraySlice_l222_1;
  wire                when_ArraySlice_l222_2;
  wire                when_ArraySlice_l222_3;
  wire                when_ArraySlice_l222_4;
  wire                when_ArraySlice_l222_5;
  wire                when_ArraySlice_l222_6;
  wire                when_ArraySlice_l222_7;
  wire                when_ArraySlice_l376;
  wire                when_ArraySlice_l377;
  wire       [7:0]    _zz_outputStreamArrayData_0_valid;
  wire                _zz_io_pop_ready;
  wire       [127:0]  _zz_3;
  wire                when_ArraySlice_l382;
  wire                outputStreamArrayData_0_fire;
  wire                when_ArraySlice_l383;
  wire                when_ArraySlice_l384;
  wire                when_ArraySlice_l387;
  wire                outputStreamArrayData_0_fire_1;
  wire                when_ArraySlice_l392;
  wire                when_ArraySlice_l393;
  reg        [7:0]    realValue1_0 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0;
  wire                when_ArraySlice_l95;
  wire                when_ArraySlice_l395;
  reg                 debug_0_1 /* verilator public */ ;
  reg                 debug_1_1 /* verilator public */ ;
  reg                 debug_2_1 /* verilator public */ ;
  reg                 debug_3_1 /* verilator public */ ;
  reg                 debug_4_1 /* verilator public */ ;
  reg                 debug_5_1 /* verilator public */ ;
  reg                 debug_6_1 /* verilator public */ ;
  reg                 debug_7_1 /* verilator public */ ;
  wire                when_ArraySlice_l158_8;
  wire                when_ArraySlice_l159_8;
  reg        [7:0]    realValue_0_8 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_8;
  wire                when_ArraySlice_l110_8;
  wire                when_ArraySlice_l166_8;
  wire                when_ArraySlice_l158_9;
  wire                when_ArraySlice_l159_9;
  reg        [7:0]    realValue_0_9 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_9;
  wire                when_ArraySlice_l110_9;
  wire                when_ArraySlice_l166_9;
  wire                when_ArraySlice_l158_10;
  wire                when_ArraySlice_l159_10;
  reg        [7:0]    realValue_0_10 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_10;
  wire                when_ArraySlice_l110_10;
  wire                when_ArraySlice_l166_10;
  wire                when_ArraySlice_l158_11;
  wire                when_ArraySlice_l159_11;
  reg        [7:0]    realValue_0_11 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_11;
  wire                when_ArraySlice_l110_11;
  wire                when_ArraySlice_l166_11;
  wire                when_ArraySlice_l158_12;
  wire                when_ArraySlice_l159_12;
  reg        [7:0]    realValue_0_12 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_12;
  wire                when_ArraySlice_l110_12;
  wire                when_ArraySlice_l166_12;
  wire                when_ArraySlice_l158_13;
  wire                when_ArraySlice_l159_13;
  reg        [7:0]    realValue_0_13 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_13;
  wire                when_ArraySlice_l110_13;
  wire                when_ArraySlice_l166_13;
  wire                when_ArraySlice_l158_14;
  wire                when_ArraySlice_l159_14;
  reg        [7:0]    realValue_0_14 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_14;
  wire                when_ArraySlice_l110_14;
  wire                when_ArraySlice_l166_14;
  wire                when_ArraySlice_l158_15;
  wire                when_ArraySlice_l159_15;
  reg        [7:0]    realValue_0_15 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_15;
  wire                when_ArraySlice_l110_15;
  wire                when_ArraySlice_l166_15;
  wire                when_ArraySlice_l400;
  wire                when_ArraySlice_l403;
  wire                when_ArraySlice_l406;
  wire                when_ArraySlice_l413;
  wire                when_ArraySlice_l417;
  wire                outputStreamArrayData_0_fire_2;
  wire                when_ArraySlice_l418;
  reg        [7:0]    realValue1_0_1 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_1;
  wire                when_ArraySlice_l95_1;
  wire                when_ArraySlice_l420;
  reg                 debug_0_2 /* verilator public */ ;
  reg                 debug_1_2 /* verilator public */ ;
  reg                 debug_2_2 /* verilator public */ ;
  reg                 debug_3_2 /* verilator public */ ;
  reg                 debug_4_2 /* verilator public */ ;
  reg                 debug_5_2 /* verilator public */ ;
  reg                 debug_6_2 /* verilator public */ ;
  reg                 debug_7_2 /* verilator public */ ;
  wire                when_ArraySlice_l158_16;
  wire                when_ArraySlice_l159_16;
  reg        [7:0]    realValue_0_16 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_16;
  wire                when_ArraySlice_l110_16;
  wire                when_ArraySlice_l166_16;
  wire                when_ArraySlice_l158_17;
  wire                when_ArraySlice_l159_17;
  reg        [7:0]    realValue_0_17 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_17;
  wire                when_ArraySlice_l110_17;
  wire                when_ArraySlice_l166_17;
  wire                when_ArraySlice_l158_18;
  wire                when_ArraySlice_l159_18;
  reg        [7:0]    realValue_0_18 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_18;
  wire                when_ArraySlice_l110_18;
  wire                when_ArraySlice_l166_18;
  wire                when_ArraySlice_l158_19;
  wire                when_ArraySlice_l159_19;
  reg        [7:0]    realValue_0_19 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_19;
  wire                when_ArraySlice_l110_19;
  wire                when_ArraySlice_l166_19;
  wire                when_ArraySlice_l158_20;
  wire                when_ArraySlice_l159_20;
  reg        [7:0]    realValue_0_20 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_20;
  wire                when_ArraySlice_l110_20;
  wire                when_ArraySlice_l166_20;
  wire                when_ArraySlice_l158_21;
  wire                when_ArraySlice_l159_21;
  reg        [7:0]    realValue_0_21 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_21;
  wire                when_ArraySlice_l110_21;
  wire                when_ArraySlice_l166_21;
  wire                when_ArraySlice_l158_22;
  wire                when_ArraySlice_l159_22;
  reg        [7:0]    realValue_0_22 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_22;
  wire                when_ArraySlice_l110_22;
  wire                when_ArraySlice_l166_22;
  wire                when_ArraySlice_l158_23;
  wire                when_ArraySlice_l159_23;
  reg        [7:0]    realValue_0_23 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_23;
  wire                when_ArraySlice_l110_23;
  wire                when_ArraySlice_l166_23;
  wire                when_ArraySlice_l425;
  wire                when_ArraySlice_l428;
  wire                when_ArraySlice_l431;
  wire                outputStreamArrayData_0_fire_3;
  wire                when_ArraySlice_l438;
  wire                outputStreamArrayData_0_fire_4;
  wire                when_ArraySlice_l449;
  reg        [7:0]    realValue1_0_2 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_2;
  wire                when_ArraySlice_l95_2;
  wire                when_ArraySlice_l450;
  reg                 debug_0_3 /* verilator public */ ;
  reg                 debug_1_3 /* verilator public */ ;
  reg                 debug_2_3 /* verilator public */ ;
  reg                 debug_3_3 /* verilator public */ ;
  reg                 debug_4_3 /* verilator public */ ;
  reg                 debug_5_3 /* verilator public */ ;
  reg                 debug_6_3 /* verilator public */ ;
  reg                 debug_7_3 /* verilator public */ ;
  wire                when_ArraySlice_l158_24;
  wire                when_ArraySlice_l159_24;
  reg        [7:0]    realValue_0_24 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_24;
  wire                when_ArraySlice_l110_24;
  wire                when_ArraySlice_l166_24;
  wire                when_ArraySlice_l158_25;
  wire                when_ArraySlice_l159_25;
  reg        [7:0]    realValue_0_25 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_25;
  wire                when_ArraySlice_l110_25;
  wire                when_ArraySlice_l166_25;
  wire                when_ArraySlice_l158_26;
  wire                when_ArraySlice_l159_26;
  reg        [7:0]    realValue_0_26 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_26;
  wire                when_ArraySlice_l110_26;
  wire                when_ArraySlice_l166_26;
  wire                when_ArraySlice_l158_27;
  wire                when_ArraySlice_l159_27;
  reg        [7:0]    realValue_0_27 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_27;
  wire                when_ArraySlice_l110_27;
  wire                when_ArraySlice_l166_27;
  wire                when_ArraySlice_l158_28;
  wire                when_ArraySlice_l159_28;
  reg        [7:0]    realValue_0_28 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_28;
  wire                when_ArraySlice_l110_28;
  wire                when_ArraySlice_l166_28;
  wire                when_ArraySlice_l158_29;
  wire                when_ArraySlice_l159_29;
  reg        [7:0]    realValue_0_29 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_29;
  wire                when_ArraySlice_l110_29;
  wire                when_ArraySlice_l166_29;
  wire                when_ArraySlice_l158_30;
  wire                when_ArraySlice_l159_30;
  reg        [7:0]    realValue_0_30 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_30;
  wire                when_ArraySlice_l110_30;
  wire                when_ArraySlice_l166_30;
  wire                when_ArraySlice_l158_31;
  wire                when_ArraySlice_l159_31;
  reg        [7:0]    realValue_0_31 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_31;
  wire                when_ArraySlice_l110_31;
  wire                when_ArraySlice_l166_31;
  wire                when_ArraySlice_l457;
  wire                outputStreamArrayData_0_fire_5;
  wire                when_ArraySlice_l461;
  wire                when_ArraySlice_l447;
  wire                outputStreamArrayData_0_fire_6;
  wire                when_ArraySlice_l468;
  wire                when_ArraySlice_l376_1;
  wire                when_ArraySlice_l377_1;
  wire       [7:0]    _zz_outputStreamArrayData_1_valid;
  wire                _zz_io_pop_ready_1;
  wire       [127:0]  _zz_4;
  wire                when_ArraySlice_l382_1;
  wire                outputStreamArrayData_1_fire;
  wire                when_ArraySlice_l383_1;
  wire                when_ArraySlice_l384_1;
  wire                when_ArraySlice_l387_1;
  wire                outputStreamArrayData_1_fire_1;
  wire                when_ArraySlice_l392_1;
  wire                when_ArraySlice_l393_1;
  reg        [7:0]    realValue1_0_3 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_3;
  wire                when_ArraySlice_l95_3;
  wire                when_ArraySlice_l395_1;
  reg                 debug_0_4 /* verilator public */ ;
  reg                 debug_1_4 /* verilator public */ ;
  reg                 debug_2_4 /* verilator public */ ;
  reg                 debug_3_4 /* verilator public */ ;
  reg                 debug_4_4 /* verilator public */ ;
  reg                 debug_5_4 /* verilator public */ ;
  reg                 debug_6_4 /* verilator public */ ;
  reg                 debug_7_4 /* verilator public */ ;
  wire                when_ArraySlice_l158_32;
  wire                when_ArraySlice_l159_32;
  reg        [7:0]    realValue_0_32 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_32;
  wire                when_ArraySlice_l110_32;
  wire                when_ArraySlice_l166_32;
  wire                when_ArraySlice_l158_33;
  wire                when_ArraySlice_l159_33;
  reg        [7:0]    realValue_0_33 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_33;
  wire                when_ArraySlice_l110_33;
  wire                when_ArraySlice_l166_33;
  wire                when_ArraySlice_l158_34;
  wire                when_ArraySlice_l159_34;
  reg        [7:0]    realValue_0_34 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_34;
  wire                when_ArraySlice_l110_34;
  wire                when_ArraySlice_l166_34;
  wire                when_ArraySlice_l158_35;
  wire                when_ArraySlice_l159_35;
  reg        [7:0]    realValue_0_35 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_35;
  wire                when_ArraySlice_l110_35;
  wire                when_ArraySlice_l166_35;
  wire                when_ArraySlice_l158_36;
  wire                when_ArraySlice_l159_36;
  reg        [7:0]    realValue_0_36 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_36;
  wire                when_ArraySlice_l110_36;
  wire                when_ArraySlice_l166_36;
  wire                when_ArraySlice_l158_37;
  wire                when_ArraySlice_l159_37;
  reg        [7:0]    realValue_0_37 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_37;
  wire                when_ArraySlice_l110_37;
  wire                when_ArraySlice_l166_37;
  wire                when_ArraySlice_l158_38;
  wire                when_ArraySlice_l159_38;
  reg        [7:0]    realValue_0_38 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_38;
  wire                when_ArraySlice_l110_38;
  wire                when_ArraySlice_l166_38;
  wire                when_ArraySlice_l158_39;
  wire                when_ArraySlice_l159_39;
  reg        [7:0]    realValue_0_39 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_39;
  wire                when_ArraySlice_l110_39;
  wire                when_ArraySlice_l166_39;
  wire                when_ArraySlice_l400_1;
  wire                when_ArraySlice_l403_1;
  wire                when_ArraySlice_l406_1;
  wire                when_ArraySlice_l413_1;
  wire                when_ArraySlice_l417_1;
  wire                outputStreamArrayData_1_fire_2;
  wire                when_ArraySlice_l418_1;
  reg        [7:0]    realValue1_0_4 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_4;
  wire                when_ArraySlice_l95_4;
  wire                when_ArraySlice_l420_1;
  reg                 debug_0_5 /* verilator public */ ;
  reg                 debug_1_5 /* verilator public */ ;
  reg                 debug_2_5 /* verilator public */ ;
  reg                 debug_3_5 /* verilator public */ ;
  reg                 debug_4_5 /* verilator public */ ;
  reg                 debug_5_5 /* verilator public */ ;
  reg                 debug_6_5 /* verilator public */ ;
  reg                 debug_7_5 /* verilator public */ ;
  wire                when_ArraySlice_l158_40;
  wire                when_ArraySlice_l159_40;
  reg        [7:0]    realValue_0_40 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_40;
  wire                when_ArraySlice_l110_40;
  wire                when_ArraySlice_l166_40;
  wire                when_ArraySlice_l158_41;
  wire                when_ArraySlice_l159_41;
  reg        [7:0]    realValue_0_41 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_41;
  wire                when_ArraySlice_l110_41;
  wire                when_ArraySlice_l166_41;
  wire                when_ArraySlice_l158_42;
  wire                when_ArraySlice_l159_42;
  reg        [7:0]    realValue_0_42 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_42;
  wire                when_ArraySlice_l110_42;
  wire                when_ArraySlice_l166_42;
  wire                when_ArraySlice_l158_43;
  wire                when_ArraySlice_l159_43;
  reg        [7:0]    realValue_0_43 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_43;
  wire                when_ArraySlice_l110_43;
  wire                when_ArraySlice_l166_43;
  wire                when_ArraySlice_l158_44;
  wire                when_ArraySlice_l159_44;
  reg        [7:0]    realValue_0_44 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_44;
  wire                when_ArraySlice_l110_44;
  wire                when_ArraySlice_l166_44;
  wire                when_ArraySlice_l158_45;
  wire                when_ArraySlice_l159_45;
  reg        [7:0]    realValue_0_45 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_45;
  wire                when_ArraySlice_l110_45;
  wire                when_ArraySlice_l166_45;
  wire                when_ArraySlice_l158_46;
  wire                when_ArraySlice_l159_46;
  reg        [7:0]    realValue_0_46 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_46;
  wire                when_ArraySlice_l110_46;
  wire                when_ArraySlice_l166_46;
  wire                when_ArraySlice_l158_47;
  wire                when_ArraySlice_l159_47;
  reg        [7:0]    realValue_0_47 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_47;
  wire                when_ArraySlice_l110_47;
  wire                when_ArraySlice_l166_47;
  wire                when_ArraySlice_l425_1;
  wire                when_ArraySlice_l428_1;
  wire                when_ArraySlice_l431_1;
  wire                outputStreamArrayData_1_fire_3;
  wire                when_ArraySlice_l438_1;
  wire                outputStreamArrayData_1_fire_4;
  wire                when_ArraySlice_l449_1;
  reg        [7:0]    realValue1_0_5 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_5;
  wire                when_ArraySlice_l95_5;
  wire                when_ArraySlice_l450_1;
  reg                 debug_0_6 /* verilator public */ ;
  reg                 debug_1_6 /* verilator public */ ;
  reg                 debug_2_6 /* verilator public */ ;
  reg                 debug_3_6 /* verilator public */ ;
  reg                 debug_4_6 /* verilator public */ ;
  reg                 debug_5_6 /* verilator public */ ;
  reg                 debug_6_6 /* verilator public */ ;
  reg                 debug_7_6 /* verilator public */ ;
  wire                when_ArraySlice_l158_48;
  wire                when_ArraySlice_l159_48;
  reg        [7:0]    realValue_0_48 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_48;
  wire                when_ArraySlice_l110_48;
  wire                when_ArraySlice_l166_48;
  wire                when_ArraySlice_l158_49;
  wire                when_ArraySlice_l159_49;
  reg        [7:0]    realValue_0_49 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_49;
  wire                when_ArraySlice_l110_49;
  wire                when_ArraySlice_l166_49;
  wire                when_ArraySlice_l158_50;
  wire                when_ArraySlice_l159_50;
  reg        [7:0]    realValue_0_50 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_50;
  wire                when_ArraySlice_l110_50;
  wire                when_ArraySlice_l166_50;
  wire                when_ArraySlice_l158_51;
  wire                when_ArraySlice_l159_51;
  reg        [7:0]    realValue_0_51 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_51;
  wire                when_ArraySlice_l110_51;
  wire                when_ArraySlice_l166_51;
  wire                when_ArraySlice_l158_52;
  wire                when_ArraySlice_l159_52;
  reg        [7:0]    realValue_0_52 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_52;
  wire                when_ArraySlice_l110_52;
  wire                when_ArraySlice_l166_52;
  wire                when_ArraySlice_l158_53;
  wire                when_ArraySlice_l159_53;
  reg        [7:0]    realValue_0_53 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_53;
  wire                when_ArraySlice_l110_53;
  wire                when_ArraySlice_l166_53;
  wire                when_ArraySlice_l158_54;
  wire                when_ArraySlice_l159_54;
  reg        [7:0]    realValue_0_54 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_54;
  wire                when_ArraySlice_l110_54;
  wire                when_ArraySlice_l166_54;
  wire                when_ArraySlice_l158_55;
  wire                when_ArraySlice_l159_55;
  reg        [7:0]    realValue_0_55 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_55;
  wire                when_ArraySlice_l110_55;
  wire                when_ArraySlice_l166_55;
  wire                when_ArraySlice_l457_1;
  wire                outputStreamArrayData_1_fire_5;
  wire                when_ArraySlice_l461_1;
  wire                when_ArraySlice_l447_1;
  wire                outputStreamArrayData_1_fire_6;
  wire                when_ArraySlice_l468_1;
  wire                when_ArraySlice_l376_2;
  wire                when_ArraySlice_l377_2;
  wire       [7:0]    _zz_outputStreamArrayData_2_valid;
  wire                _zz_io_pop_ready_2;
  wire       [127:0]  _zz_5;
  wire                when_ArraySlice_l382_2;
  wire                outputStreamArrayData_2_fire;
  wire                when_ArraySlice_l383_2;
  wire                when_ArraySlice_l384_2;
  wire                when_ArraySlice_l387_2;
  wire                outputStreamArrayData_2_fire_1;
  wire                when_ArraySlice_l392_2;
  wire                when_ArraySlice_l393_2;
  reg        [7:0]    realValue1_0_6 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_6;
  wire                when_ArraySlice_l95_6;
  wire                when_ArraySlice_l395_2;
  reg                 debug_0_7 /* verilator public */ ;
  reg                 debug_1_7 /* verilator public */ ;
  reg                 debug_2_7 /* verilator public */ ;
  reg                 debug_3_7 /* verilator public */ ;
  reg                 debug_4_7 /* verilator public */ ;
  reg                 debug_5_7 /* verilator public */ ;
  reg                 debug_6_7 /* verilator public */ ;
  reg                 debug_7_7 /* verilator public */ ;
  wire                when_ArraySlice_l158_56;
  wire                when_ArraySlice_l159_56;
  reg        [7:0]    realValue_0_56 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_56;
  wire                when_ArraySlice_l110_56;
  wire                when_ArraySlice_l166_56;
  wire                when_ArraySlice_l158_57;
  wire                when_ArraySlice_l159_57;
  reg        [7:0]    realValue_0_57 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_57;
  wire                when_ArraySlice_l110_57;
  wire                when_ArraySlice_l166_57;
  wire                when_ArraySlice_l158_58;
  wire                when_ArraySlice_l159_58;
  reg        [7:0]    realValue_0_58 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_58;
  wire                when_ArraySlice_l110_58;
  wire                when_ArraySlice_l166_58;
  wire                when_ArraySlice_l158_59;
  wire                when_ArraySlice_l159_59;
  reg        [7:0]    realValue_0_59 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_59;
  wire                when_ArraySlice_l110_59;
  wire                when_ArraySlice_l166_59;
  wire                when_ArraySlice_l158_60;
  wire                when_ArraySlice_l159_60;
  reg        [7:0]    realValue_0_60 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_60;
  wire                when_ArraySlice_l110_60;
  wire                when_ArraySlice_l166_60;
  wire                when_ArraySlice_l158_61;
  wire                when_ArraySlice_l159_61;
  reg        [7:0]    realValue_0_61 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_61;
  wire                when_ArraySlice_l110_61;
  wire                when_ArraySlice_l166_61;
  wire                when_ArraySlice_l158_62;
  wire                when_ArraySlice_l159_62;
  reg        [7:0]    realValue_0_62 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_62;
  wire                when_ArraySlice_l110_62;
  wire                when_ArraySlice_l166_62;
  wire                when_ArraySlice_l158_63;
  wire                when_ArraySlice_l159_63;
  reg        [7:0]    realValue_0_63 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_63;
  wire                when_ArraySlice_l110_63;
  wire                when_ArraySlice_l166_63;
  wire                when_ArraySlice_l400_2;
  wire                when_ArraySlice_l403_2;
  wire                when_ArraySlice_l406_2;
  wire                when_ArraySlice_l413_2;
  wire                when_ArraySlice_l417_2;
  wire                outputStreamArrayData_2_fire_2;
  wire                when_ArraySlice_l418_2;
  reg        [7:0]    realValue1_0_7 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_7;
  wire                when_ArraySlice_l95_7;
  wire                when_ArraySlice_l420_2;
  reg                 debug_0_8 /* verilator public */ ;
  reg                 debug_1_8 /* verilator public */ ;
  reg                 debug_2_8 /* verilator public */ ;
  reg                 debug_3_8 /* verilator public */ ;
  reg                 debug_4_8 /* verilator public */ ;
  reg                 debug_5_8 /* verilator public */ ;
  reg                 debug_6_8 /* verilator public */ ;
  reg                 debug_7_8 /* verilator public */ ;
  wire                when_ArraySlice_l158_64;
  wire                when_ArraySlice_l159_64;
  reg        [7:0]    realValue_0_64 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_64;
  wire                when_ArraySlice_l110_64;
  wire                when_ArraySlice_l166_64;
  wire                when_ArraySlice_l158_65;
  wire                when_ArraySlice_l159_65;
  reg        [7:0]    realValue_0_65 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_65;
  wire                when_ArraySlice_l110_65;
  wire                when_ArraySlice_l166_65;
  wire                when_ArraySlice_l158_66;
  wire                when_ArraySlice_l159_66;
  reg        [7:0]    realValue_0_66 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_66;
  wire                when_ArraySlice_l110_66;
  wire                when_ArraySlice_l166_66;
  wire                when_ArraySlice_l158_67;
  wire                when_ArraySlice_l159_67;
  reg        [7:0]    realValue_0_67 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_67;
  wire                when_ArraySlice_l110_67;
  wire                when_ArraySlice_l166_67;
  wire                when_ArraySlice_l158_68;
  wire                when_ArraySlice_l159_68;
  reg        [7:0]    realValue_0_68 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_68;
  wire                when_ArraySlice_l110_68;
  wire                when_ArraySlice_l166_68;
  wire                when_ArraySlice_l158_69;
  wire                when_ArraySlice_l159_69;
  reg        [7:0]    realValue_0_69 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_69;
  wire                when_ArraySlice_l110_69;
  wire                when_ArraySlice_l166_69;
  wire                when_ArraySlice_l158_70;
  wire                when_ArraySlice_l159_70;
  reg        [7:0]    realValue_0_70 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_70;
  wire                when_ArraySlice_l110_70;
  wire                when_ArraySlice_l166_70;
  wire                when_ArraySlice_l158_71;
  wire                when_ArraySlice_l159_71;
  reg        [7:0]    realValue_0_71 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_71;
  wire                when_ArraySlice_l110_71;
  wire                when_ArraySlice_l166_71;
  wire                when_ArraySlice_l425_2;
  wire                when_ArraySlice_l428_2;
  wire                when_ArraySlice_l431_2;
  wire                outputStreamArrayData_2_fire_3;
  wire                when_ArraySlice_l438_2;
  wire                outputStreamArrayData_2_fire_4;
  wire                when_ArraySlice_l449_2;
  reg        [7:0]    realValue1_0_8 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_8;
  wire                when_ArraySlice_l95_8;
  wire                when_ArraySlice_l450_2;
  reg                 debug_0_9 /* verilator public */ ;
  reg                 debug_1_9 /* verilator public */ ;
  reg                 debug_2_9 /* verilator public */ ;
  reg                 debug_3_9 /* verilator public */ ;
  reg                 debug_4_9 /* verilator public */ ;
  reg                 debug_5_9 /* verilator public */ ;
  reg                 debug_6_9 /* verilator public */ ;
  reg                 debug_7_9 /* verilator public */ ;
  wire                when_ArraySlice_l158_72;
  wire                when_ArraySlice_l159_72;
  reg        [7:0]    realValue_0_72 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_72;
  wire                when_ArraySlice_l110_72;
  wire                when_ArraySlice_l166_72;
  wire                when_ArraySlice_l158_73;
  wire                when_ArraySlice_l159_73;
  reg        [7:0]    realValue_0_73 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_73;
  wire                when_ArraySlice_l110_73;
  wire                when_ArraySlice_l166_73;
  wire                when_ArraySlice_l158_74;
  wire                when_ArraySlice_l159_74;
  reg        [7:0]    realValue_0_74 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_74;
  wire                when_ArraySlice_l110_74;
  wire                when_ArraySlice_l166_74;
  wire                when_ArraySlice_l158_75;
  wire                when_ArraySlice_l159_75;
  reg        [7:0]    realValue_0_75 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_75;
  wire                when_ArraySlice_l110_75;
  wire                when_ArraySlice_l166_75;
  wire                when_ArraySlice_l158_76;
  wire                when_ArraySlice_l159_76;
  reg        [7:0]    realValue_0_76 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_76;
  wire                when_ArraySlice_l110_76;
  wire                when_ArraySlice_l166_76;
  wire                when_ArraySlice_l158_77;
  wire                when_ArraySlice_l159_77;
  reg        [7:0]    realValue_0_77 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_77;
  wire                when_ArraySlice_l110_77;
  wire                when_ArraySlice_l166_77;
  wire                when_ArraySlice_l158_78;
  wire                when_ArraySlice_l159_78;
  reg        [7:0]    realValue_0_78 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_78;
  wire                when_ArraySlice_l110_78;
  wire                when_ArraySlice_l166_78;
  wire                when_ArraySlice_l158_79;
  wire                when_ArraySlice_l159_79;
  reg        [7:0]    realValue_0_79 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_79;
  wire                when_ArraySlice_l110_79;
  wire                when_ArraySlice_l166_79;
  wire                when_ArraySlice_l457_2;
  wire                outputStreamArrayData_2_fire_5;
  wire                when_ArraySlice_l461_2;
  wire                when_ArraySlice_l447_2;
  wire                outputStreamArrayData_2_fire_6;
  wire                when_ArraySlice_l468_2;
  wire                when_ArraySlice_l376_3;
  wire                when_ArraySlice_l377_3;
  wire       [7:0]    _zz_outputStreamArrayData_3_valid;
  wire                _zz_io_pop_ready_3;
  wire       [127:0]  _zz_6;
  wire                when_ArraySlice_l382_3;
  wire                outputStreamArrayData_3_fire;
  wire                when_ArraySlice_l383_3;
  wire                when_ArraySlice_l384_3;
  wire                when_ArraySlice_l387_3;
  wire                outputStreamArrayData_3_fire_1;
  wire                when_ArraySlice_l392_3;
  wire                when_ArraySlice_l393_3;
  reg        [7:0]    realValue1_0_9 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_9;
  wire                when_ArraySlice_l95_9;
  wire                when_ArraySlice_l395_3;
  reg                 debug_0_10 /* verilator public */ ;
  reg                 debug_1_10 /* verilator public */ ;
  reg                 debug_2_10 /* verilator public */ ;
  reg                 debug_3_10 /* verilator public */ ;
  reg                 debug_4_10 /* verilator public */ ;
  reg                 debug_5_10 /* verilator public */ ;
  reg                 debug_6_10 /* verilator public */ ;
  reg                 debug_7_10 /* verilator public */ ;
  wire                when_ArraySlice_l158_80;
  wire                when_ArraySlice_l159_80;
  reg        [7:0]    realValue_0_80 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_80;
  wire                when_ArraySlice_l110_80;
  wire                when_ArraySlice_l166_80;
  wire                when_ArraySlice_l158_81;
  wire                when_ArraySlice_l159_81;
  reg        [7:0]    realValue_0_81 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_81;
  wire                when_ArraySlice_l110_81;
  wire                when_ArraySlice_l166_81;
  wire                when_ArraySlice_l158_82;
  wire                when_ArraySlice_l159_82;
  reg        [7:0]    realValue_0_82 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_82;
  wire                when_ArraySlice_l110_82;
  wire                when_ArraySlice_l166_82;
  wire                when_ArraySlice_l158_83;
  wire                when_ArraySlice_l159_83;
  reg        [7:0]    realValue_0_83 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_83;
  wire                when_ArraySlice_l110_83;
  wire                when_ArraySlice_l166_83;
  wire                when_ArraySlice_l158_84;
  wire                when_ArraySlice_l159_84;
  reg        [7:0]    realValue_0_84 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_84;
  wire                when_ArraySlice_l110_84;
  wire                when_ArraySlice_l166_84;
  wire                when_ArraySlice_l158_85;
  wire                when_ArraySlice_l159_85;
  reg        [7:0]    realValue_0_85 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_85;
  wire                when_ArraySlice_l110_85;
  wire                when_ArraySlice_l166_85;
  wire                when_ArraySlice_l158_86;
  wire                when_ArraySlice_l159_86;
  reg        [7:0]    realValue_0_86 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_86;
  wire                when_ArraySlice_l110_86;
  wire                when_ArraySlice_l166_86;
  wire                when_ArraySlice_l158_87;
  wire                when_ArraySlice_l159_87;
  reg        [7:0]    realValue_0_87 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_87;
  wire                when_ArraySlice_l110_87;
  wire                when_ArraySlice_l166_87;
  wire                when_ArraySlice_l400_3;
  wire                when_ArraySlice_l403_3;
  wire                when_ArraySlice_l406_3;
  wire                when_ArraySlice_l413_3;
  wire                when_ArraySlice_l417_3;
  wire                outputStreamArrayData_3_fire_2;
  wire                when_ArraySlice_l418_3;
  reg        [7:0]    realValue1_0_10 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_10;
  wire                when_ArraySlice_l95_10;
  wire                when_ArraySlice_l420_3;
  reg                 debug_0_11 /* verilator public */ ;
  reg                 debug_1_11 /* verilator public */ ;
  reg                 debug_2_11 /* verilator public */ ;
  reg                 debug_3_11 /* verilator public */ ;
  reg                 debug_4_11 /* verilator public */ ;
  reg                 debug_5_11 /* verilator public */ ;
  reg                 debug_6_11 /* verilator public */ ;
  reg                 debug_7_11 /* verilator public */ ;
  wire                when_ArraySlice_l158_88;
  wire                when_ArraySlice_l159_88;
  reg        [7:0]    realValue_0_88 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_88;
  wire                when_ArraySlice_l110_88;
  wire                when_ArraySlice_l166_88;
  wire                when_ArraySlice_l158_89;
  wire                when_ArraySlice_l159_89;
  reg        [7:0]    realValue_0_89 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_89;
  wire                when_ArraySlice_l110_89;
  wire                when_ArraySlice_l166_89;
  wire                when_ArraySlice_l158_90;
  wire                when_ArraySlice_l159_90;
  reg        [7:0]    realValue_0_90 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_90;
  wire                when_ArraySlice_l110_90;
  wire                when_ArraySlice_l166_90;
  wire                when_ArraySlice_l158_91;
  wire                when_ArraySlice_l159_91;
  reg        [7:0]    realValue_0_91 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_91;
  wire                when_ArraySlice_l110_91;
  wire                when_ArraySlice_l166_91;
  wire                when_ArraySlice_l158_92;
  wire                when_ArraySlice_l159_92;
  reg        [7:0]    realValue_0_92 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_92;
  wire                when_ArraySlice_l110_92;
  wire                when_ArraySlice_l166_92;
  wire                when_ArraySlice_l158_93;
  wire                when_ArraySlice_l159_93;
  reg        [7:0]    realValue_0_93 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_93;
  wire                when_ArraySlice_l110_93;
  wire                when_ArraySlice_l166_93;
  wire                when_ArraySlice_l158_94;
  wire                when_ArraySlice_l159_94;
  reg        [7:0]    realValue_0_94 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_94;
  wire                when_ArraySlice_l110_94;
  wire                when_ArraySlice_l166_94;
  wire                when_ArraySlice_l158_95;
  wire                when_ArraySlice_l159_95;
  reg        [7:0]    realValue_0_95 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_95;
  wire                when_ArraySlice_l110_95;
  wire                when_ArraySlice_l166_95;
  wire                when_ArraySlice_l425_3;
  wire                when_ArraySlice_l428_3;
  wire                when_ArraySlice_l431_3;
  wire                outputStreamArrayData_3_fire_3;
  wire                when_ArraySlice_l438_3;
  wire                outputStreamArrayData_3_fire_4;
  wire                when_ArraySlice_l449_3;
  reg        [7:0]    realValue1_0_11 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_11;
  wire                when_ArraySlice_l95_11;
  wire                when_ArraySlice_l450_3;
  reg                 debug_0_12 /* verilator public */ ;
  reg                 debug_1_12 /* verilator public */ ;
  reg                 debug_2_12 /* verilator public */ ;
  reg                 debug_3_12 /* verilator public */ ;
  reg                 debug_4_12 /* verilator public */ ;
  reg                 debug_5_12 /* verilator public */ ;
  reg                 debug_6_12 /* verilator public */ ;
  reg                 debug_7_12 /* verilator public */ ;
  wire                when_ArraySlice_l158_96;
  wire                when_ArraySlice_l159_96;
  reg        [7:0]    realValue_0_96 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_96;
  wire                when_ArraySlice_l110_96;
  wire                when_ArraySlice_l166_96;
  wire                when_ArraySlice_l158_97;
  wire                when_ArraySlice_l159_97;
  reg        [7:0]    realValue_0_97 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_97;
  wire                when_ArraySlice_l110_97;
  wire                when_ArraySlice_l166_97;
  wire                when_ArraySlice_l158_98;
  wire                when_ArraySlice_l159_98;
  reg        [7:0]    realValue_0_98 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_98;
  wire                when_ArraySlice_l110_98;
  wire                when_ArraySlice_l166_98;
  wire                when_ArraySlice_l158_99;
  wire                when_ArraySlice_l159_99;
  reg        [7:0]    realValue_0_99 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_99;
  wire                when_ArraySlice_l110_99;
  wire                when_ArraySlice_l166_99;
  wire                when_ArraySlice_l158_100;
  wire                when_ArraySlice_l159_100;
  reg        [7:0]    realValue_0_100 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_100;
  wire                when_ArraySlice_l110_100;
  wire                when_ArraySlice_l166_100;
  wire                when_ArraySlice_l158_101;
  wire                when_ArraySlice_l159_101;
  reg        [7:0]    realValue_0_101 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_101;
  wire                when_ArraySlice_l110_101;
  wire                when_ArraySlice_l166_101;
  wire                when_ArraySlice_l158_102;
  wire                when_ArraySlice_l159_102;
  reg        [7:0]    realValue_0_102 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_102;
  wire                when_ArraySlice_l110_102;
  wire                when_ArraySlice_l166_102;
  wire                when_ArraySlice_l158_103;
  wire                when_ArraySlice_l159_103;
  reg        [7:0]    realValue_0_103 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_103;
  wire                when_ArraySlice_l110_103;
  wire                when_ArraySlice_l166_103;
  wire                when_ArraySlice_l457_3;
  wire                outputStreamArrayData_3_fire_5;
  wire                when_ArraySlice_l461_3;
  wire                when_ArraySlice_l447_3;
  wire                outputStreamArrayData_3_fire_6;
  wire                when_ArraySlice_l468_3;
  wire                when_ArraySlice_l376_4;
  wire                when_ArraySlice_l377_4;
  wire       [7:0]    _zz_outputStreamArrayData_4_valid;
  wire                _zz_io_pop_ready_4;
  wire       [127:0]  _zz_7;
  wire                when_ArraySlice_l382_4;
  wire                outputStreamArrayData_4_fire;
  wire                when_ArraySlice_l383_4;
  wire                when_ArraySlice_l384_4;
  wire                when_ArraySlice_l387_4;
  wire                outputStreamArrayData_4_fire_1;
  wire                when_ArraySlice_l392_4;
  wire                when_ArraySlice_l393_4;
  reg        [7:0]    realValue1_0_12 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_12;
  wire                when_ArraySlice_l95_12;
  wire                when_ArraySlice_l395_4;
  reg                 debug_0_13 /* verilator public */ ;
  reg                 debug_1_13 /* verilator public */ ;
  reg                 debug_2_13 /* verilator public */ ;
  reg                 debug_3_13 /* verilator public */ ;
  reg                 debug_4_13 /* verilator public */ ;
  reg                 debug_5_13 /* verilator public */ ;
  reg                 debug_6_13 /* verilator public */ ;
  reg                 debug_7_13 /* verilator public */ ;
  wire                when_ArraySlice_l158_104;
  wire                when_ArraySlice_l159_104;
  reg        [7:0]    realValue_0_104 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_104;
  wire                when_ArraySlice_l110_104;
  wire                when_ArraySlice_l166_104;
  wire                when_ArraySlice_l158_105;
  wire                when_ArraySlice_l159_105;
  reg        [7:0]    realValue_0_105 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_105;
  wire                when_ArraySlice_l110_105;
  wire                when_ArraySlice_l166_105;
  wire                when_ArraySlice_l158_106;
  wire                when_ArraySlice_l159_106;
  reg        [7:0]    realValue_0_106 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_106;
  wire                when_ArraySlice_l110_106;
  wire                when_ArraySlice_l166_106;
  wire                when_ArraySlice_l158_107;
  wire                when_ArraySlice_l159_107;
  reg        [7:0]    realValue_0_107 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_107;
  wire                when_ArraySlice_l110_107;
  wire                when_ArraySlice_l166_107;
  wire                when_ArraySlice_l158_108;
  wire                when_ArraySlice_l159_108;
  reg        [7:0]    realValue_0_108 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_108;
  wire                when_ArraySlice_l110_108;
  wire                when_ArraySlice_l166_108;
  wire                when_ArraySlice_l158_109;
  wire                when_ArraySlice_l159_109;
  reg        [7:0]    realValue_0_109 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_109;
  wire                when_ArraySlice_l110_109;
  wire                when_ArraySlice_l166_109;
  wire                when_ArraySlice_l158_110;
  wire                when_ArraySlice_l159_110;
  reg        [7:0]    realValue_0_110 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_110;
  wire                when_ArraySlice_l110_110;
  wire                when_ArraySlice_l166_110;
  wire                when_ArraySlice_l158_111;
  wire                when_ArraySlice_l159_111;
  reg        [7:0]    realValue_0_111 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_111;
  wire                when_ArraySlice_l110_111;
  wire                when_ArraySlice_l166_111;
  wire                when_ArraySlice_l400_4;
  wire                when_ArraySlice_l403_4;
  wire                when_ArraySlice_l406_4;
  wire                when_ArraySlice_l413_4;
  wire                when_ArraySlice_l417_4;
  wire                outputStreamArrayData_4_fire_2;
  wire                when_ArraySlice_l418_4;
  reg        [7:0]    realValue1_0_13 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_13;
  wire                when_ArraySlice_l95_13;
  wire                when_ArraySlice_l420_4;
  reg                 debug_0_14 /* verilator public */ ;
  reg                 debug_1_14 /* verilator public */ ;
  reg                 debug_2_14 /* verilator public */ ;
  reg                 debug_3_14 /* verilator public */ ;
  reg                 debug_4_14 /* verilator public */ ;
  reg                 debug_5_14 /* verilator public */ ;
  reg                 debug_6_14 /* verilator public */ ;
  reg                 debug_7_14 /* verilator public */ ;
  wire                when_ArraySlice_l158_112;
  wire                when_ArraySlice_l159_112;
  reg        [7:0]    realValue_0_112 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_112;
  wire                when_ArraySlice_l110_112;
  wire                when_ArraySlice_l166_112;
  wire                when_ArraySlice_l158_113;
  wire                when_ArraySlice_l159_113;
  reg        [7:0]    realValue_0_113 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_113;
  wire                when_ArraySlice_l110_113;
  wire                when_ArraySlice_l166_113;
  wire                when_ArraySlice_l158_114;
  wire                when_ArraySlice_l159_114;
  reg        [7:0]    realValue_0_114 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_114;
  wire                when_ArraySlice_l110_114;
  wire                when_ArraySlice_l166_114;
  wire                when_ArraySlice_l158_115;
  wire                when_ArraySlice_l159_115;
  reg        [7:0]    realValue_0_115 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_115;
  wire                when_ArraySlice_l110_115;
  wire                when_ArraySlice_l166_115;
  wire                when_ArraySlice_l158_116;
  wire                when_ArraySlice_l159_116;
  reg        [7:0]    realValue_0_116 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_116;
  wire                when_ArraySlice_l110_116;
  wire                when_ArraySlice_l166_116;
  wire                when_ArraySlice_l158_117;
  wire                when_ArraySlice_l159_117;
  reg        [7:0]    realValue_0_117 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_117;
  wire                when_ArraySlice_l110_117;
  wire                when_ArraySlice_l166_117;
  wire                when_ArraySlice_l158_118;
  wire                when_ArraySlice_l159_118;
  reg        [7:0]    realValue_0_118 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_118;
  wire                when_ArraySlice_l110_118;
  wire                when_ArraySlice_l166_118;
  wire                when_ArraySlice_l158_119;
  wire                when_ArraySlice_l159_119;
  reg        [7:0]    realValue_0_119 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_119;
  wire                when_ArraySlice_l110_119;
  wire                when_ArraySlice_l166_119;
  wire                when_ArraySlice_l425_4;
  wire                when_ArraySlice_l428_4;
  wire                when_ArraySlice_l431_4;
  wire                outputStreamArrayData_4_fire_3;
  wire                when_ArraySlice_l438_4;
  wire                outputStreamArrayData_4_fire_4;
  wire                when_ArraySlice_l449_4;
  reg        [7:0]    realValue1_0_14 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_14;
  wire                when_ArraySlice_l95_14;
  wire                when_ArraySlice_l450_4;
  reg                 debug_0_15 /* verilator public */ ;
  reg                 debug_1_15 /* verilator public */ ;
  reg                 debug_2_15 /* verilator public */ ;
  reg                 debug_3_15 /* verilator public */ ;
  reg                 debug_4_15 /* verilator public */ ;
  reg                 debug_5_15 /* verilator public */ ;
  reg                 debug_6_15 /* verilator public */ ;
  reg                 debug_7_15 /* verilator public */ ;
  wire                when_ArraySlice_l158_120;
  wire                when_ArraySlice_l159_120;
  reg        [7:0]    realValue_0_120 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_120;
  wire                when_ArraySlice_l110_120;
  wire                when_ArraySlice_l166_120;
  wire                when_ArraySlice_l158_121;
  wire                when_ArraySlice_l159_121;
  reg        [7:0]    realValue_0_121 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_121;
  wire                when_ArraySlice_l110_121;
  wire                when_ArraySlice_l166_121;
  wire                when_ArraySlice_l158_122;
  wire                when_ArraySlice_l159_122;
  reg        [7:0]    realValue_0_122 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_122;
  wire                when_ArraySlice_l110_122;
  wire                when_ArraySlice_l166_122;
  wire                when_ArraySlice_l158_123;
  wire                when_ArraySlice_l159_123;
  reg        [7:0]    realValue_0_123 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_123;
  wire                when_ArraySlice_l110_123;
  wire                when_ArraySlice_l166_123;
  wire                when_ArraySlice_l158_124;
  wire                when_ArraySlice_l159_124;
  reg        [7:0]    realValue_0_124 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_124;
  wire                when_ArraySlice_l110_124;
  wire                when_ArraySlice_l166_124;
  wire                when_ArraySlice_l158_125;
  wire                when_ArraySlice_l159_125;
  reg        [7:0]    realValue_0_125 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_125;
  wire                when_ArraySlice_l110_125;
  wire                when_ArraySlice_l166_125;
  wire                when_ArraySlice_l158_126;
  wire                when_ArraySlice_l159_126;
  reg        [7:0]    realValue_0_126 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_126;
  wire                when_ArraySlice_l110_126;
  wire                when_ArraySlice_l166_126;
  wire                when_ArraySlice_l158_127;
  wire                when_ArraySlice_l159_127;
  reg        [7:0]    realValue_0_127 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_127;
  wire                when_ArraySlice_l110_127;
  wire                when_ArraySlice_l166_127;
  wire                when_ArraySlice_l457_4;
  wire                outputStreamArrayData_4_fire_5;
  wire                when_ArraySlice_l461_4;
  wire                when_ArraySlice_l447_4;
  wire                outputStreamArrayData_4_fire_6;
  wire                when_ArraySlice_l468_4;
  wire                when_ArraySlice_l376_5;
  wire                when_ArraySlice_l377_5;
  wire       [7:0]    _zz_outputStreamArrayData_5_valid;
  wire                _zz_io_pop_ready_5;
  wire       [127:0]  _zz_8;
  wire                when_ArraySlice_l382_5;
  wire                outputStreamArrayData_5_fire;
  wire                when_ArraySlice_l383_5;
  wire                when_ArraySlice_l384_5;
  wire                when_ArraySlice_l387_5;
  wire                outputStreamArrayData_5_fire_1;
  wire                when_ArraySlice_l392_5;
  wire                when_ArraySlice_l393_5;
  reg        [7:0]    realValue1_0_15 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_15;
  wire                when_ArraySlice_l95_15;
  wire                when_ArraySlice_l395_5;
  reg                 debug_0_16 /* verilator public */ ;
  reg                 debug_1_16 /* verilator public */ ;
  reg                 debug_2_16 /* verilator public */ ;
  reg                 debug_3_16 /* verilator public */ ;
  reg                 debug_4_16 /* verilator public */ ;
  reg                 debug_5_16 /* verilator public */ ;
  reg                 debug_6_16 /* verilator public */ ;
  reg                 debug_7_16 /* verilator public */ ;
  wire                when_ArraySlice_l158_128;
  wire                when_ArraySlice_l159_128;
  reg        [7:0]    realValue_0_128 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_128;
  wire                when_ArraySlice_l110_128;
  wire                when_ArraySlice_l166_128;
  wire                when_ArraySlice_l158_129;
  wire                when_ArraySlice_l159_129;
  reg        [7:0]    realValue_0_129 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_129;
  wire                when_ArraySlice_l110_129;
  wire                when_ArraySlice_l166_129;
  wire                when_ArraySlice_l158_130;
  wire                when_ArraySlice_l159_130;
  reg        [7:0]    realValue_0_130 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_130;
  wire                when_ArraySlice_l110_130;
  wire                when_ArraySlice_l166_130;
  wire                when_ArraySlice_l158_131;
  wire                when_ArraySlice_l159_131;
  reg        [7:0]    realValue_0_131 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_131;
  wire                when_ArraySlice_l110_131;
  wire                when_ArraySlice_l166_131;
  wire                when_ArraySlice_l158_132;
  wire                when_ArraySlice_l159_132;
  reg        [7:0]    realValue_0_132 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_132;
  wire                when_ArraySlice_l110_132;
  wire                when_ArraySlice_l166_132;
  wire                when_ArraySlice_l158_133;
  wire                when_ArraySlice_l159_133;
  reg        [7:0]    realValue_0_133 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_133;
  wire                when_ArraySlice_l110_133;
  wire                when_ArraySlice_l166_133;
  wire                when_ArraySlice_l158_134;
  wire                when_ArraySlice_l159_134;
  reg        [7:0]    realValue_0_134 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_134;
  wire                when_ArraySlice_l110_134;
  wire                when_ArraySlice_l166_134;
  wire                when_ArraySlice_l158_135;
  wire                when_ArraySlice_l159_135;
  reg        [7:0]    realValue_0_135 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_135;
  wire                when_ArraySlice_l110_135;
  wire                when_ArraySlice_l166_135;
  wire                when_ArraySlice_l400_5;
  wire                when_ArraySlice_l403_5;
  wire                when_ArraySlice_l406_5;
  wire                when_ArraySlice_l413_5;
  wire                when_ArraySlice_l417_5;
  wire                outputStreamArrayData_5_fire_2;
  wire                when_ArraySlice_l418_5;
  reg        [7:0]    realValue1_0_16 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_16;
  wire                when_ArraySlice_l95_16;
  wire                when_ArraySlice_l420_5;
  reg                 debug_0_17 /* verilator public */ ;
  reg                 debug_1_17 /* verilator public */ ;
  reg                 debug_2_17 /* verilator public */ ;
  reg                 debug_3_17 /* verilator public */ ;
  reg                 debug_4_17 /* verilator public */ ;
  reg                 debug_5_17 /* verilator public */ ;
  reg                 debug_6_17 /* verilator public */ ;
  reg                 debug_7_17 /* verilator public */ ;
  wire                when_ArraySlice_l158_136;
  wire                when_ArraySlice_l159_136;
  reg        [7:0]    realValue_0_136 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_136;
  wire                when_ArraySlice_l110_136;
  wire                when_ArraySlice_l166_136;
  wire                when_ArraySlice_l158_137;
  wire                when_ArraySlice_l159_137;
  reg        [7:0]    realValue_0_137 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_137;
  wire                when_ArraySlice_l110_137;
  wire                when_ArraySlice_l166_137;
  wire                when_ArraySlice_l158_138;
  wire                when_ArraySlice_l159_138;
  reg        [7:0]    realValue_0_138 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_138;
  wire                when_ArraySlice_l110_138;
  wire                when_ArraySlice_l166_138;
  wire                when_ArraySlice_l158_139;
  wire                when_ArraySlice_l159_139;
  reg        [7:0]    realValue_0_139 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_139;
  wire                when_ArraySlice_l110_139;
  wire                when_ArraySlice_l166_139;
  wire                when_ArraySlice_l158_140;
  wire                when_ArraySlice_l159_140;
  reg        [7:0]    realValue_0_140 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_140;
  wire                when_ArraySlice_l110_140;
  wire                when_ArraySlice_l166_140;
  wire                when_ArraySlice_l158_141;
  wire                when_ArraySlice_l159_141;
  reg        [7:0]    realValue_0_141 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_141;
  wire                when_ArraySlice_l110_141;
  wire                when_ArraySlice_l166_141;
  wire                when_ArraySlice_l158_142;
  wire                when_ArraySlice_l159_142;
  reg        [7:0]    realValue_0_142 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_142;
  wire                when_ArraySlice_l110_142;
  wire                when_ArraySlice_l166_142;
  wire                when_ArraySlice_l158_143;
  wire                when_ArraySlice_l159_143;
  reg        [7:0]    realValue_0_143 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_143;
  wire                when_ArraySlice_l110_143;
  wire                when_ArraySlice_l166_143;
  wire                when_ArraySlice_l425_5;
  wire                when_ArraySlice_l428_5;
  wire                when_ArraySlice_l431_5;
  wire                outputStreamArrayData_5_fire_3;
  wire                when_ArraySlice_l438_5;
  wire                outputStreamArrayData_5_fire_4;
  wire                when_ArraySlice_l449_5;
  reg        [7:0]    realValue1_0_17 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_17;
  wire                when_ArraySlice_l95_17;
  wire                when_ArraySlice_l450_5;
  reg                 debug_0_18 /* verilator public */ ;
  reg                 debug_1_18 /* verilator public */ ;
  reg                 debug_2_18 /* verilator public */ ;
  reg                 debug_3_18 /* verilator public */ ;
  reg                 debug_4_18 /* verilator public */ ;
  reg                 debug_5_18 /* verilator public */ ;
  reg                 debug_6_18 /* verilator public */ ;
  reg                 debug_7_18 /* verilator public */ ;
  wire                when_ArraySlice_l158_144;
  wire                when_ArraySlice_l159_144;
  reg        [7:0]    realValue_0_144 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_144;
  wire                when_ArraySlice_l110_144;
  wire                when_ArraySlice_l166_144;
  wire                when_ArraySlice_l158_145;
  wire                when_ArraySlice_l159_145;
  reg        [7:0]    realValue_0_145 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_145;
  wire                when_ArraySlice_l110_145;
  wire                when_ArraySlice_l166_145;
  wire                when_ArraySlice_l158_146;
  wire                when_ArraySlice_l159_146;
  reg        [7:0]    realValue_0_146 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_146;
  wire                when_ArraySlice_l110_146;
  wire                when_ArraySlice_l166_146;
  wire                when_ArraySlice_l158_147;
  wire                when_ArraySlice_l159_147;
  reg        [7:0]    realValue_0_147 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_147;
  wire                when_ArraySlice_l110_147;
  wire                when_ArraySlice_l166_147;
  wire                when_ArraySlice_l158_148;
  wire                when_ArraySlice_l159_148;
  reg        [7:0]    realValue_0_148 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_148;
  wire                when_ArraySlice_l110_148;
  wire                when_ArraySlice_l166_148;
  wire                when_ArraySlice_l158_149;
  wire                when_ArraySlice_l159_149;
  reg        [7:0]    realValue_0_149 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_149;
  wire                when_ArraySlice_l110_149;
  wire                when_ArraySlice_l166_149;
  wire                when_ArraySlice_l158_150;
  wire                when_ArraySlice_l159_150;
  reg        [7:0]    realValue_0_150 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_150;
  wire                when_ArraySlice_l110_150;
  wire                when_ArraySlice_l166_150;
  wire                when_ArraySlice_l158_151;
  wire                when_ArraySlice_l159_151;
  reg        [7:0]    realValue_0_151 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_151;
  wire                when_ArraySlice_l110_151;
  wire                when_ArraySlice_l166_151;
  wire                when_ArraySlice_l457_5;
  wire                outputStreamArrayData_5_fire_5;
  wire                when_ArraySlice_l461_5;
  wire                when_ArraySlice_l447_5;
  wire                outputStreamArrayData_5_fire_6;
  wire                when_ArraySlice_l468_5;
  wire                when_ArraySlice_l376_6;
  wire                when_ArraySlice_l377_6;
  wire       [7:0]    _zz_outputStreamArrayData_6_valid;
  wire                _zz_io_pop_ready_6;
  wire       [127:0]  _zz_9;
  wire                when_ArraySlice_l382_6;
  wire                outputStreamArrayData_6_fire;
  wire                when_ArraySlice_l383_6;
  wire                when_ArraySlice_l384_6;
  wire                when_ArraySlice_l387_6;
  wire                outputStreamArrayData_6_fire_1;
  wire                when_ArraySlice_l392_6;
  wire                when_ArraySlice_l393_6;
  reg        [7:0]    realValue1_0_18 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_18;
  wire                when_ArraySlice_l95_18;
  wire                when_ArraySlice_l395_6;
  reg                 debug_0_19 /* verilator public */ ;
  reg                 debug_1_19 /* verilator public */ ;
  reg                 debug_2_19 /* verilator public */ ;
  reg                 debug_3_19 /* verilator public */ ;
  reg                 debug_4_19 /* verilator public */ ;
  reg                 debug_5_19 /* verilator public */ ;
  reg                 debug_6_19 /* verilator public */ ;
  reg                 debug_7_19 /* verilator public */ ;
  wire                when_ArraySlice_l158_152;
  wire                when_ArraySlice_l159_152;
  reg        [7:0]    realValue_0_152 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_152;
  wire                when_ArraySlice_l110_152;
  wire                when_ArraySlice_l166_152;
  wire                when_ArraySlice_l158_153;
  wire                when_ArraySlice_l159_153;
  reg        [7:0]    realValue_0_153 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_153;
  wire                when_ArraySlice_l110_153;
  wire                when_ArraySlice_l166_153;
  wire                when_ArraySlice_l158_154;
  wire                when_ArraySlice_l159_154;
  reg        [7:0]    realValue_0_154 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_154;
  wire                when_ArraySlice_l110_154;
  wire                when_ArraySlice_l166_154;
  wire                when_ArraySlice_l158_155;
  wire                when_ArraySlice_l159_155;
  reg        [7:0]    realValue_0_155 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_155;
  wire                when_ArraySlice_l110_155;
  wire                when_ArraySlice_l166_155;
  wire                when_ArraySlice_l158_156;
  wire                when_ArraySlice_l159_156;
  reg        [7:0]    realValue_0_156 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_156;
  wire                when_ArraySlice_l110_156;
  wire                when_ArraySlice_l166_156;
  wire                when_ArraySlice_l158_157;
  wire                when_ArraySlice_l159_157;
  reg        [7:0]    realValue_0_157 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_157;
  wire                when_ArraySlice_l110_157;
  wire                when_ArraySlice_l166_157;
  wire                when_ArraySlice_l158_158;
  wire                when_ArraySlice_l159_158;
  reg        [7:0]    realValue_0_158 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_158;
  wire                when_ArraySlice_l110_158;
  wire                when_ArraySlice_l166_158;
  wire                when_ArraySlice_l158_159;
  wire                when_ArraySlice_l159_159;
  reg        [7:0]    realValue_0_159 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_159;
  wire                when_ArraySlice_l110_159;
  wire                when_ArraySlice_l166_159;
  wire                when_ArraySlice_l400_6;
  wire                when_ArraySlice_l403_6;
  wire                when_ArraySlice_l406_6;
  wire                when_ArraySlice_l413_6;
  wire                when_ArraySlice_l417_6;
  wire                outputStreamArrayData_6_fire_2;
  wire                when_ArraySlice_l418_6;
  reg        [7:0]    realValue1_0_19 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_19;
  wire                when_ArraySlice_l95_19;
  wire                when_ArraySlice_l420_6;
  reg                 debug_0_20 /* verilator public */ ;
  reg                 debug_1_20 /* verilator public */ ;
  reg                 debug_2_20 /* verilator public */ ;
  reg                 debug_3_20 /* verilator public */ ;
  reg                 debug_4_20 /* verilator public */ ;
  reg                 debug_5_20 /* verilator public */ ;
  reg                 debug_6_20 /* verilator public */ ;
  reg                 debug_7_20 /* verilator public */ ;
  wire                when_ArraySlice_l158_160;
  wire                when_ArraySlice_l159_160;
  reg        [7:0]    realValue_0_160 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_160;
  wire                when_ArraySlice_l110_160;
  wire                when_ArraySlice_l166_160;
  wire                when_ArraySlice_l158_161;
  wire                when_ArraySlice_l159_161;
  reg        [7:0]    realValue_0_161 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_161;
  wire                when_ArraySlice_l110_161;
  wire                when_ArraySlice_l166_161;
  wire                when_ArraySlice_l158_162;
  wire                when_ArraySlice_l159_162;
  reg        [7:0]    realValue_0_162 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_162;
  wire                when_ArraySlice_l110_162;
  wire                when_ArraySlice_l166_162;
  wire                when_ArraySlice_l158_163;
  wire                when_ArraySlice_l159_163;
  reg        [7:0]    realValue_0_163 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_163;
  wire                when_ArraySlice_l110_163;
  wire                when_ArraySlice_l166_163;
  wire                when_ArraySlice_l158_164;
  wire                when_ArraySlice_l159_164;
  reg        [7:0]    realValue_0_164 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_164;
  wire                when_ArraySlice_l110_164;
  wire                when_ArraySlice_l166_164;
  wire                when_ArraySlice_l158_165;
  wire                when_ArraySlice_l159_165;
  reg        [7:0]    realValue_0_165 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_165;
  wire                when_ArraySlice_l110_165;
  wire                when_ArraySlice_l166_165;
  wire                when_ArraySlice_l158_166;
  wire                when_ArraySlice_l159_166;
  reg        [7:0]    realValue_0_166 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_166;
  wire                when_ArraySlice_l110_166;
  wire                when_ArraySlice_l166_166;
  wire                when_ArraySlice_l158_167;
  wire                when_ArraySlice_l159_167;
  reg        [7:0]    realValue_0_167 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_167;
  wire                when_ArraySlice_l110_167;
  wire                when_ArraySlice_l166_167;
  wire                when_ArraySlice_l425_6;
  wire                when_ArraySlice_l428_6;
  wire                when_ArraySlice_l431_6;
  wire                outputStreamArrayData_6_fire_3;
  wire                when_ArraySlice_l438_6;
  wire                outputStreamArrayData_6_fire_4;
  wire                when_ArraySlice_l449_6;
  reg        [7:0]    realValue1_0_20 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_20;
  wire                when_ArraySlice_l95_20;
  wire                when_ArraySlice_l450_6;
  reg                 debug_0_21 /* verilator public */ ;
  reg                 debug_1_21 /* verilator public */ ;
  reg                 debug_2_21 /* verilator public */ ;
  reg                 debug_3_21 /* verilator public */ ;
  reg                 debug_4_21 /* verilator public */ ;
  reg                 debug_5_21 /* verilator public */ ;
  reg                 debug_6_21 /* verilator public */ ;
  reg                 debug_7_21 /* verilator public */ ;
  wire                when_ArraySlice_l158_168;
  wire                when_ArraySlice_l159_168;
  reg        [7:0]    realValue_0_168 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_168;
  wire                when_ArraySlice_l110_168;
  wire                when_ArraySlice_l166_168;
  wire                when_ArraySlice_l158_169;
  wire                when_ArraySlice_l159_169;
  reg        [7:0]    realValue_0_169 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_169;
  wire                when_ArraySlice_l110_169;
  wire                when_ArraySlice_l166_169;
  wire                when_ArraySlice_l158_170;
  wire                when_ArraySlice_l159_170;
  reg        [7:0]    realValue_0_170 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_170;
  wire                when_ArraySlice_l110_170;
  wire                when_ArraySlice_l166_170;
  wire                when_ArraySlice_l158_171;
  wire                when_ArraySlice_l159_171;
  reg        [7:0]    realValue_0_171 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_171;
  wire                when_ArraySlice_l110_171;
  wire                when_ArraySlice_l166_171;
  wire                when_ArraySlice_l158_172;
  wire                when_ArraySlice_l159_172;
  reg        [7:0]    realValue_0_172 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_172;
  wire                when_ArraySlice_l110_172;
  wire                when_ArraySlice_l166_172;
  wire                when_ArraySlice_l158_173;
  wire                when_ArraySlice_l159_173;
  reg        [7:0]    realValue_0_173 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_173;
  wire                when_ArraySlice_l110_173;
  wire                when_ArraySlice_l166_173;
  wire                when_ArraySlice_l158_174;
  wire                when_ArraySlice_l159_174;
  reg        [7:0]    realValue_0_174 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_174;
  wire                when_ArraySlice_l110_174;
  wire                when_ArraySlice_l166_174;
  wire                when_ArraySlice_l158_175;
  wire                when_ArraySlice_l159_175;
  reg        [7:0]    realValue_0_175 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_175;
  wire                when_ArraySlice_l110_175;
  wire                when_ArraySlice_l166_175;
  wire                when_ArraySlice_l457_6;
  wire                outputStreamArrayData_6_fire_5;
  wire                when_ArraySlice_l461_6;
  wire                when_ArraySlice_l447_6;
  wire                outputStreamArrayData_6_fire_6;
  wire                when_ArraySlice_l468_6;
  wire                when_ArraySlice_l376_7;
  wire                when_ArraySlice_l377_7;
  wire       [7:0]    _zz_outputStreamArrayData_7_valid;
  wire                _zz_io_pop_ready_7;
  wire       [127:0]  _zz_10;
  wire                when_ArraySlice_l382_7;
  wire                outputStreamArrayData_7_fire;
  wire                when_ArraySlice_l383_7;
  wire                when_ArraySlice_l384_7;
  wire                when_ArraySlice_l387_7;
  wire                outputStreamArrayData_7_fire_1;
  wire                when_ArraySlice_l392_7;
  wire                when_ArraySlice_l393_7;
  reg        [7:0]    realValue1_0_21 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_21;
  wire                when_ArraySlice_l95_21;
  wire                when_ArraySlice_l395_7;
  reg                 debug_0_22 /* verilator public */ ;
  reg                 debug_1_22 /* verilator public */ ;
  reg                 debug_2_22 /* verilator public */ ;
  reg                 debug_3_22 /* verilator public */ ;
  reg                 debug_4_22 /* verilator public */ ;
  reg                 debug_5_22 /* verilator public */ ;
  reg                 debug_6_22 /* verilator public */ ;
  reg                 debug_7_22 /* verilator public */ ;
  wire                when_ArraySlice_l158_176;
  wire                when_ArraySlice_l159_176;
  reg        [7:0]    realValue_0_176 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_176;
  wire                when_ArraySlice_l110_176;
  wire                when_ArraySlice_l166_176;
  wire                when_ArraySlice_l158_177;
  wire                when_ArraySlice_l159_177;
  reg        [7:0]    realValue_0_177 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_177;
  wire                when_ArraySlice_l110_177;
  wire                when_ArraySlice_l166_177;
  wire                when_ArraySlice_l158_178;
  wire                when_ArraySlice_l159_178;
  reg        [7:0]    realValue_0_178 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_178;
  wire                when_ArraySlice_l110_178;
  wire                when_ArraySlice_l166_178;
  wire                when_ArraySlice_l158_179;
  wire                when_ArraySlice_l159_179;
  reg        [7:0]    realValue_0_179 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_179;
  wire                when_ArraySlice_l110_179;
  wire                when_ArraySlice_l166_179;
  wire                when_ArraySlice_l158_180;
  wire                when_ArraySlice_l159_180;
  reg        [7:0]    realValue_0_180 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_180;
  wire                when_ArraySlice_l110_180;
  wire                when_ArraySlice_l166_180;
  wire                when_ArraySlice_l158_181;
  wire                when_ArraySlice_l159_181;
  reg        [7:0]    realValue_0_181 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_181;
  wire                when_ArraySlice_l110_181;
  wire                when_ArraySlice_l166_181;
  wire                when_ArraySlice_l158_182;
  wire                when_ArraySlice_l159_182;
  reg        [7:0]    realValue_0_182 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_182;
  wire                when_ArraySlice_l110_182;
  wire                when_ArraySlice_l166_182;
  wire                when_ArraySlice_l158_183;
  wire                when_ArraySlice_l159_183;
  reg        [7:0]    realValue_0_183 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_183;
  wire                when_ArraySlice_l110_183;
  wire                when_ArraySlice_l166_183;
  wire                when_ArraySlice_l400_7;
  wire                when_ArraySlice_l403_7;
  wire                when_ArraySlice_l406_7;
  wire                when_ArraySlice_l413_7;
  wire                when_ArraySlice_l417_7;
  wire                outputStreamArrayData_7_fire_2;
  wire                when_ArraySlice_l418_7;
  reg        [7:0]    realValue1_0_22 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_22;
  wire                when_ArraySlice_l95_22;
  wire                when_ArraySlice_l420_7;
  reg                 debug_0_23 /* verilator public */ ;
  reg                 debug_1_23 /* verilator public */ ;
  reg                 debug_2_23 /* verilator public */ ;
  reg                 debug_3_23 /* verilator public */ ;
  reg                 debug_4_23 /* verilator public */ ;
  reg                 debug_5_23 /* verilator public */ ;
  reg                 debug_6_23 /* verilator public */ ;
  reg                 debug_7_23 /* verilator public */ ;
  wire                when_ArraySlice_l158_184;
  wire                when_ArraySlice_l159_184;
  reg        [7:0]    realValue_0_184 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_184;
  wire                when_ArraySlice_l110_184;
  wire                when_ArraySlice_l166_184;
  wire                when_ArraySlice_l158_185;
  wire                when_ArraySlice_l159_185;
  reg        [7:0]    realValue_0_185 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_185;
  wire                when_ArraySlice_l110_185;
  wire                when_ArraySlice_l166_185;
  wire                when_ArraySlice_l158_186;
  wire                when_ArraySlice_l159_186;
  reg        [7:0]    realValue_0_186 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_186;
  wire                when_ArraySlice_l110_186;
  wire                when_ArraySlice_l166_186;
  wire                when_ArraySlice_l158_187;
  wire                when_ArraySlice_l159_187;
  reg        [7:0]    realValue_0_187 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_187;
  wire                when_ArraySlice_l110_187;
  wire                when_ArraySlice_l166_187;
  wire                when_ArraySlice_l158_188;
  wire                when_ArraySlice_l159_188;
  reg        [7:0]    realValue_0_188 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_188;
  wire                when_ArraySlice_l110_188;
  wire                when_ArraySlice_l166_188;
  wire                when_ArraySlice_l158_189;
  wire                when_ArraySlice_l159_189;
  reg        [7:0]    realValue_0_189 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_189;
  wire                when_ArraySlice_l110_189;
  wire                when_ArraySlice_l166_189;
  wire                when_ArraySlice_l158_190;
  wire                when_ArraySlice_l159_190;
  reg        [7:0]    realValue_0_190 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_190;
  wire                when_ArraySlice_l110_190;
  wire                when_ArraySlice_l166_190;
  wire                when_ArraySlice_l158_191;
  wire                when_ArraySlice_l159_191;
  reg        [7:0]    realValue_0_191 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_191;
  wire                when_ArraySlice_l110_191;
  wire                when_ArraySlice_l166_191;
  wire                when_ArraySlice_l425_7;
  wire                when_ArraySlice_l428_7;
  wire                when_ArraySlice_l431_7;
  wire                outputStreamArrayData_7_fire_3;
  wire                when_ArraySlice_l438_7;
  wire                outputStreamArrayData_7_fire_4;
  wire                when_ArraySlice_l449_7;
  reg        [7:0]    realValue1_0_23 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_23;
  wire                when_ArraySlice_l95_23;
  wire                when_ArraySlice_l450_7;
  reg                 debug_0_24 /* verilator public */ ;
  reg                 debug_1_24 /* verilator public */ ;
  reg                 debug_2_24 /* verilator public */ ;
  reg                 debug_3_24 /* verilator public */ ;
  reg                 debug_4_24 /* verilator public */ ;
  reg                 debug_5_24 /* verilator public */ ;
  reg                 debug_6_24 /* verilator public */ ;
  reg                 debug_7_24 /* verilator public */ ;
  wire                when_ArraySlice_l158_192;
  wire                when_ArraySlice_l159_192;
  reg        [7:0]    realValue_0_192 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_192;
  wire                when_ArraySlice_l110_192;
  wire                when_ArraySlice_l166_192;
  wire                when_ArraySlice_l158_193;
  wire                when_ArraySlice_l159_193;
  reg        [7:0]    realValue_0_193 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_193;
  wire                when_ArraySlice_l110_193;
  wire                when_ArraySlice_l166_193;
  wire                when_ArraySlice_l158_194;
  wire                when_ArraySlice_l159_194;
  reg        [7:0]    realValue_0_194 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_194;
  wire                when_ArraySlice_l110_194;
  wire                when_ArraySlice_l166_194;
  wire                when_ArraySlice_l158_195;
  wire                when_ArraySlice_l159_195;
  reg        [7:0]    realValue_0_195 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_195;
  wire                when_ArraySlice_l110_195;
  wire                when_ArraySlice_l166_195;
  wire                when_ArraySlice_l158_196;
  wire                when_ArraySlice_l159_196;
  reg        [7:0]    realValue_0_196 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_196;
  wire                when_ArraySlice_l110_196;
  wire                when_ArraySlice_l166_196;
  wire                when_ArraySlice_l158_197;
  wire                when_ArraySlice_l159_197;
  reg        [7:0]    realValue_0_197 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_197;
  wire                when_ArraySlice_l110_197;
  wire                when_ArraySlice_l166_197;
  wire                when_ArraySlice_l158_198;
  wire                when_ArraySlice_l159_198;
  reg        [7:0]    realValue_0_198 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_198;
  wire                when_ArraySlice_l110_198;
  wire                when_ArraySlice_l166_198;
  wire                when_ArraySlice_l158_199;
  wire                when_ArraySlice_l159_199;
  reg        [7:0]    realValue_0_199 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_199;
  wire                when_ArraySlice_l110_199;
  wire                when_ArraySlice_l166_199;
  wire                when_ArraySlice_l457_7;
  wire                outputStreamArrayData_7_fire_5;
  wire                when_ArraySlice_l461_7;
  wire                when_ArraySlice_l447_7;
  wire                outputStreamArrayData_7_fire_6;
  wire                when_ArraySlice_l468_7;
  reg                 debug_0_25 /* verilator public */ ;
  reg                 debug_1_25 /* verilator public */ ;
  reg                 debug_2_25 /* verilator public */ ;
  reg                 debug_3_25 /* verilator public */ ;
  reg                 debug_4_25 /* verilator public */ ;
  reg                 debug_5_25 /* verilator public */ ;
  reg                 debug_6_25 /* verilator public */ ;
  reg                 debug_7_25 /* verilator public */ ;
  wire                when_ArraySlice_l158_200;
  wire                when_ArraySlice_l159_200;
  reg        [7:0]    realValue_0_200 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_200;
  wire                when_ArraySlice_l110_200;
  wire                when_ArraySlice_l166_200;
  wire                when_ArraySlice_l158_201;
  wire                when_ArraySlice_l159_201;
  reg        [7:0]    realValue_0_201 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_201;
  wire                when_ArraySlice_l110_201;
  wire                when_ArraySlice_l166_201;
  wire                when_ArraySlice_l158_202;
  wire                when_ArraySlice_l159_202;
  reg        [7:0]    realValue_0_202 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_202;
  wire                when_ArraySlice_l110_202;
  wire                when_ArraySlice_l166_202;
  wire                when_ArraySlice_l158_203;
  wire                when_ArraySlice_l159_203;
  reg        [7:0]    realValue_0_203 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_203;
  wire                when_ArraySlice_l110_203;
  wire                when_ArraySlice_l166_203;
  wire                when_ArraySlice_l158_204;
  wire                when_ArraySlice_l159_204;
  reg        [7:0]    realValue_0_204 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_204;
  wire                when_ArraySlice_l110_204;
  wire                when_ArraySlice_l166_204;
  wire                when_ArraySlice_l158_205;
  wire                when_ArraySlice_l159_205;
  reg        [7:0]    realValue_0_205 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_205;
  wire                when_ArraySlice_l110_205;
  wire                when_ArraySlice_l166_205;
  wire                when_ArraySlice_l158_206;
  wire                when_ArraySlice_l159_206;
  reg        [7:0]    realValue_0_206 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_206;
  wire                when_ArraySlice_l110_206;
  wire                when_ArraySlice_l166_206;
  wire                when_ArraySlice_l158_207;
  wire                when_ArraySlice_l159_207;
  reg        [7:0]    realValue_0_207 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_207;
  wire                when_ArraySlice_l110_207;
  wire                when_ArraySlice_l166_207;
  wire                when_ArraySlice_l478;
  wire                when_ArraySlice_l481;
  wire                when_ArraySlice_l481_1;
  wire                when_ArraySlice_l481_2;
  wire                when_ArraySlice_l481_3;
  wire                when_ArraySlice_l481_4;
  wire                when_ArraySlice_l481_5;
  wire                when_ArraySlice_l481_6;
  wire                when_ArraySlice_l481_7;
  wire                when_ArraySlice_l233;
  wire                when_ArraySlice_l234;
  wire       [7:0]    _zz_outputStreamArrayData_0_valid_1;
  wire                _zz_io_pop_ready_8;
  wire       [127:0]  _zz_11;
  wire                when_ArraySlice_l239;
  wire                outputStreamArrayData_0_fire_7;
  wire                when_ArraySlice_l240;
  wire                when_ArraySlice_l241;
  wire                when_ArraySlice_l244;
  wire                outputStreamArrayData_0_fire_8;
  wire                when_ArraySlice_l249;
  wire                when_ArraySlice_l250;
  reg        [7:0]    realValue1_0_24 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_24;
  wire                when_ArraySlice_l95_24;
  wire                when_ArraySlice_l252;
  reg                 debug_0_26 /* verilator public */ ;
  reg                 debug_1_26 /* verilator public */ ;
  reg                 debug_2_26 /* verilator public */ ;
  reg                 debug_3_26 /* verilator public */ ;
  reg                 debug_4_26 /* verilator public */ ;
  reg                 debug_5_26 /* verilator public */ ;
  reg                 debug_6_26 /* verilator public */ ;
  reg                 debug_7_26 /* verilator public */ ;
  wire                when_ArraySlice_l158_208;
  wire                when_ArraySlice_l159_208;
  reg        [7:0]    realValue_0_208 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_208;
  wire                when_ArraySlice_l110_208;
  wire                when_ArraySlice_l166_208;
  wire                when_ArraySlice_l158_209;
  wire                when_ArraySlice_l159_209;
  reg        [7:0]    realValue_0_209 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_209;
  wire                when_ArraySlice_l110_209;
  wire                when_ArraySlice_l166_209;
  wire                when_ArraySlice_l158_210;
  wire                when_ArraySlice_l159_210;
  reg        [7:0]    realValue_0_210 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_210;
  wire                when_ArraySlice_l110_210;
  wire                when_ArraySlice_l166_210;
  wire                when_ArraySlice_l158_211;
  wire                when_ArraySlice_l159_211;
  reg        [7:0]    realValue_0_211 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_211;
  wire                when_ArraySlice_l110_211;
  wire                when_ArraySlice_l166_211;
  wire                when_ArraySlice_l158_212;
  wire                when_ArraySlice_l159_212;
  reg        [7:0]    realValue_0_212 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_212;
  wire                when_ArraySlice_l110_212;
  wire                when_ArraySlice_l166_212;
  wire                when_ArraySlice_l158_213;
  wire                when_ArraySlice_l159_213;
  reg        [7:0]    realValue_0_213 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_213;
  wire                when_ArraySlice_l110_213;
  wire                when_ArraySlice_l166_213;
  wire                when_ArraySlice_l158_214;
  wire                when_ArraySlice_l159_214;
  reg        [7:0]    realValue_0_214 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_214;
  wire                when_ArraySlice_l110_214;
  wire                when_ArraySlice_l166_214;
  wire                when_ArraySlice_l158_215;
  wire                when_ArraySlice_l159_215;
  reg        [7:0]    realValue_0_215 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_215;
  wire                when_ArraySlice_l110_215;
  wire                when_ArraySlice_l166_215;
  wire                when_ArraySlice_l257;
  wire                when_ArraySlice_l260;
  wire                when_ArraySlice_l263;
  wire                when_ArraySlice_l270;
  wire                when_ArraySlice_l274;
  wire                outputStreamArrayData_0_fire_9;
  wire                when_ArraySlice_l275;
  reg        [7:0]    realValue1_0_25 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_25;
  wire                when_ArraySlice_l95_25;
  wire                when_ArraySlice_l277;
  reg                 debug_0_27 /* verilator public */ ;
  reg                 debug_1_27 /* verilator public */ ;
  reg                 debug_2_27 /* verilator public */ ;
  reg                 debug_3_27 /* verilator public */ ;
  reg                 debug_4_27 /* verilator public */ ;
  reg                 debug_5_27 /* verilator public */ ;
  reg                 debug_6_27 /* verilator public */ ;
  reg                 debug_7_27 /* verilator public */ ;
  wire                when_ArraySlice_l158_216;
  wire                when_ArraySlice_l159_216;
  reg        [7:0]    realValue_0_216 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_216;
  wire                when_ArraySlice_l110_216;
  wire                when_ArraySlice_l166_216;
  wire                when_ArraySlice_l158_217;
  wire                when_ArraySlice_l159_217;
  reg        [7:0]    realValue_0_217 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_217;
  wire                when_ArraySlice_l110_217;
  wire                when_ArraySlice_l166_217;
  wire                when_ArraySlice_l158_218;
  wire                when_ArraySlice_l159_218;
  reg        [7:0]    realValue_0_218 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_218;
  wire                when_ArraySlice_l110_218;
  wire                when_ArraySlice_l166_218;
  wire                when_ArraySlice_l158_219;
  wire                when_ArraySlice_l159_219;
  reg        [7:0]    realValue_0_219 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_219;
  wire                when_ArraySlice_l110_219;
  wire                when_ArraySlice_l166_219;
  wire                when_ArraySlice_l158_220;
  wire                when_ArraySlice_l159_220;
  reg        [7:0]    realValue_0_220 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_220;
  wire                when_ArraySlice_l110_220;
  wire                when_ArraySlice_l166_220;
  wire                when_ArraySlice_l158_221;
  wire                when_ArraySlice_l159_221;
  reg        [7:0]    realValue_0_221 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_221;
  wire                when_ArraySlice_l110_221;
  wire                when_ArraySlice_l166_221;
  wire                when_ArraySlice_l158_222;
  wire                when_ArraySlice_l159_222;
  reg        [7:0]    realValue_0_222 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_222;
  wire                when_ArraySlice_l110_222;
  wire                when_ArraySlice_l166_222;
  wire                when_ArraySlice_l158_223;
  wire                when_ArraySlice_l159_223;
  reg        [7:0]    realValue_0_223 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_223;
  wire                when_ArraySlice_l110_223;
  wire                when_ArraySlice_l166_223;
  wire                when_ArraySlice_l282;
  wire                when_ArraySlice_l285;
  wire                when_ArraySlice_l288;
  wire                outputStreamArrayData_0_fire_10;
  wire                when_ArraySlice_l295;
  wire                outputStreamArrayData_0_fire_11;
  wire                when_ArraySlice_l306;
  reg        [7:0]    realValue1_0_26 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_26;
  wire                when_ArraySlice_l95_26;
  wire                when_ArraySlice_l307;
  reg                 debug_0_28 /* verilator public */ ;
  reg                 debug_1_28 /* verilator public */ ;
  reg                 debug_2_28 /* verilator public */ ;
  reg                 debug_3_28 /* verilator public */ ;
  reg                 debug_4_28 /* verilator public */ ;
  reg                 debug_5_28 /* verilator public */ ;
  reg                 debug_6_28 /* verilator public */ ;
  reg                 debug_7_28 /* verilator public */ ;
  wire                when_ArraySlice_l158_224;
  wire                when_ArraySlice_l159_224;
  reg        [7:0]    realValue_0_224 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_224;
  wire                when_ArraySlice_l110_224;
  wire                when_ArraySlice_l166_224;
  wire                when_ArraySlice_l158_225;
  wire                when_ArraySlice_l159_225;
  reg        [7:0]    realValue_0_225 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_225;
  wire                when_ArraySlice_l110_225;
  wire                when_ArraySlice_l166_225;
  wire                when_ArraySlice_l158_226;
  wire                when_ArraySlice_l159_226;
  reg        [7:0]    realValue_0_226 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_226;
  wire                when_ArraySlice_l110_226;
  wire                when_ArraySlice_l166_226;
  wire                when_ArraySlice_l158_227;
  wire                when_ArraySlice_l159_227;
  reg        [7:0]    realValue_0_227 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_227;
  wire                when_ArraySlice_l110_227;
  wire                when_ArraySlice_l166_227;
  wire                when_ArraySlice_l158_228;
  wire                when_ArraySlice_l159_228;
  reg        [7:0]    realValue_0_228 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_228;
  wire                when_ArraySlice_l110_228;
  wire                when_ArraySlice_l166_228;
  wire                when_ArraySlice_l158_229;
  wire                when_ArraySlice_l159_229;
  reg        [7:0]    realValue_0_229 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_229;
  wire                when_ArraySlice_l110_229;
  wire                when_ArraySlice_l166_229;
  wire                when_ArraySlice_l158_230;
  wire                when_ArraySlice_l159_230;
  reg        [7:0]    realValue_0_230 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_230;
  wire                when_ArraySlice_l110_230;
  wire                when_ArraySlice_l166_230;
  wire                when_ArraySlice_l158_231;
  wire                when_ArraySlice_l159_231;
  reg        [7:0]    realValue_0_231 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_231;
  wire                when_ArraySlice_l110_231;
  wire                when_ArraySlice_l166_231;
  wire                when_ArraySlice_l314;
  wire                outputStreamArrayData_0_fire_12;
  wire                when_ArraySlice_l318;
  wire                when_ArraySlice_l304;
  wire                outputStreamArrayData_0_fire_13;
  wire                when_ArraySlice_l325;
  wire                when_ArraySlice_l233_1;
  wire                when_ArraySlice_l234_1;
  wire       [7:0]    _zz_outputStreamArrayData_1_valid_1;
  wire                _zz_io_pop_ready_9;
  wire       [127:0]  _zz_12;
  wire                when_ArraySlice_l239_1;
  wire                outputStreamArrayData_1_fire_7;
  wire                when_ArraySlice_l240_1;
  wire                when_ArraySlice_l241_1;
  wire                when_ArraySlice_l244_1;
  wire                outputStreamArrayData_1_fire_8;
  wire                when_ArraySlice_l249_1;
  wire                when_ArraySlice_l250_1;
  reg        [7:0]    realValue1_0_27 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_27;
  wire                when_ArraySlice_l95_27;
  wire                when_ArraySlice_l252_1;
  reg                 debug_0_29 /* verilator public */ ;
  reg                 debug_1_29 /* verilator public */ ;
  reg                 debug_2_29 /* verilator public */ ;
  reg                 debug_3_29 /* verilator public */ ;
  reg                 debug_4_29 /* verilator public */ ;
  reg                 debug_5_29 /* verilator public */ ;
  reg                 debug_6_29 /* verilator public */ ;
  reg                 debug_7_29 /* verilator public */ ;
  wire                when_ArraySlice_l158_232;
  wire                when_ArraySlice_l159_232;
  reg        [7:0]    realValue_0_232 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_232;
  wire                when_ArraySlice_l110_232;
  wire                when_ArraySlice_l166_232;
  wire                when_ArraySlice_l158_233;
  wire                when_ArraySlice_l159_233;
  reg        [7:0]    realValue_0_233 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_233;
  wire                when_ArraySlice_l110_233;
  wire                when_ArraySlice_l166_233;
  wire                when_ArraySlice_l158_234;
  wire                when_ArraySlice_l159_234;
  reg        [7:0]    realValue_0_234 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_234;
  wire                when_ArraySlice_l110_234;
  wire                when_ArraySlice_l166_234;
  wire                when_ArraySlice_l158_235;
  wire                when_ArraySlice_l159_235;
  reg        [7:0]    realValue_0_235 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_235;
  wire                when_ArraySlice_l110_235;
  wire                when_ArraySlice_l166_235;
  wire                when_ArraySlice_l158_236;
  wire                when_ArraySlice_l159_236;
  reg        [7:0]    realValue_0_236 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_236;
  wire                when_ArraySlice_l110_236;
  wire                when_ArraySlice_l166_236;
  wire                when_ArraySlice_l158_237;
  wire                when_ArraySlice_l159_237;
  reg        [7:0]    realValue_0_237 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_237;
  wire                when_ArraySlice_l110_237;
  wire                when_ArraySlice_l166_237;
  wire                when_ArraySlice_l158_238;
  wire                when_ArraySlice_l159_238;
  reg        [7:0]    realValue_0_238 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_238;
  wire                when_ArraySlice_l110_238;
  wire                when_ArraySlice_l166_238;
  wire                when_ArraySlice_l158_239;
  wire                when_ArraySlice_l159_239;
  reg        [7:0]    realValue_0_239 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_239;
  wire                when_ArraySlice_l110_239;
  wire                when_ArraySlice_l166_239;
  wire                when_ArraySlice_l257_1;
  wire                when_ArraySlice_l260_1;
  wire                when_ArraySlice_l263_1;
  wire                when_ArraySlice_l270_1;
  wire                when_ArraySlice_l274_1;
  wire                outputStreamArrayData_1_fire_9;
  wire                when_ArraySlice_l275_1;
  reg        [7:0]    realValue1_0_28 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_28;
  wire                when_ArraySlice_l95_28;
  wire                when_ArraySlice_l277_1;
  reg                 debug_0_30 /* verilator public */ ;
  reg                 debug_1_30 /* verilator public */ ;
  reg                 debug_2_30 /* verilator public */ ;
  reg                 debug_3_30 /* verilator public */ ;
  reg                 debug_4_30 /* verilator public */ ;
  reg                 debug_5_30 /* verilator public */ ;
  reg                 debug_6_30 /* verilator public */ ;
  reg                 debug_7_30 /* verilator public */ ;
  wire                when_ArraySlice_l158_240;
  wire                when_ArraySlice_l159_240;
  reg        [7:0]    realValue_0_240 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_240;
  wire                when_ArraySlice_l110_240;
  wire                when_ArraySlice_l166_240;
  wire                when_ArraySlice_l158_241;
  wire                when_ArraySlice_l159_241;
  reg        [7:0]    realValue_0_241 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_241;
  wire                when_ArraySlice_l110_241;
  wire                when_ArraySlice_l166_241;
  wire                when_ArraySlice_l158_242;
  wire                when_ArraySlice_l159_242;
  reg        [7:0]    realValue_0_242 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_242;
  wire                when_ArraySlice_l110_242;
  wire                when_ArraySlice_l166_242;
  wire                when_ArraySlice_l158_243;
  wire                when_ArraySlice_l159_243;
  reg        [7:0]    realValue_0_243 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_243;
  wire                when_ArraySlice_l110_243;
  wire                when_ArraySlice_l166_243;
  wire                when_ArraySlice_l158_244;
  wire                when_ArraySlice_l159_244;
  reg        [7:0]    realValue_0_244 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_244;
  wire                when_ArraySlice_l110_244;
  wire                when_ArraySlice_l166_244;
  wire                when_ArraySlice_l158_245;
  wire                when_ArraySlice_l159_245;
  reg        [7:0]    realValue_0_245 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_245;
  wire                when_ArraySlice_l110_245;
  wire                when_ArraySlice_l166_245;
  wire                when_ArraySlice_l158_246;
  wire                when_ArraySlice_l159_246;
  reg        [7:0]    realValue_0_246 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_246;
  wire                when_ArraySlice_l110_246;
  wire                when_ArraySlice_l166_246;
  wire                when_ArraySlice_l158_247;
  wire                when_ArraySlice_l159_247;
  reg        [7:0]    realValue_0_247 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_247;
  wire                when_ArraySlice_l110_247;
  wire                when_ArraySlice_l166_247;
  wire                when_ArraySlice_l282_1;
  wire                when_ArraySlice_l285_1;
  wire                when_ArraySlice_l288_1;
  wire                outputStreamArrayData_1_fire_10;
  wire                when_ArraySlice_l295_1;
  wire                outputStreamArrayData_1_fire_11;
  wire                when_ArraySlice_l306_1;
  reg        [7:0]    realValue1_0_29 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_29;
  wire                when_ArraySlice_l95_29;
  wire                when_ArraySlice_l307_1;
  reg                 debug_0_31 /* verilator public */ ;
  reg                 debug_1_31 /* verilator public */ ;
  reg                 debug_2_31 /* verilator public */ ;
  reg                 debug_3_31 /* verilator public */ ;
  reg                 debug_4_31 /* verilator public */ ;
  reg                 debug_5_31 /* verilator public */ ;
  reg                 debug_6_31 /* verilator public */ ;
  reg                 debug_7_31 /* verilator public */ ;
  wire                when_ArraySlice_l158_248;
  wire                when_ArraySlice_l159_248;
  reg        [7:0]    realValue_0_248 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_248;
  wire                when_ArraySlice_l110_248;
  wire                when_ArraySlice_l166_248;
  wire                when_ArraySlice_l158_249;
  wire                when_ArraySlice_l159_249;
  reg        [7:0]    realValue_0_249 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_249;
  wire                when_ArraySlice_l110_249;
  wire                when_ArraySlice_l166_249;
  wire                when_ArraySlice_l158_250;
  wire                when_ArraySlice_l159_250;
  reg        [7:0]    realValue_0_250 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_250;
  wire                when_ArraySlice_l110_250;
  wire                when_ArraySlice_l166_250;
  wire                when_ArraySlice_l158_251;
  wire                when_ArraySlice_l159_251;
  reg        [7:0]    realValue_0_251 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_251;
  wire                when_ArraySlice_l110_251;
  wire                when_ArraySlice_l166_251;
  wire                when_ArraySlice_l158_252;
  wire                when_ArraySlice_l159_252;
  reg        [7:0]    realValue_0_252 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_252;
  wire                when_ArraySlice_l110_252;
  wire                when_ArraySlice_l166_252;
  wire                when_ArraySlice_l158_253;
  wire                when_ArraySlice_l159_253;
  reg        [7:0]    realValue_0_253 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_253;
  wire                when_ArraySlice_l110_253;
  wire                when_ArraySlice_l166_253;
  wire                when_ArraySlice_l158_254;
  wire                when_ArraySlice_l159_254;
  reg        [7:0]    realValue_0_254 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_254;
  wire                when_ArraySlice_l110_254;
  wire                when_ArraySlice_l166_254;
  wire                when_ArraySlice_l158_255;
  wire                when_ArraySlice_l159_255;
  reg        [7:0]    realValue_0_255 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_255;
  wire                when_ArraySlice_l110_255;
  wire                when_ArraySlice_l166_255;
  wire                when_ArraySlice_l314_1;
  wire                outputStreamArrayData_1_fire_12;
  wire                when_ArraySlice_l318_1;
  wire                when_ArraySlice_l304_1;
  wire                outputStreamArrayData_1_fire_13;
  wire                when_ArraySlice_l325_1;
  wire                when_ArraySlice_l233_2;
  wire                when_ArraySlice_l234_2;
  wire       [7:0]    _zz_outputStreamArrayData_2_valid_1;
  wire                _zz_io_pop_ready_10;
  wire       [127:0]  _zz_13;
  wire                when_ArraySlice_l239_2;
  wire                outputStreamArrayData_2_fire_7;
  wire                when_ArraySlice_l240_2;
  wire                when_ArraySlice_l241_2;
  wire                when_ArraySlice_l244_2;
  wire                outputStreamArrayData_2_fire_8;
  wire                when_ArraySlice_l249_2;
  wire                when_ArraySlice_l250_2;
  reg        [7:0]    realValue1_0_30 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_30;
  wire                when_ArraySlice_l95_30;
  wire                when_ArraySlice_l252_2;
  reg                 debug_0_32 /* verilator public */ ;
  reg                 debug_1_32 /* verilator public */ ;
  reg                 debug_2_32 /* verilator public */ ;
  reg                 debug_3_32 /* verilator public */ ;
  reg                 debug_4_32 /* verilator public */ ;
  reg                 debug_5_32 /* verilator public */ ;
  reg                 debug_6_32 /* verilator public */ ;
  reg                 debug_7_32 /* verilator public */ ;
  wire                when_ArraySlice_l158_256;
  wire                when_ArraySlice_l159_256;
  reg        [7:0]    realValue_0_256 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_256;
  wire                when_ArraySlice_l110_256;
  wire                when_ArraySlice_l166_256;
  wire                when_ArraySlice_l158_257;
  wire                when_ArraySlice_l159_257;
  reg        [7:0]    realValue_0_257 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_257;
  wire                when_ArraySlice_l110_257;
  wire                when_ArraySlice_l166_257;
  wire                when_ArraySlice_l158_258;
  wire                when_ArraySlice_l159_258;
  reg        [7:0]    realValue_0_258 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_258;
  wire                when_ArraySlice_l110_258;
  wire                when_ArraySlice_l166_258;
  wire                when_ArraySlice_l158_259;
  wire                when_ArraySlice_l159_259;
  reg        [7:0]    realValue_0_259 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_259;
  wire                when_ArraySlice_l110_259;
  wire                when_ArraySlice_l166_259;
  wire                when_ArraySlice_l158_260;
  wire                when_ArraySlice_l159_260;
  reg        [7:0]    realValue_0_260 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_260;
  wire                when_ArraySlice_l110_260;
  wire                when_ArraySlice_l166_260;
  wire                when_ArraySlice_l158_261;
  wire                when_ArraySlice_l159_261;
  reg        [7:0]    realValue_0_261 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_261;
  wire                when_ArraySlice_l110_261;
  wire                when_ArraySlice_l166_261;
  wire                when_ArraySlice_l158_262;
  wire                when_ArraySlice_l159_262;
  reg        [7:0]    realValue_0_262 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_262;
  wire                when_ArraySlice_l110_262;
  wire                when_ArraySlice_l166_262;
  wire                when_ArraySlice_l158_263;
  wire                when_ArraySlice_l159_263;
  reg        [7:0]    realValue_0_263 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_263;
  wire                when_ArraySlice_l110_263;
  wire                when_ArraySlice_l166_263;
  wire                when_ArraySlice_l257_2;
  wire                when_ArraySlice_l260_2;
  wire                when_ArraySlice_l263_2;
  wire                when_ArraySlice_l270_2;
  wire                when_ArraySlice_l274_2;
  wire                outputStreamArrayData_2_fire_9;
  wire                when_ArraySlice_l275_2;
  reg        [7:0]    realValue1_0_31 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_31;
  wire                when_ArraySlice_l95_31;
  wire                when_ArraySlice_l277_2;
  reg                 debug_0_33 /* verilator public */ ;
  reg                 debug_1_33 /* verilator public */ ;
  reg                 debug_2_33 /* verilator public */ ;
  reg                 debug_3_33 /* verilator public */ ;
  reg                 debug_4_33 /* verilator public */ ;
  reg                 debug_5_33 /* verilator public */ ;
  reg                 debug_6_33 /* verilator public */ ;
  reg                 debug_7_33 /* verilator public */ ;
  wire                when_ArraySlice_l158_264;
  wire                when_ArraySlice_l159_264;
  reg        [7:0]    realValue_0_264 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_264;
  wire                when_ArraySlice_l110_264;
  wire                when_ArraySlice_l166_264;
  wire                when_ArraySlice_l158_265;
  wire                when_ArraySlice_l159_265;
  reg        [7:0]    realValue_0_265 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_265;
  wire                when_ArraySlice_l110_265;
  wire                when_ArraySlice_l166_265;
  wire                when_ArraySlice_l158_266;
  wire                when_ArraySlice_l159_266;
  reg        [7:0]    realValue_0_266 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_266;
  wire                when_ArraySlice_l110_266;
  wire                when_ArraySlice_l166_266;
  wire                when_ArraySlice_l158_267;
  wire                when_ArraySlice_l159_267;
  reg        [7:0]    realValue_0_267 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_267;
  wire                when_ArraySlice_l110_267;
  wire                when_ArraySlice_l166_267;
  wire                when_ArraySlice_l158_268;
  wire                when_ArraySlice_l159_268;
  reg        [7:0]    realValue_0_268 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_268;
  wire                when_ArraySlice_l110_268;
  wire                when_ArraySlice_l166_268;
  wire                when_ArraySlice_l158_269;
  wire                when_ArraySlice_l159_269;
  reg        [7:0]    realValue_0_269 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_269;
  wire                when_ArraySlice_l110_269;
  wire                when_ArraySlice_l166_269;
  wire                when_ArraySlice_l158_270;
  wire                when_ArraySlice_l159_270;
  reg        [7:0]    realValue_0_270 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_270;
  wire                when_ArraySlice_l110_270;
  wire                when_ArraySlice_l166_270;
  wire                when_ArraySlice_l158_271;
  wire                when_ArraySlice_l159_271;
  reg        [7:0]    realValue_0_271 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_271;
  wire                when_ArraySlice_l110_271;
  wire                when_ArraySlice_l166_271;
  wire                when_ArraySlice_l282_2;
  wire                when_ArraySlice_l285_2;
  wire                when_ArraySlice_l288_2;
  wire                outputStreamArrayData_2_fire_10;
  wire                when_ArraySlice_l295_2;
  wire                outputStreamArrayData_2_fire_11;
  wire                when_ArraySlice_l306_2;
  reg        [7:0]    realValue1_0_32 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_32;
  wire                when_ArraySlice_l95_32;
  wire                when_ArraySlice_l307_2;
  reg                 debug_0_34 /* verilator public */ ;
  reg                 debug_1_34 /* verilator public */ ;
  reg                 debug_2_34 /* verilator public */ ;
  reg                 debug_3_34 /* verilator public */ ;
  reg                 debug_4_34 /* verilator public */ ;
  reg                 debug_5_34 /* verilator public */ ;
  reg                 debug_6_34 /* verilator public */ ;
  reg                 debug_7_34 /* verilator public */ ;
  wire                when_ArraySlice_l158_272;
  wire                when_ArraySlice_l159_272;
  reg        [7:0]    realValue_0_272 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_272;
  wire                when_ArraySlice_l110_272;
  wire                when_ArraySlice_l166_272;
  wire                when_ArraySlice_l158_273;
  wire                when_ArraySlice_l159_273;
  reg        [7:0]    realValue_0_273 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_273;
  wire                when_ArraySlice_l110_273;
  wire                when_ArraySlice_l166_273;
  wire                when_ArraySlice_l158_274;
  wire                when_ArraySlice_l159_274;
  reg        [7:0]    realValue_0_274 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_274;
  wire                when_ArraySlice_l110_274;
  wire                when_ArraySlice_l166_274;
  wire                when_ArraySlice_l158_275;
  wire                when_ArraySlice_l159_275;
  reg        [7:0]    realValue_0_275 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_275;
  wire                when_ArraySlice_l110_275;
  wire                when_ArraySlice_l166_275;
  wire                when_ArraySlice_l158_276;
  wire                when_ArraySlice_l159_276;
  reg        [7:0]    realValue_0_276 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_276;
  wire                when_ArraySlice_l110_276;
  wire                when_ArraySlice_l166_276;
  wire                when_ArraySlice_l158_277;
  wire                when_ArraySlice_l159_277;
  reg        [7:0]    realValue_0_277 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_277;
  wire                when_ArraySlice_l110_277;
  wire                when_ArraySlice_l166_277;
  wire                when_ArraySlice_l158_278;
  wire                when_ArraySlice_l159_278;
  reg        [7:0]    realValue_0_278 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_278;
  wire                when_ArraySlice_l110_278;
  wire                when_ArraySlice_l166_278;
  wire                when_ArraySlice_l158_279;
  wire                when_ArraySlice_l159_279;
  reg        [7:0]    realValue_0_279 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_279;
  wire                when_ArraySlice_l110_279;
  wire                when_ArraySlice_l166_279;
  wire                when_ArraySlice_l314_2;
  wire                outputStreamArrayData_2_fire_12;
  wire                when_ArraySlice_l318_2;
  wire                when_ArraySlice_l304_2;
  wire                outputStreamArrayData_2_fire_13;
  wire                when_ArraySlice_l325_2;
  wire                when_ArraySlice_l233_3;
  wire                when_ArraySlice_l234_3;
  wire       [7:0]    _zz_outputStreamArrayData_3_valid_1;
  wire                _zz_io_pop_ready_11;
  wire       [127:0]  _zz_14;
  wire                when_ArraySlice_l239_3;
  wire                outputStreamArrayData_3_fire_7;
  wire                when_ArraySlice_l240_3;
  wire                when_ArraySlice_l241_3;
  wire                when_ArraySlice_l244_3;
  wire                outputStreamArrayData_3_fire_8;
  wire                when_ArraySlice_l249_3;
  wire                when_ArraySlice_l250_3;
  reg        [7:0]    realValue1_0_33 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_33;
  wire                when_ArraySlice_l95_33;
  wire                when_ArraySlice_l252_3;
  reg                 debug_0_35 /* verilator public */ ;
  reg                 debug_1_35 /* verilator public */ ;
  reg                 debug_2_35 /* verilator public */ ;
  reg                 debug_3_35 /* verilator public */ ;
  reg                 debug_4_35 /* verilator public */ ;
  reg                 debug_5_35 /* verilator public */ ;
  reg                 debug_6_35 /* verilator public */ ;
  reg                 debug_7_35 /* verilator public */ ;
  wire                when_ArraySlice_l158_280;
  wire                when_ArraySlice_l159_280;
  reg        [7:0]    realValue_0_280 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_280;
  wire                when_ArraySlice_l110_280;
  wire                when_ArraySlice_l166_280;
  wire                when_ArraySlice_l158_281;
  wire                when_ArraySlice_l159_281;
  reg        [7:0]    realValue_0_281 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_281;
  wire                when_ArraySlice_l110_281;
  wire                when_ArraySlice_l166_281;
  wire                when_ArraySlice_l158_282;
  wire                when_ArraySlice_l159_282;
  reg        [7:0]    realValue_0_282 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_282;
  wire                when_ArraySlice_l110_282;
  wire                when_ArraySlice_l166_282;
  wire                when_ArraySlice_l158_283;
  wire                when_ArraySlice_l159_283;
  reg        [7:0]    realValue_0_283 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_283;
  wire                when_ArraySlice_l110_283;
  wire                when_ArraySlice_l166_283;
  wire                when_ArraySlice_l158_284;
  wire                when_ArraySlice_l159_284;
  reg        [7:0]    realValue_0_284 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_284;
  wire                when_ArraySlice_l110_284;
  wire                when_ArraySlice_l166_284;
  wire                when_ArraySlice_l158_285;
  wire                when_ArraySlice_l159_285;
  reg        [7:0]    realValue_0_285 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_285;
  wire                when_ArraySlice_l110_285;
  wire                when_ArraySlice_l166_285;
  wire                when_ArraySlice_l158_286;
  wire                when_ArraySlice_l159_286;
  reg        [7:0]    realValue_0_286 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_286;
  wire                when_ArraySlice_l110_286;
  wire                when_ArraySlice_l166_286;
  wire                when_ArraySlice_l158_287;
  wire                when_ArraySlice_l159_287;
  reg        [7:0]    realValue_0_287 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_287;
  wire                when_ArraySlice_l110_287;
  wire                when_ArraySlice_l166_287;
  wire                when_ArraySlice_l257_3;
  wire                when_ArraySlice_l260_3;
  wire                when_ArraySlice_l263_3;
  wire                when_ArraySlice_l270_3;
  wire                when_ArraySlice_l274_3;
  wire                outputStreamArrayData_3_fire_9;
  wire                when_ArraySlice_l275_3;
  reg        [7:0]    realValue1_0_34 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_34;
  wire                when_ArraySlice_l95_34;
  wire                when_ArraySlice_l277_3;
  reg                 debug_0_36 /* verilator public */ ;
  reg                 debug_1_36 /* verilator public */ ;
  reg                 debug_2_36 /* verilator public */ ;
  reg                 debug_3_36 /* verilator public */ ;
  reg                 debug_4_36 /* verilator public */ ;
  reg                 debug_5_36 /* verilator public */ ;
  reg                 debug_6_36 /* verilator public */ ;
  reg                 debug_7_36 /* verilator public */ ;
  wire                when_ArraySlice_l158_288;
  wire                when_ArraySlice_l159_288;
  reg        [7:0]    realValue_0_288 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_288;
  wire                when_ArraySlice_l110_288;
  wire                when_ArraySlice_l166_288;
  wire                when_ArraySlice_l158_289;
  wire                when_ArraySlice_l159_289;
  reg        [7:0]    realValue_0_289 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_289;
  wire                when_ArraySlice_l110_289;
  wire                when_ArraySlice_l166_289;
  wire                when_ArraySlice_l158_290;
  wire                when_ArraySlice_l159_290;
  reg        [7:0]    realValue_0_290 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_290;
  wire                when_ArraySlice_l110_290;
  wire                when_ArraySlice_l166_290;
  wire                when_ArraySlice_l158_291;
  wire                when_ArraySlice_l159_291;
  reg        [7:0]    realValue_0_291 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_291;
  wire                when_ArraySlice_l110_291;
  wire                when_ArraySlice_l166_291;
  wire                when_ArraySlice_l158_292;
  wire                when_ArraySlice_l159_292;
  reg        [7:0]    realValue_0_292 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_292;
  wire                when_ArraySlice_l110_292;
  wire                when_ArraySlice_l166_292;
  wire                when_ArraySlice_l158_293;
  wire                when_ArraySlice_l159_293;
  reg        [7:0]    realValue_0_293 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_293;
  wire                when_ArraySlice_l110_293;
  wire                when_ArraySlice_l166_293;
  wire                when_ArraySlice_l158_294;
  wire                when_ArraySlice_l159_294;
  reg        [7:0]    realValue_0_294 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_294;
  wire                when_ArraySlice_l110_294;
  wire                when_ArraySlice_l166_294;
  wire                when_ArraySlice_l158_295;
  wire                when_ArraySlice_l159_295;
  reg        [7:0]    realValue_0_295 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_295;
  wire                when_ArraySlice_l110_295;
  wire                when_ArraySlice_l166_295;
  wire                when_ArraySlice_l282_3;
  wire                when_ArraySlice_l285_3;
  wire                when_ArraySlice_l288_3;
  wire                outputStreamArrayData_3_fire_10;
  wire                when_ArraySlice_l295_3;
  wire                outputStreamArrayData_3_fire_11;
  wire                when_ArraySlice_l306_3;
  reg        [7:0]    realValue1_0_35 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_35;
  wire                when_ArraySlice_l95_35;
  wire                when_ArraySlice_l307_3;
  reg                 debug_0_37 /* verilator public */ ;
  reg                 debug_1_37 /* verilator public */ ;
  reg                 debug_2_37 /* verilator public */ ;
  reg                 debug_3_37 /* verilator public */ ;
  reg                 debug_4_37 /* verilator public */ ;
  reg                 debug_5_37 /* verilator public */ ;
  reg                 debug_6_37 /* verilator public */ ;
  reg                 debug_7_37 /* verilator public */ ;
  wire                when_ArraySlice_l158_296;
  wire                when_ArraySlice_l159_296;
  reg        [7:0]    realValue_0_296 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_296;
  wire                when_ArraySlice_l110_296;
  wire                when_ArraySlice_l166_296;
  wire                when_ArraySlice_l158_297;
  wire                when_ArraySlice_l159_297;
  reg        [7:0]    realValue_0_297 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_297;
  wire                when_ArraySlice_l110_297;
  wire                when_ArraySlice_l166_297;
  wire                when_ArraySlice_l158_298;
  wire                when_ArraySlice_l159_298;
  reg        [7:0]    realValue_0_298 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_298;
  wire                when_ArraySlice_l110_298;
  wire                when_ArraySlice_l166_298;
  wire                when_ArraySlice_l158_299;
  wire                when_ArraySlice_l159_299;
  reg        [7:0]    realValue_0_299 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_299;
  wire                when_ArraySlice_l110_299;
  wire                when_ArraySlice_l166_299;
  wire                when_ArraySlice_l158_300;
  wire                when_ArraySlice_l159_300;
  reg        [7:0]    realValue_0_300 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_300;
  wire                when_ArraySlice_l110_300;
  wire                when_ArraySlice_l166_300;
  wire                when_ArraySlice_l158_301;
  wire                when_ArraySlice_l159_301;
  reg        [7:0]    realValue_0_301 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_301;
  wire                when_ArraySlice_l110_301;
  wire                when_ArraySlice_l166_301;
  wire                when_ArraySlice_l158_302;
  wire                when_ArraySlice_l159_302;
  reg        [7:0]    realValue_0_302 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_302;
  wire                when_ArraySlice_l110_302;
  wire                when_ArraySlice_l166_302;
  wire                when_ArraySlice_l158_303;
  wire                when_ArraySlice_l159_303;
  reg        [7:0]    realValue_0_303 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_303;
  wire                when_ArraySlice_l110_303;
  wire                when_ArraySlice_l166_303;
  wire                when_ArraySlice_l314_3;
  wire                outputStreamArrayData_3_fire_12;
  wire                when_ArraySlice_l318_3;
  wire                when_ArraySlice_l304_3;
  wire                outputStreamArrayData_3_fire_13;
  wire                when_ArraySlice_l325_3;
  wire                when_ArraySlice_l233_4;
  wire                when_ArraySlice_l234_4;
  wire       [7:0]    _zz_outputStreamArrayData_4_valid_1;
  wire                _zz_io_pop_ready_12;
  wire       [127:0]  _zz_15;
  wire                when_ArraySlice_l239_4;
  wire                outputStreamArrayData_4_fire_7;
  wire                when_ArraySlice_l240_4;
  wire                when_ArraySlice_l241_4;
  wire                when_ArraySlice_l244_4;
  wire                outputStreamArrayData_4_fire_8;
  wire                when_ArraySlice_l249_4;
  wire                when_ArraySlice_l250_4;
  reg        [7:0]    realValue1_0_36 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_36;
  wire                when_ArraySlice_l95_36;
  wire                when_ArraySlice_l252_4;
  reg                 debug_0_38 /* verilator public */ ;
  reg                 debug_1_38 /* verilator public */ ;
  reg                 debug_2_38 /* verilator public */ ;
  reg                 debug_3_38 /* verilator public */ ;
  reg                 debug_4_38 /* verilator public */ ;
  reg                 debug_5_38 /* verilator public */ ;
  reg                 debug_6_38 /* verilator public */ ;
  reg                 debug_7_38 /* verilator public */ ;
  wire                when_ArraySlice_l158_304;
  wire                when_ArraySlice_l159_304;
  reg        [7:0]    realValue_0_304 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_304;
  wire                when_ArraySlice_l110_304;
  wire                when_ArraySlice_l166_304;
  wire                when_ArraySlice_l158_305;
  wire                when_ArraySlice_l159_305;
  reg        [7:0]    realValue_0_305 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_305;
  wire                when_ArraySlice_l110_305;
  wire                when_ArraySlice_l166_305;
  wire                when_ArraySlice_l158_306;
  wire                when_ArraySlice_l159_306;
  reg        [7:0]    realValue_0_306 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_306;
  wire                when_ArraySlice_l110_306;
  wire                when_ArraySlice_l166_306;
  wire                when_ArraySlice_l158_307;
  wire                when_ArraySlice_l159_307;
  reg        [7:0]    realValue_0_307 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_307;
  wire                when_ArraySlice_l110_307;
  wire                when_ArraySlice_l166_307;
  wire                when_ArraySlice_l158_308;
  wire                when_ArraySlice_l159_308;
  reg        [7:0]    realValue_0_308 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_308;
  wire                when_ArraySlice_l110_308;
  wire                when_ArraySlice_l166_308;
  wire                when_ArraySlice_l158_309;
  wire                when_ArraySlice_l159_309;
  reg        [7:0]    realValue_0_309 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_309;
  wire                when_ArraySlice_l110_309;
  wire                when_ArraySlice_l166_309;
  wire                when_ArraySlice_l158_310;
  wire                when_ArraySlice_l159_310;
  reg        [7:0]    realValue_0_310 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_310;
  wire                when_ArraySlice_l110_310;
  wire                when_ArraySlice_l166_310;
  wire                when_ArraySlice_l158_311;
  wire                when_ArraySlice_l159_311;
  reg        [7:0]    realValue_0_311 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_311;
  wire                when_ArraySlice_l110_311;
  wire                when_ArraySlice_l166_311;
  wire                when_ArraySlice_l257_4;
  wire                when_ArraySlice_l260_4;
  wire                when_ArraySlice_l263_4;
  wire                when_ArraySlice_l270_4;
  wire                when_ArraySlice_l274_4;
  wire                outputStreamArrayData_4_fire_9;
  wire                when_ArraySlice_l275_4;
  reg        [7:0]    realValue1_0_37 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_37;
  wire                when_ArraySlice_l95_37;
  wire                when_ArraySlice_l277_4;
  reg                 debug_0_39 /* verilator public */ ;
  reg                 debug_1_39 /* verilator public */ ;
  reg                 debug_2_39 /* verilator public */ ;
  reg                 debug_3_39 /* verilator public */ ;
  reg                 debug_4_39 /* verilator public */ ;
  reg                 debug_5_39 /* verilator public */ ;
  reg                 debug_6_39 /* verilator public */ ;
  reg                 debug_7_39 /* verilator public */ ;
  wire                when_ArraySlice_l158_312;
  wire                when_ArraySlice_l159_312;
  reg        [7:0]    realValue_0_312 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_312;
  wire                when_ArraySlice_l110_312;
  wire                when_ArraySlice_l166_312;
  wire                when_ArraySlice_l158_313;
  wire                when_ArraySlice_l159_313;
  reg        [7:0]    realValue_0_313 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_313;
  wire                when_ArraySlice_l110_313;
  wire                when_ArraySlice_l166_313;
  wire                when_ArraySlice_l158_314;
  wire                when_ArraySlice_l159_314;
  reg        [7:0]    realValue_0_314 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_314;
  wire                when_ArraySlice_l110_314;
  wire                when_ArraySlice_l166_314;
  wire                when_ArraySlice_l158_315;
  wire                when_ArraySlice_l159_315;
  reg        [7:0]    realValue_0_315 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_315;
  wire                when_ArraySlice_l110_315;
  wire                when_ArraySlice_l166_315;
  wire                when_ArraySlice_l158_316;
  wire                when_ArraySlice_l159_316;
  reg        [7:0]    realValue_0_316 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_316;
  wire                when_ArraySlice_l110_316;
  wire                when_ArraySlice_l166_316;
  wire                when_ArraySlice_l158_317;
  wire                when_ArraySlice_l159_317;
  reg        [7:0]    realValue_0_317 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_317;
  wire                when_ArraySlice_l110_317;
  wire                when_ArraySlice_l166_317;
  wire                when_ArraySlice_l158_318;
  wire                when_ArraySlice_l159_318;
  reg        [7:0]    realValue_0_318 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_318;
  wire                when_ArraySlice_l110_318;
  wire                when_ArraySlice_l166_318;
  wire                when_ArraySlice_l158_319;
  wire                when_ArraySlice_l159_319;
  reg        [7:0]    realValue_0_319 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_319;
  wire                when_ArraySlice_l110_319;
  wire                when_ArraySlice_l166_319;
  wire                when_ArraySlice_l282_4;
  wire                when_ArraySlice_l285_4;
  wire                when_ArraySlice_l288_4;
  wire                outputStreamArrayData_4_fire_10;
  wire                when_ArraySlice_l295_4;
  wire                outputStreamArrayData_4_fire_11;
  wire                when_ArraySlice_l306_4;
  reg        [7:0]    realValue1_0_38 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_38;
  wire                when_ArraySlice_l95_38;
  wire                when_ArraySlice_l307_4;
  reg                 debug_0_40 /* verilator public */ ;
  reg                 debug_1_40 /* verilator public */ ;
  reg                 debug_2_40 /* verilator public */ ;
  reg                 debug_3_40 /* verilator public */ ;
  reg                 debug_4_40 /* verilator public */ ;
  reg                 debug_5_40 /* verilator public */ ;
  reg                 debug_6_40 /* verilator public */ ;
  reg                 debug_7_40 /* verilator public */ ;
  wire                when_ArraySlice_l158_320;
  wire                when_ArraySlice_l159_320;
  reg        [7:0]    realValue_0_320 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_320;
  wire                when_ArraySlice_l110_320;
  wire                when_ArraySlice_l166_320;
  wire                when_ArraySlice_l158_321;
  wire                when_ArraySlice_l159_321;
  reg        [7:0]    realValue_0_321 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_321;
  wire                when_ArraySlice_l110_321;
  wire                when_ArraySlice_l166_321;
  wire                when_ArraySlice_l158_322;
  wire                when_ArraySlice_l159_322;
  reg        [7:0]    realValue_0_322 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_322;
  wire                when_ArraySlice_l110_322;
  wire                when_ArraySlice_l166_322;
  wire                when_ArraySlice_l158_323;
  wire                when_ArraySlice_l159_323;
  reg        [7:0]    realValue_0_323 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_323;
  wire                when_ArraySlice_l110_323;
  wire                when_ArraySlice_l166_323;
  wire                when_ArraySlice_l158_324;
  wire                when_ArraySlice_l159_324;
  reg        [7:0]    realValue_0_324 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_324;
  wire                when_ArraySlice_l110_324;
  wire                when_ArraySlice_l166_324;
  wire                when_ArraySlice_l158_325;
  wire                when_ArraySlice_l159_325;
  reg        [7:0]    realValue_0_325 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_325;
  wire                when_ArraySlice_l110_325;
  wire                when_ArraySlice_l166_325;
  wire                when_ArraySlice_l158_326;
  wire                when_ArraySlice_l159_326;
  reg        [7:0]    realValue_0_326 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_326;
  wire                when_ArraySlice_l110_326;
  wire                when_ArraySlice_l166_326;
  wire                when_ArraySlice_l158_327;
  wire                when_ArraySlice_l159_327;
  reg        [7:0]    realValue_0_327 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_327;
  wire                when_ArraySlice_l110_327;
  wire                when_ArraySlice_l166_327;
  wire                when_ArraySlice_l314_4;
  wire                outputStreamArrayData_4_fire_12;
  wire                when_ArraySlice_l318_4;
  wire                when_ArraySlice_l304_4;
  wire                outputStreamArrayData_4_fire_13;
  wire                when_ArraySlice_l325_4;
  wire                when_ArraySlice_l233_5;
  wire                when_ArraySlice_l234_5;
  wire       [7:0]    _zz_outputStreamArrayData_5_valid_1;
  wire                _zz_io_pop_ready_13;
  wire       [127:0]  _zz_16;
  wire                when_ArraySlice_l239_5;
  wire                outputStreamArrayData_5_fire_7;
  wire                when_ArraySlice_l240_5;
  wire                when_ArraySlice_l241_5;
  wire                when_ArraySlice_l244_5;
  wire                outputStreamArrayData_5_fire_8;
  wire                when_ArraySlice_l249_5;
  wire                when_ArraySlice_l250_5;
  reg        [7:0]    realValue1_0_39 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_39;
  wire                when_ArraySlice_l95_39;
  wire                when_ArraySlice_l252_5;
  reg                 debug_0_41 /* verilator public */ ;
  reg                 debug_1_41 /* verilator public */ ;
  reg                 debug_2_41 /* verilator public */ ;
  reg                 debug_3_41 /* verilator public */ ;
  reg                 debug_4_41 /* verilator public */ ;
  reg                 debug_5_41 /* verilator public */ ;
  reg                 debug_6_41 /* verilator public */ ;
  reg                 debug_7_41 /* verilator public */ ;
  wire                when_ArraySlice_l158_328;
  wire                when_ArraySlice_l159_328;
  reg        [7:0]    realValue_0_328 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_328;
  wire                when_ArraySlice_l110_328;
  wire                when_ArraySlice_l166_328;
  wire                when_ArraySlice_l158_329;
  wire                when_ArraySlice_l159_329;
  reg        [7:0]    realValue_0_329 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_329;
  wire                when_ArraySlice_l110_329;
  wire                when_ArraySlice_l166_329;
  wire                when_ArraySlice_l158_330;
  wire                when_ArraySlice_l159_330;
  reg        [7:0]    realValue_0_330 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_330;
  wire                when_ArraySlice_l110_330;
  wire                when_ArraySlice_l166_330;
  wire                when_ArraySlice_l158_331;
  wire                when_ArraySlice_l159_331;
  reg        [7:0]    realValue_0_331 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_331;
  wire                when_ArraySlice_l110_331;
  wire                when_ArraySlice_l166_331;
  wire                when_ArraySlice_l158_332;
  wire                when_ArraySlice_l159_332;
  reg        [7:0]    realValue_0_332 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_332;
  wire                when_ArraySlice_l110_332;
  wire                when_ArraySlice_l166_332;
  wire                when_ArraySlice_l158_333;
  wire                when_ArraySlice_l159_333;
  reg        [7:0]    realValue_0_333 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_333;
  wire                when_ArraySlice_l110_333;
  wire                when_ArraySlice_l166_333;
  wire                when_ArraySlice_l158_334;
  wire                when_ArraySlice_l159_334;
  reg        [7:0]    realValue_0_334 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_334;
  wire                when_ArraySlice_l110_334;
  wire                when_ArraySlice_l166_334;
  wire                when_ArraySlice_l158_335;
  wire                when_ArraySlice_l159_335;
  reg        [7:0]    realValue_0_335 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_335;
  wire                when_ArraySlice_l110_335;
  wire                when_ArraySlice_l166_335;
  wire                when_ArraySlice_l257_5;
  wire                when_ArraySlice_l260_5;
  wire                when_ArraySlice_l263_5;
  wire                when_ArraySlice_l270_5;
  wire                when_ArraySlice_l274_5;
  wire                outputStreamArrayData_5_fire_9;
  wire                when_ArraySlice_l275_5;
  reg        [7:0]    realValue1_0_40 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_40;
  wire                when_ArraySlice_l95_40;
  wire                when_ArraySlice_l277_5;
  reg                 debug_0_42 /* verilator public */ ;
  reg                 debug_1_42 /* verilator public */ ;
  reg                 debug_2_42 /* verilator public */ ;
  reg                 debug_3_42 /* verilator public */ ;
  reg                 debug_4_42 /* verilator public */ ;
  reg                 debug_5_42 /* verilator public */ ;
  reg                 debug_6_42 /* verilator public */ ;
  reg                 debug_7_42 /* verilator public */ ;
  wire                when_ArraySlice_l158_336;
  wire                when_ArraySlice_l159_336;
  reg        [7:0]    realValue_0_336 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_336;
  wire                when_ArraySlice_l110_336;
  wire                when_ArraySlice_l166_336;
  wire                when_ArraySlice_l158_337;
  wire                when_ArraySlice_l159_337;
  reg        [7:0]    realValue_0_337 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_337;
  wire                when_ArraySlice_l110_337;
  wire                when_ArraySlice_l166_337;
  wire                when_ArraySlice_l158_338;
  wire                when_ArraySlice_l159_338;
  reg        [7:0]    realValue_0_338 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_338;
  wire                when_ArraySlice_l110_338;
  wire                when_ArraySlice_l166_338;
  wire                when_ArraySlice_l158_339;
  wire                when_ArraySlice_l159_339;
  reg        [7:0]    realValue_0_339 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_339;
  wire                when_ArraySlice_l110_339;
  wire                when_ArraySlice_l166_339;
  wire                when_ArraySlice_l158_340;
  wire                when_ArraySlice_l159_340;
  reg        [7:0]    realValue_0_340 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_340;
  wire                when_ArraySlice_l110_340;
  wire                when_ArraySlice_l166_340;
  wire                when_ArraySlice_l158_341;
  wire                when_ArraySlice_l159_341;
  reg        [7:0]    realValue_0_341 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_341;
  wire                when_ArraySlice_l110_341;
  wire                when_ArraySlice_l166_341;
  wire                when_ArraySlice_l158_342;
  wire                when_ArraySlice_l159_342;
  reg        [7:0]    realValue_0_342 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_342;
  wire                when_ArraySlice_l110_342;
  wire                when_ArraySlice_l166_342;
  wire                when_ArraySlice_l158_343;
  wire                when_ArraySlice_l159_343;
  reg        [7:0]    realValue_0_343 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_343;
  wire                when_ArraySlice_l110_343;
  wire                when_ArraySlice_l166_343;
  wire                when_ArraySlice_l282_5;
  wire                when_ArraySlice_l285_5;
  wire                when_ArraySlice_l288_5;
  wire                outputStreamArrayData_5_fire_10;
  wire                when_ArraySlice_l295_5;
  wire                outputStreamArrayData_5_fire_11;
  wire                when_ArraySlice_l306_5;
  reg        [7:0]    realValue1_0_41 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_41;
  wire                when_ArraySlice_l95_41;
  wire                when_ArraySlice_l307_5;
  reg                 debug_0_43 /* verilator public */ ;
  reg                 debug_1_43 /* verilator public */ ;
  reg                 debug_2_43 /* verilator public */ ;
  reg                 debug_3_43 /* verilator public */ ;
  reg                 debug_4_43 /* verilator public */ ;
  reg                 debug_5_43 /* verilator public */ ;
  reg                 debug_6_43 /* verilator public */ ;
  reg                 debug_7_43 /* verilator public */ ;
  wire                when_ArraySlice_l158_344;
  wire                when_ArraySlice_l159_344;
  reg        [7:0]    realValue_0_344 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_344;
  wire                when_ArraySlice_l110_344;
  wire                when_ArraySlice_l166_344;
  wire                when_ArraySlice_l158_345;
  wire                when_ArraySlice_l159_345;
  reg        [7:0]    realValue_0_345 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_345;
  wire                when_ArraySlice_l110_345;
  wire                when_ArraySlice_l166_345;
  wire                when_ArraySlice_l158_346;
  wire                when_ArraySlice_l159_346;
  reg        [7:0]    realValue_0_346 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_346;
  wire                when_ArraySlice_l110_346;
  wire                when_ArraySlice_l166_346;
  wire                when_ArraySlice_l158_347;
  wire                when_ArraySlice_l159_347;
  reg        [7:0]    realValue_0_347 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_347;
  wire                when_ArraySlice_l110_347;
  wire                when_ArraySlice_l166_347;
  wire                when_ArraySlice_l158_348;
  wire                when_ArraySlice_l159_348;
  reg        [7:0]    realValue_0_348 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_348;
  wire                when_ArraySlice_l110_348;
  wire                when_ArraySlice_l166_348;
  wire                when_ArraySlice_l158_349;
  wire                when_ArraySlice_l159_349;
  reg        [7:0]    realValue_0_349 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_349;
  wire                when_ArraySlice_l110_349;
  wire                when_ArraySlice_l166_349;
  wire                when_ArraySlice_l158_350;
  wire                when_ArraySlice_l159_350;
  reg        [7:0]    realValue_0_350 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_350;
  wire                when_ArraySlice_l110_350;
  wire                when_ArraySlice_l166_350;
  wire                when_ArraySlice_l158_351;
  wire                when_ArraySlice_l159_351;
  reg        [7:0]    realValue_0_351 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_351;
  wire                when_ArraySlice_l110_351;
  wire                when_ArraySlice_l166_351;
  wire                when_ArraySlice_l314_5;
  wire                outputStreamArrayData_5_fire_12;
  wire                when_ArraySlice_l318_5;
  wire                when_ArraySlice_l304_5;
  wire                outputStreamArrayData_5_fire_13;
  wire                when_ArraySlice_l325_5;
  wire                when_ArraySlice_l233_6;
  wire                when_ArraySlice_l234_6;
  wire       [7:0]    _zz_outputStreamArrayData_6_valid_1;
  wire                _zz_io_pop_ready_14;
  wire       [127:0]  _zz_17;
  wire                when_ArraySlice_l239_6;
  wire                outputStreamArrayData_6_fire_7;
  wire                when_ArraySlice_l240_6;
  wire                when_ArraySlice_l241_6;
  wire                when_ArraySlice_l244_6;
  wire                outputStreamArrayData_6_fire_8;
  wire                when_ArraySlice_l249_6;
  wire                when_ArraySlice_l250_6;
  reg        [7:0]    realValue1_0_42 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_42;
  wire                when_ArraySlice_l95_42;
  wire                when_ArraySlice_l252_6;
  reg                 debug_0_44 /* verilator public */ ;
  reg                 debug_1_44 /* verilator public */ ;
  reg                 debug_2_44 /* verilator public */ ;
  reg                 debug_3_44 /* verilator public */ ;
  reg                 debug_4_44 /* verilator public */ ;
  reg                 debug_5_44 /* verilator public */ ;
  reg                 debug_6_44 /* verilator public */ ;
  reg                 debug_7_44 /* verilator public */ ;
  wire                when_ArraySlice_l158_352;
  wire                when_ArraySlice_l159_352;
  reg        [7:0]    realValue_0_352 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_352;
  wire                when_ArraySlice_l110_352;
  wire                when_ArraySlice_l166_352;
  wire                when_ArraySlice_l158_353;
  wire                when_ArraySlice_l159_353;
  reg        [7:0]    realValue_0_353 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_353;
  wire                when_ArraySlice_l110_353;
  wire                when_ArraySlice_l166_353;
  wire                when_ArraySlice_l158_354;
  wire                when_ArraySlice_l159_354;
  reg        [7:0]    realValue_0_354 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_354;
  wire                when_ArraySlice_l110_354;
  wire                when_ArraySlice_l166_354;
  wire                when_ArraySlice_l158_355;
  wire                when_ArraySlice_l159_355;
  reg        [7:0]    realValue_0_355 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_355;
  wire                when_ArraySlice_l110_355;
  wire                when_ArraySlice_l166_355;
  wire                when_ArraySlice_l158_356;
  wire                when_ArraySlice_l159_356;
  reg        [7:0]    realValue_0_356 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_356;
  wire                when_ArraySlice_l110_356;
  wire                when_ArraySlice_l166_356;
  wire                when_ArraySlice_l158_357;
  wire                when_ArraySlice_l159_357;
  reg        [7:0]    realValue_0_357 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_357;
  wire                when_ArraySlice_l110_357;
  wire                when_ArraySlice_l166_357;
  wire                when_ArraySlice_l158_358;
  wire                when_ArraySlice_l159_358;
  reg        [7:0]    realValue_0_358 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_358;
  wire                when_ArraySlice_l110_358;
  wire                when_ArraySlice_l166_358;
  wire                when_ArraySlice_l158_359;
  wire                when_ArraySlice_l159_359;
  reg        [7:0]    realValue_0_359 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_359;
  wire                when_ArraySlice_l110_359;
  wire                when_ArraySlice_l166_359;
  wire                when_ArraySlice_l257_6;
  wire                when_ArraySlice_l260_6;
  wire                when_ArraySlice_l263_6;
  wire                when_ArraySlice_l270_6;
  wire                when_ArraySlice_l274_6;
  wire                outputStreamArrayData_6_fire_9;
  wire                when_ArraySlice_l275_6;
  reg        [7:0]    realValue1_0_43 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_43;
  wire                when_ArraySlice_l95_43;
  wire                when_ArraySlice_l277_6;
  reg                 debug_0_45 /* verilator public */ ;
  reg                 debug_1_45 /* verilator public */ ;
  reg                 debug_2_45 /* verilator public */ ;
  reg                 debug_3_45 /* verilator public */ ;
  reg                 debug_4_45 /* verilator public */ ;
  reg                 debug_5_45 /* verilator public */ ;
  reg                 debug_6_45 /* verilator public */ ;
  reg                 debug_7_45 /* verilator public */ ;
  wire                when_ArraySlice_l158_360;
  wire                when_ArraySlice_l159_360;
  reg        [7:0]    realValue_0_360 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_360;
  wire                when_ArraySlice_l110_360;
  wire                when_ArraySlice_l166_360;
  wire                when_ArraySlice_l158_361;
  wire                when_ArraySlice_l159_361;
  reg        [7:0]    realValue_0_361 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_361;
  wire                when_ArraySlice_l110_361;
  wire                when_ArraySlice_l166_361;
  wire                when_ArraySlice_l158_362;
  wire                when_ArraySlice_l159_362;
  reg        [7:0]    realValue_0_362 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_362;
  wire                when_ArraySlice_l110_362;
  wire                when_ArraySlice_l166_362;
  wire                when_ArraySlice_l158_363;
  wire                when_ArraySlice_l159_363;
  reg        [7:0]    realValue_0_363 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_363;
  wire                when_ArraySlice_l110_363;
  wire                when_ArraySlice_l166_363;
  wire                when_ArraySlice_l158_364;
  wire                when_ArraySlice_l159_364;
  reg        [7:0]    realValue_0_364 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_364;
  wire                when_ArraySlice_l110_364;
  wire                when_ArraySlice_l166_364;
  wire                when_ArraySlice_l158_365;
  wire                when_ArraySlice_l159_365;
  reg        [7:0]    realValue_0_365 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_365;
  wire                when_ArraySlice_l110_365;
  wire                when_ArraySlice_l166_365;
  wire                when_ArraySlice_l158_366;
  wire                when_ArraySlice_l159_366;
  reg        [7:0]    realValue_0_366 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_366;
  wire                when_ArraySlice_l110_366;
  wire                when_ArraySlice_l166_366;
  wire                when_ArraySlice_l158_367;
  wire                when_ArraySlice_l159_367;
  reg        [7:0]    realValue_0_367 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_367;
  wire                when_ArraySlice_l110_367;
  wire                when_ArraySlice_l166_367;
  wire                when_ArraySlice_l282_6;
  wire                when_ArraySlice_l285_6;
  wire                when_ArraySlice_l288_6;
  wire                outputStreamArrayData_6_fire_10;
  wire                when_ArraySlice_l295_6;
  wire                outputStreamArrayData_6_fire_11;
  wire                when_ArraySlice_l306_6;
  reg        [7:0]    realValue1_0_44 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_44;
  wire                when_ArraySlice_l95_44;
  wire                when_ArraySlice_l307_6;
  reg                 debug_0_46 /* verilator public */ ;
  reg                 debug_1_46 /* verilator public */ ;
  reg                 debug_2_46 /* verilator public */ ;
  reg                 debug_3_46 /* verilator public */ ;
  reg                 debug_4_46 /* verilator public */ ;
  reg                 debug_5_46 /* verilator public */ ;
  reg                 debug_6_46 /* verilator public */ ;
  reg                 debug_7_46 /* verilator public */ ;
  wire                when_ArraySlice_l158_368;
  wire                when_ArraySlice_l159_368;
  reg        [7:0]    realValue_0_368 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_368;
  wire                when_ArraySlice_l110_368;
  wire                when_ArraySlice_l166_368;
  wire                when_ArraySlice_l158_369;
  wire                when_ArraySlice_l159_369;
  reg        [7:0]    realValue_0_369 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_369;
  wire                when_ArraySlice_l110_369;
  wire                when_ArraySlice_l166_369;
  wire                when_ArraySlice_l158_370;
  wire                when_ArraySlice_l159_370;
  reg        [7:0]    realValue_0_370 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_370;
  wire                when_ArraySlice_l110_370;
  wire                when_ArraySlice_l166_370;
  wire                when_ArraySlice_l158_371;
  wire                when_ArraySlice_l159_371;
  reg        [7:0]    realValue_0_371 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_371;
  wire                when_ArraySlice_l110_371;
  wire                when_ArraySlice_l166_371;
  wire                when_ArraySlice_l158_372;
  wire                when_ArraySlice_l159_372;
  reg        [7:0]    realValue_0_372 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_372;
  wire                when_ArraySlice_l110_372;
  wire                when_ArraySlice_l166_372;
  wire                when_ArraySlice_l158_373;
  wire                when_ArraySlice_l159_373;
  reg        [7:0]    realValue_0_373 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_373;
  wire                when_ArraySlice_l110_373;
  wire                when_ArraySlice_l166_373;
  wire                when_ArraySlice_l158_374;
  wire                when_ArraySlice_l159_374;
  reg        [7:0]    realValue_0_374 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_374;
  wire                when_ArraySlice_l110_374;
  wire                when_ArraySlice_l166_374;
  wire                when_ArraySlice_l158_375;
  wire                when_ArraySlice_l159_375;
  reg        [7:0]    realValue_0_375 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_375;
  wire                when_ArraySlice_l110_375;
  wire                when_ArraySlice_l166_375;
  wire                when_ArraySlice_l314_6;
  wire                outputStreamArrayData_6_fire_12;
  wire                when_ArraySlice_l318_6;
  wire                when_ArraySlice_l304_6;
  wire                outputStreamArrayData_6_fire_13;
  wire                when_ArraySlice_l325_6;
  wire                when_ArraySlice_l233_7;
  wire                when_ArraySlice_l234_7;
  wire       [7:0]    _zz_outputStreamArrayData_7_valid_1;
  wire                _zz_io_pop_ready_15;
  wire       [127:0]  _zz_18;
  wire                when_ArraySlice_l239_7;
  wire                outputStreamArrayData_7_fire_7;
  wire                when_ArraySlice_l240_7;
  wire                when_ArraySlice_l241_7;
  wire                when_ArraySlice_l244_7;
  wire                outputStreamArrayData_7_fire_8;
  wire                when_ArraySlice_l249_7;
  wire                when_ArraySlice_l250_7;
  reg        [7:0]    realValue1_0_45 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_45;
  wire                when_ArraySlice_l95_45;
  wire                when_ArraySlice_l252_7;
  reg                 debug_0_47 /* verilator public */ ;
  reg                 debug_1_47 /* verilator public */ ;
  reg                 debug_2_47 /* verilator public */ ;
  reg                 debug_3_47 /* verilator public */ ;
  reg                 debug_4_47 /* verilator public */ ;
  reg                 debug_5_47 /* verilator public */ ;
  reg                 debug_6_47 /* verilator public */ ;
  reg                 debug_7_47 /* verilator public */ ;
  wire                when_ArraySlice_l158_376;
  wire                when_ArraySlice_l159_376;
  reg        [7:0]    realValue_0_376 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_376;
  wire                when_ArraySlice_l110_376;
  wire                when_ArraySlice_l166_376;
  wire                when_ArraySlice_l158_377;
  wire                when_ArraySlice_l159_377;
  reg        [7:0]    realValue_0_377 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_377;
  wire                when_ArraySlice_l110_377;
  wire                when_ArraySlice_l166_377;
  wire                when_ArraySlice_l158_378;
  wire                when_ArraySlice_l159_378;
  reg        [7:0]    realValue_0_378 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_378;
  wire                when_ArraySlice_l110_378;
  wire                when_ArraySlice_l166_378;
  wire                when_ArraySlice_l158_379;
  wire                when_ArraySlice_l159_379;
  reg        [7:0]    realValue_0_379 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_379;
  wire                when_ArraySlice_l110_379;
  wire                when_ArraySlice_l166_379;
  wire                when_ArraySlice_l158_380;
  wire                when_ArraySlice_l159_380;
  reg        [7:0]    realValue_0_380 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_380;
  wire                when_ArraySlice_l110_380;
  wire                when_ArraySlice_l166_380;
  wire                when_ArraySlice_l158_381;
  wire                when_ArraySlice_l159_381;
  reg        [7:0]    realValue_0_381 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_381;
  wire                when_ArraySlice_l110_381;
  wire                when_ArraySlice_l166_381;
  wire                when_ArraySlice_l158_382;
  wire                when_ArraySlice_l159_382;
  reg        [7:0]    realValue_0_382 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_382;
  wire                when_ArraySlice_l110_382;
  wire                when_ArraySlice_l166_382;
  wire                when_ArraySlice_l158_383;
  wire                when_ArraySlice_l159_383;
  reg        [7:0]    realValue_0_383 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_383;
  wire                when_ArraySlice_l110_383;
  wire                when_ArraySlice_l166_383;
  wire                when_ArraySlice_l257_7;
  wire                when_ArraySlice_l260_7;
  wire                when_ArraySlice_l263_7;
  wire                when_ArraySlice_l270_7;
  wire                when_ArraySlice_l274_7;
  wire                outputStreamArrayData_7_fire_9;
  wire                when_ArraySlice_l275_7;
  reg        [7:0]    realValue1_0_46 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_46;
  wire                when_ArraySlice_l95_46;
  wire                when_ArraySlice_l277_7;
  reg                 debug_0_48 /* verilator public */ ;
  reg                 debug_1_48 /* verilator public */ ;
  reg                 debug_2_48 /* verilator public */ ;
  reg                 debug_3_48 /* verilator public */ ;
  reg                 debug_4_48 /* verilator public */ ;
  reg                 debug_5_48 /* verilator public */ ;
  reg                 debug_6_48 /* verilator public */ ;
  reg                 debug_7_48 /* verilator public */ ;
  wire                when_ArraySlice_l158_384;
  wire                when_ArraySlice_l159_384;
  reg        [7:0]    realValue_0_384 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_384;
  wire                when_ArraySlice_l110_384;
  wire                when_ArraySlice_l166_384;
  wire                when_ArraySlice_l158_385;
  wire                when_ArraySlice_l159_385;
  reg        [7:0]    realValue_0_385 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_385;
  wire                when_ArraySlice_l110_385;
  wire                when_ArraySlice_l166_385;
  wire                when_ArraySlice_l158_386;
  wire                when_ArraySlice_l159_386;
  reg        [7:0]    realValue_0_386 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_386;
  wire                when_ArraySlice_l110_386;
  wire                when_ArraySlice_l166_386;
  wire                when_ArraySlice_l158_387;
  wire                when_ArraySlice_l159_387;
  reg        [7:0]    realValue_0_387 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_387;
  wire                when_ArraySlice_l110_387;
  wire                when_ArraySlice_l166_387;
  wire                when_ArraySlice_l158_388;
  wire                when_ArraySlice_l159_388;
  reg        [7:0]    realValue_0_388 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_388;
  wire                when_ArraySlice_l110_388;
  wire                when_ArraySlice_l166_388;
  wire                when_ArraySlice_l158_389;
  wire                when_ArraySlice_l159_389;
  reg        [7:0]    realValue_0_389 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_389;
  wire                when_ArraySlice_l110_389;
  wire                when_ArraySlice_l166_389;
  wire                when_ArraySlice_l158_390;
  wire                when_ArraySlice_l159_390;
  reg        [7:0]    realValue_0_390 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_390;
  wire                when_ArraySlice_l110_390;
  wire                when_ArraySlice_l166_390;
  wire                when_ArraySlice_l158_391;
  wire                when_ArraySlice_l159_391;
  reg        [7:0]    realValue_0_391 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_391;
  wire                when_ArraySlice_l110_391;
  wire                when_ArraySlice_l166_391;
  wire                when_ArraySlice_l282_7;
  wire                when_ArraySlice_l285_7;
  wire                when_ArraySlice_l288_7;
  wire                outputStreamArrayData_7_fire_10;
  wire                when_ArraySlice_l295_7;
  wire                outputStreamArrayData_7_fire_11;
  wire                when_ArraySlice_l306_7;
  reg        [7:0]    realValue1_0_47 /* verilator public */ ;
  wire       [7:0]    _zz_realValue1_0_47;
  wire                when_ArraySlice_l95_47;
  wire                when_ArraySlice_l307_7;
  reg                 debug_0_49 /* verilator public */ ;
  reg                 debug_1_49 /* verilator public */ ;
  reg                 debug_2_49 /* verilator public */ ;
  reg                 debug_3_49 /* verilator public */ ;
  reg                 debug_4_49 /* verilator public */ ;
  reg                 debug_5_49 /* verilator public */ ;
  reg                 debug_6_49 /* verilator public */ ;
  reg                 debug_7_49 /* verilator public */ ;
  wire                when_ArraySlice_l158_392;
  wire                when_ArraySlice_l159_392;
  reg        [7:0]    realValue_0_392 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_392;
  wire                when_ArraySlice_l110_392;
  wire                when_ArraySlice_l166_392;
  wire                when_ArraySlice_l158_393;
  wire                when_ArraySlice_l159_393;
  reg        [7:0]    realValue_0_393 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_393;
  wire                when_ArraySlice_l110_393;
  wire                when_ArraySlice_l166_393;
  wire                when_ArraySlice_l158_394;
  wire                when_ArraySlice_l159_394;
  reg        [7:0]    realValue_0_394 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_394;
  wire                when_ArraySlice_l110_394;
  wire                when_ArraySlice_l166_394;
  wire                when_ArraySlice_l158_395;
  wire                when_ArraySlice_l159_395;
  reg        [7:0]    realValue_0_395 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_395;
  wire                when_ArraySlice_l110_395;
  wire                when_ArraySlice_l166_395;
  wire                when_ArraySlice_l158_396;
  wire                when_ArraySlice_l159_396;
  reg        [7:0]    realValue_0_396 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_396;
  wire                when_ArraySlice_l110_396;
  wire                when_ArraySlice_l166_396;
  wire                when_ArraySlice_l158_397;
  wire                when_ArraySlice_l159_397;
  reg        [7:0]    realValue_0_397 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_397;
  wire                when_ArraySlice_l110_397;
  wire                when_ArraySlice_l166_397;
  wire                when_ArraySlice_l158_398;
  wire                when_ArraySlice_l159_398;
  reg        [7:0]    realValue_0_398 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_398;
  wire                when_ArraySlice_l110_398;
  wire                when_ArraySlice_l166_398;
  wire                when_ArraySlice_l158_399;
  wire                when_ArraySlice_l159_399;
  reg        [7:0]    realValue_0_399 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_399;
  wire                when_ArraySlice_l110_399;
  wire                when_ArraySlice_l166_399;
  wire                when_ArraySlice_l314_7;
  wire                outputStreamArrayData_7_fire_12;
  wire                when_ArraySlice_l318_7;
  wire                when_ArraySlice_l304_7;
  wire                outputStreamArrayData_7_fire_13;
  wire                when_ArraySlice_l325_7;
  reg                 _zz_when_ArraySlice_l336;
  reg                 _zz_when_ArraySlice_l336_1;
  reg                 _zz_when_ArraySlice_l336_2;
  reg                 _zz_when_ArraySlice_l336_3;
  reg                 _zz_when_ArraySlice_l336_4;
  reg                 _zz_when_ArraySlice_l336_5;
  reg                 _zz_when_ArraySlice_l336_6;
  reg                 _zz_when_ArraySlice_l336_7;
  wire                when_ArraySlice_l182;
  wire                when_ArraySlice_l183;
  wire                when_ArraySlice_l182_1;
  wire                when_ArraySlice_l183_1;
  wire                when_ArraySlice_l182_2;
  wire                when_ArraySlice_l183_2;
  wire                when_ArraySlice_l182_3;
  wire                when_ArraySlice_l183_3;
  wire                when_ArraySlice_l182_4;
  wire                when_ArraySlice_l183_4;
  wire                when_ArraySlice_l182_5;
  wire                when_ArraySlice_l183_5;
  wire                when_ArraySlice_l182_6;
  wire                when_ArraySlice_l183_6;
  wire                when_ArraySlice_l182_7;
  wire                when_ArraySlice_l183_7;
  wire                when_ArraySlice_l336;
  wire                when_ArraySlice_l337;
  wire                _zz_io_push_valid_1;
  wire       [31:0]   _zz_io_push_payload_1;
  wire       [127:0]  _zz_19;
  wire       [127:0]  _zz_20;
  wire                inputStreamArrayData_fire_1;
  wire                when_ArraySlice_l341;
  wire                when_ArraySlice_l342;
  reg                 debug_0_50 /* verilator public */ ;
  reg                 debug_1_50 /* verilator public */ ;
  reg                 debug_2_50 /* verilator public */ ;
  reg                 debug_3_50 /* verilator public */ ;
  reg                 debug_4_50 /* verilator public */ ;
  reg                 debug_5_50 /* verilator public */ ;
  reg                 debug_6_50 /* verilator public */ ;
  reg                 debug_7_50 /* verilator public */ ;
  wire                when_ArraySlice_l158_400;
  wire                when_ArraySlice_l159_400;
  reg        [7:0]    realValue_0_400 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_400;
  wire                when_ArraySlice_l110_400;
  wire                when_ArraySlice_l166_400;
  wire                when_ArraySlice_l158_401;
  wire                when_ArraySlice_l159_401;
  reg        [7:0]    realValue_0_401 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_401;
  wire                when_ArraySlice_l110_401;
  wire                when_ArraySlice_l166_401;
  wire                when_ArraySlice_l158_402;
  wire                when_ArraySlice_l159_402;
  reg        [7:0]    realValue_0_402 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_402;
  wire                when_ArraySlice_l110_402;
  wire                when_ArraySlice_l166_402;
  wire                when_ArraySlice_l158_403;
  wire                when_ArraySlice_l159_403;
  reg        [7:0]    realValue_0_403 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_403;
  wire                when_ArraySlice_l110_403;
  wire                when_ArraySlice_l166_403;
  wire                when_ArraySlice_l158_404;
  wire                when_ArraySlice_l159_404;
  reg        [7:0]    realValue_0_404 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_404;
  wire                when_ArraySlice_l110_404;
  wire                when_ArraySlice_l166_404;
  wire                when_ArraySlice_l158_405;
  wire                when_ArraySlice_l159_405;
  reg        [7:0]    realValue_0_405 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_405;
  wire                when_ArraySlice_l110_405;
  wire                when_ArraySlice_l166_405;
  wire                when_ArraySlice_l158_406;
  wire                when_ArraySlice_l159_406;
  reg        [7:0]    realValue_0_406 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_406;
  wire                when_ArraySlice_l110_406;
  wire                when_ArraySlice_l166_406;
  wire                when_ArraySlice_l158_407;
  wire                when_ArraySlice_l159_407;
  reg        [7:0]    realValue_0_407 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_407;
  wire                when_ArraySlice_l110_407;
  wire                when_ArraySlice_l166_407;
  wire                when_ArraySlice_l353;
  reg                 debug_0_51 /* verilator public */ ;
  reg                 debug_1_51 /* verilator public */ ;
  reg                 debug_2_51 /* verilator public */ ;
  reg                 debug_3_51 /* verilator public */ ;
  reg                 debug_4_51 /* verilator public */ ;
  reg                 debug_5_51 /* verilator public */ ;
  reg                 debug_6_51 /* verilator public */ ;
  reg                 debug_7_51 /* verilator public */ ;
  wire                when_ArraySlice_l158_408;
  wire                when_ArraySlice_l159_408;
  reg        [7:0]    realValue_0_408 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_408;
  wire                when_ArraySlice_l110_408;
  wire                when_ArraySlice_l166_408;
  wire                when_ArraySlice_l158_409;
  wire                when_ArraySlice_l159_409;
  reg        [7:0]    realValue_0_409 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_409;
  wire                when_ArraySlice_l110_409;
  wire                when_ArraySlice_l166_409;
  wire                when_ArraySlice_l158_410;
  wire                when_ArraySlice_l159_410;
  reg        [7:0]    realValue_0_410 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_410;
  wire                when_ArraySlice_l110_410;
  wire                when_ArraySlice_l166_410;
  wire                when_ArraySlice_l158_411;
  wire                when_ArraySlice_l159_411;
  reg        [7:0]    realValue_0_411 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_411;
  wire                when_ArraySlice_l110_411;
  wire                when_ArraySlice_l166_411;
  wire                when_ArraySlice_l158_412;
  wire                when_ArraySlice_l159_412;
  reg        [7:0]    realValue_0_412 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_412;
  wire                when_ArraySlice_l110_412;
  wire                when_ArraySlice_l166_412;
  wire                when_ArraySlice_l158_413;
  wire                when_ArraySlice_l159_413;
  reg        [7:0]    realValue_0_413 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_413;
  wire                when_ArraySlice_l110_413;
  wire                when_ArraySlice_l166_413;
  wire                when_ArraySlice_l158_414;
  wire                when_ArraySlice_l159_414;
  reg        [7:0]    realValue_0_414 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_414;
  wire                when_ArraySlice_l110_414;
  wire                when_ArraySlice_l166_414;
  wire                when_ArraySlice_l158_415;
  wire                when_ArraySlice_l159_415;
  reg        [7:0]    realValue_0_415 /* verilator public */ ;
  wire       [7:0]    _zz_realValue_0_415;
  wire                when_ArraySlice_l110_415;
  wire                when_ArraySlice_l166_415;
  reg                 _zz_when_ArraySlice_l357;
  reg                 _zz_when_ArraySlice_l357_1;
  reg                 _zz_when_ArraySlice_l357_2;
  reg                 _zz_when_ArraySlice_l357_3;
  reg                 _zz_when_ArraySlice_l357_4;
  reg                 _zz_when_ArraySlice_l357_5;
  reg                 _zz_when_ArraySlice_l357_6;
  reg                 _zz_when_ArraySlice_l357_7;
  wire                when_ArraySlice_l182_8;
  wire                when_ArraySlice_l183_8;
  wire                when_ArraySlice_l182_9;
  wire                when_ArraySlice_l183_9;
  wire                when_ArraySlice_l182_10;
  wire                when_ArraySlice_l183_10;
  wire                when_ArraySlice_l182_11;
  wire                when_ArraySlice_l183_11;
  wire                when_ArraySlice_l182_12;
  wire                when_ArraySlice_l183_12;
  wire                when_ArraySlice_l182_13;
  wire                when_ArraySlice_l183_13;
  wire                when_ArraySlice_l182_14;
  wire                when_ArraySlice_l183_14;
  wire                when_ArraySlice_l182_15;
  wire                when_ArraySlice_l183_15;
  wire                when_ArraySlice_l357;
  reg                 _zz_when_ArraySlice_l361;
  reg                 _zz_when_ArraySlice_l361_1;
  reg                 _zz_when_ArraySlice_l361_2;
  reg                 _zz_when_ArraySlice_l361_3;
  reg                 _zz_when_ArraySlice_l361_4;
  reg                 _zz_when_ArraySlice_l361_5;
  reg                 _zz_when_ArraySlice_l361_6;
  reg                 _zz_when_ArraySlice_l361_7;
  wire                when_ArraySlice_l182_16;
  wire                when_ArraySlice_l183_16;
  wire                when_ArraySlice_l182_17;
  wire                when_ArraySlice_l183_17;
  wire                when_ArraySlice_l182_18;
  wire                when_ArraySlice_l183_18;
  wire                when_ArraySlice_l182_19;
  wire                when_ArraySlice_l183_19;
  wire                when_ArraySlice_l182_20;
  wire                when_ArraySlice_l183_20;
  wire                when_ArraySlice_l182_21;
  wire                when_ArraySlice_l183_21;
  wire                when_ArraySlice_l182_22;
  wire                when_ArraySlice_l183_22;
  wire                when_ArraySlice_l182_23;
  wire                when_ArraySlice_l183_23;
  wire                when_ArraySlice_l361;
  wire                when_ArraySlice_l364;
  wire                when_ArraySlice_l364_1;
  wire                when_ArraySlice_l364_2;
  wire                when_ArraySlice_l364_3;
  wire                when_ArraySlice_l364_4;
  wire                when_ArraySlice_l364_5;
  wire                when_ArraySlice_l364_6;
  wire                when_ArraySlice_l364_7;
  `ifndef SYNTHESIS
  reg [103:0] arraySliceStateMachine_stateReg_string;
  reg [103:0] arraySliceStateMachine_stateNext_string;
  `endif


  assign _zz_handshakeTimes_0_valueNext_1 = handshakeTimes_0_willIncrement;
  assign _zz_handshakeTimes_0_valueNext = {12'd0, _zz_handshakeTimes_0_valueNext_1};
  assign _zz_handshakeTimes_1_valueNext_1 = handshakeTimes_1_willIncrement;
  assign _zz_handshakeTimes_1_valueNext = {12'd0, _zz_handshakeTimes_1_valueNext_1};
  assign _zz_handshakeTimes_2_valueNext_1 = handshakeTimes_2_willIncrement;
  assign _zz_handshakeTimes_2_valueNext = {12'd0, _zz_handshakeTimes_2_valueNext_1};
  assign _zz_handshakeTimes_3_valueNext_1 = handshakeTimes_3_willIncrement;
  assign _zz_handshakeTimes_3_valueNext = {12'd0, _zz_handshakeTimes_3_valueNext_1};
  assign _zz_handshakeTimes_4_valueNext_1 = handshakeTimes_4_willIncrement;
  assign _zz_handshakeTimes_4_valueNext = {12'd0, _zz_handshakeTimes_4_valueNext_1};
  assign _zz_handshakeTimes_5_valueNext_1 = handshakeTimes_5_willIncrement;
  assign _zz_handshakeTimes_5_valueNext = {12'd0, _zz_handshakeTimes_5_valueNext_1};
  assign _zz_handshakeTimes_6_valueNext_1 = handshakeTimes_6_willIncrement;
  assign _zz_handshakeTimes_6_valueNext = {12'd0, _zz_handshakeTimes_6_valueNext_1};
  assign _zz_handshakeTimes_7_valueNext_1 = handshakeTimes_7_willIncrement;
  assign _zz_handshakeTimes_7_valueNext = {12'd0, _zz_handshakeTimes_7_valueNext_1};
  assign _zz_outSliceNumb_0_valueNext_1 = outSliceNumb_0_willIncrement;
  assign _zz_outSliceNumb_0_valueNext = {6'd0, _zz_outSliceNumb_0_valueNext_1};
  assign _zz_outSliceNumb_1_valueNext_1 = outSliceNumb_1_willIncrement;
  assign _zz_outSliceNumb_1_valueNext = {6'd0, _zz_outSliceNumb_1_valueNext_1};
  assign _zz_outSliceNumb_2_valueNext_1 = outSliceNumb_2_willIncrement;
  assign _zz_outSliceNumb_2_valueNext = {6'd0, _zz_outSliceNumb_2_valueNext_1};
  assign _zz_outSliceNumb_3_valueNext_1 = outSliceNumb_3_willIncrement;
  assign _zz_outSliceNumb_3_valueNext = {6'd0, _zz_outSliceNumb_3_valueNext_1};
  assign _zz_outSliceNumb_4_valueNext_1 = outSliceNumb_4_willIncrement;
  assign _zz_outSliceNumb_4_valueNext = {6'd0, _zz_outSliceNumb_4_valueNext_1};
  assign _zz_outSliceNumb_5_valueNext_1 = outSliceNumb_5_willIncrement;
  assign _zz_outSliceNumb_5_valueNext = {6'd0, _zz_outSliceNumb_5_valueNext_1};
  assign _zz_outSliceNumb_6_valueNext_1 = outSliceNumb_6_willIncrement;
  assign _zz_outSliceNumb_6_valueNext = {6'd0, _zz_outSliceNumb_6_valueNext_1};
  assign _zz_outSliceNumb_7_valueNext_1 = outSliceNumb_7_willIncrement;
  assign _zz_outSliceNumb_7_valueNext = {6'd0, _zz_outSliceNumb_7_valueNext_1};
  assign _zz_when_ArraySlice_l208_1 = (hReg - 7'h01);
  assign _zz_when_ArraySlice_l209 = (wReg - 7'h01);
  assign _zz_when_ArraySlice_l158 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_1);
  assign _zz_when_ArraySlice_l158_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_1 = {4'd0, _zz_when_ArraySlice_l158_2};
  assign _zz_when_ArraySlice_l158_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_1 = (_zz_when_ArraySlice_l159_2 - _zz_when_ArraySlice_l159_3);
  assign _zz_when_ArraySlice_l159_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_4);
  assign _zz_when_ArraySlice_l159_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_4 = {4'd0, _zz_when_ArraySlice_l159_5};
  assign _zz__zz_realValue_0 = {1'd0, wReg};
  assign _zz__zz_realValue_0_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_416 = (_zz_realValue_0_417 + _zz_realValue_0_418);
  assign _zz_realValue_0_417 = {1'd0, wReg};
  assign _zz_realValue_0_418 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_1 = (_zz_when_ArraySlice_l166_2 + _zz_when_ArraySlice_l166_6);
  assign _zz_when_ArraySlice_l166_2 = (realValue_0 - _zz_when_ArraySlice_l166_3);
  assign _zz_when_ArraySlice_l166_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_4);
  assign _zz_when_ArraySlice_l166_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_4 = {4'd0, _zz_when_ArraySlice_l166_5};
  assign _zz_when_ArraySlice_l166_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_1_2);
  assign _zz_when_ArraySlice_l158_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_1_2 = {3'd0, _zz_when_ArraySlice_l158_1_3};
  assign _zz_when_ArraySlice_l158_1_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_1_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_1_1 = {1'd0, _zz_when_ArraySlice_l159_1_2};
  assign _zz_when_ArraySlice_l159_1_3 = (_zz_when_ArraySlice_l159_1_4 - _zz_when_ArraySlice_l159_1_5);
  assign _zz_when_ArraySlice_l159_1_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_1_5 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_1_6);
  assign _zz_when_ArraySlice_l159_1_7 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_1_6 = {3'd0, _zz_when_ArraySlice_l159_1_7};
  assign _zz__zz_realValue_0_1_1 = {1'd0, wReg};
  assign _zz__zz_realValue_0_1_2 = (bReg * 4'b1000);
  assign _zz_realValue_0_1_1 = (_zz_realValue_0_1_2 + _zz_realValue_0_1_3);
  assign _zz_realValue_0_1_2 = {1'd0, wReg};
  assign _zz_realValue_0_1_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_1_2 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_1_1 = {1'd0, _zz_when_ArraySlice_l166_1_2};
  assign _zz_when_ArraySlice_l166_1_3 = (_zz_when_ArraySlice_l166_1_4 + _zz_when_ArraySlice_l166_1_8);
  assign _zz_when_ArraySlice_l166_1_4 = (realValue_0_1 - _zz_when_ArraySlice_l166_1_5);
  assign _zz_when_ArraySlice_l166_1_5 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_1_6);
  assign _zz_when_ArraySlice_l166_1_7 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_1_6 = {3'd0, _zz_when_ArraySlice_l166_1_7};
  assign _zz_when_ArraySlice_l166_1_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_2_2);
  assign _zz_when_ArraySlice_l158_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_2_2 = {2'd0, _zz_when_ArraySlice_l158_2_3};
  assign _zz_when_ArraySlice_l158_2_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_2_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_2_1 = {1'd0, _zz_when_ArraySlice_l159_2_2};
  assign _zz_when_ArraySlice_l159_2_3 = (_zz_when_ArraySlice_l159_2_4 - _zz_when_ArraySlice_l159_2_5);
  assign _zz_when_ArraySlice_l159_2_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_2_5 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_2_6);
  assign _zz_when_ArraySlice_l159_2_7 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_2_6 = {2'd0, _zz_when_ArraySlice_l159_2_7};
  assign _zz__zz_realValue_0_2 = {1'd0, wReg};
  assign _zz__zz_realValue_0_2_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_2_1 = (_zz_realValue_0_2_2 + _zz_realValue_0_2_3);
  assign _zz_realValue_0_2_2 = {1'd0, wReg};
  assign _zz_realValue_0_2_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_2_2 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_2_1 = {1'd0, _zz_when_ArraySlice_l166_2_2};
  assign _zz_when_ArraySlice_l166_2_3 = (_zz_when_ArraySlice_l166_2_4 + _zz_when_ArraySlice_l166_2_8);
  assign _zz_when_ArraySlice_l166_2_4 = (realValue_0_2 - _zz_when_ArraySlice_l166_2_5);
  assign _zz_when_ArraySlice_l166_2_5 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_2_6);
  assign _zz_when_ArraySlice_l166_2_7 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_2_6 = {2'd0, _zz_when_ArraySlice_l166_2_7};
  assign _zz_when_ArraySlice_l166_2_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_3_1 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_3_2);
  assign _zz_when_ArraySlice_l158_3_3 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_3_2 = {2'd0, _zz_when_ArraySlice_l158_3_3};
  assign _zz_when_ArraySlice_l158_3_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_3_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_3_1 = {1'd0, _zz_when_ArraySlice_l159_3_2};
  assign _zz_when_ArraySlice_l159_3_3 = (_zz_when_ArraySlice_l159_3_4 - _zz_when_ArraySlice_l159_3_5);
  assign _zz_when_ArraySlice_l159_3_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_3_5 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_3_6);
  assign _zz_when_ArraySlice_l159_3_7 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_3_6 = {2'd0, _zz_when_ArraySlice_l159_3_7};
  assign _zz__zz_realValue_0_3 = {1'd0, wReg};
  assign _zz__zz_realValue_0_3_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_3_1 = (_zz_realValue_0_3_2 + _zz_realValue_0_3_3);
  assign _zz_realValue_0_3_2 = {1'd0, wReg};
  assign _zz_realValue_0_3_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_3_2 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_3_1 = {1'd0, _zz_when_ArraySlice_l166_3_2};
  assign _zz_when_ArraySlice_l166_3_3 = (_zz_when_ArraySlice_l166_3_4 + _zz_when_ArraySlice_l166_3_8);
  assign _zz_when_ArraySlice_l166_3_4 = (realValue_0_3 - _zz_when_ArraySlice_l166_3_5);
  assign _zz_when_ArraySlice_l166_3_5 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_3_6);
  assign _zz_when_ArraySlice_l166_3_7 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_3_6 = {2'd0, _zz_when_ArraySlice_l166_3_7};
  assign _zz_when_ArraySlice_l166_3_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_4_1);
  assign _zz_when_ArraySlice_l158_4_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_4_1 = {1'd0, _zz_when_ArraySlice_l158_4_2};
  assign _zz_when_ArraySlice_l158_4_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_4_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_4_1 = {1'd0, _zz_when_ArraySlice_l159_4_2};
  assign _zz_when_ArraySlice_l159_4_3 = (_zz_when_ArraySlice_l159_4_4 - _zz_when_ArraySlice_l159_4_5);
  assign _zz_when_ArraySlice_l159_4_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_4_5 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_4_6);
  assign _zz_when_ArraySlice_l159_4_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_4_6 = {1'd0, _zz_when_ArraySlice_l159_4_7};
  assign _zz__zz_realValue_0_4 = {1'd0, wReg};
  assign _zz__zz_realValue_0_4_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_4_1 = (_zz_realValue_0_4_2 + _zz_realValue_0_4_3);
  assign _zz_realValue_0_4_2 = {1'd0, wReg};
  assign _zz_realValue_0_4_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_4_2 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_4_1 = {1'd0, _zz_when_ArraySlice_l166_4_2};
  assign _zz_when_ArraySlice_l166_4_3 = (_zz_when_ArraySlice_l166_4_4 + _zz_when_ArraySlice_l166_4_8);
  assign _zz_when_ArraySlice_l166_4_4 = (realValue_0_4 - _zz_when_ArraySlice_l166_4_5);
  assign _zz_when_ArraySlice_l166_4_5 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_4_6);
  assign _zz_when_ArraySlice_l166_4_7 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_4_6 = {1'd0, _zz_when_ArraySlice_l166_4_7};
  assign _zz_when_ArraySlice_l166_4_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_5_1);
  assign _zz_when_ArraySlice_l158_5_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_5_1 = {1'd0, _zz_when_ArraySlice_l158_5_2};
  assign _zz_when_ArraySlice_l158_5_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_5_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_5_1 = {2'd0, _zz_when_ArraySlice_l159_5_2};
  assign _zz_when_ArraySlice_l159_5_3 = (_zz_when_ArraySlice_l159_5_4 - _zz_when_ArraySlice_l159_5_5);
  assign _zz_when_ArraySlice_l159_5_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_5_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_5_6);
  assign _zz_when_ArraySlice_l159_5_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_5_6 = {1'd0, _zz_when_ArraySlice_l159_5_7};
  assign _zz__zz_realValue_0_5 = {1'd0, wReg};
  assign _zz__zz_realValue_0_5_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_5_1 = (_zz_realValue_0_5_2 + _zz_realValue_0_5_3);
  assign _zz_realValue_0_5_2 = {1'd0, wReg};
  assign _zz_realValue_0_5_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_5_2 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_5_1 = {2'd0, _zz_when_ArraySlice_l166_5_2};
  assign _zz_when_ArraySlice_l166_5_3 = (_zz_when_ArraySlice_l166_5_4 + _zz_when_ArraySlice_l166_5_8);
  assign _zz_when_ArraySlice_l166_5_4 = (realValue_0_5 - _zz_when_ArraySlice_l166_5_5);
  assign _zz_when_ArraySlice_l166_5_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_5_6);
  assign _zz_when_ArraySlice_l166_5_7 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_5_6 = {1'd0, _zz_when_ArraySlice_l166_5_7};
  assign _zz_when_ArraySlice_l166_5_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_6_1);
  assign _zz_when_ArraySlice_l158_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_6_1 = {1'd0, _zz_when_ArraySlice_l158_6_2};
  assign _zz_when_ArraySlice_l158_6_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_6_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_6 = {2'd0, _zz_when_ArraySlice_l159_6_1};
  assign _zz_when_ArraySlice_l159_6_2 = (_zz_when_ArraySlice_l159_6_3 - _zz_when_ArraySlice_l159_6_4);
  assign _zz_when_ArraySlice_l159_6_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_6_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_6_5);
  assign _zz_when_ArraySlice_l159_6_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_6_5 = {1'd0, _zz_when_ArraySlice_l159_6_6};
  assign _zz__zz_realValue_0_6 = {1'd0, wReg};
  assign _zz__zz_realValue_0_6_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_6_1 = (_zz_realValue_0_6_2 + _zz_realValue_0_6_3);
  assign _zz_realValue_0_6_2 = {1'd0, wReg};
  assign _zz_realValue_0_6_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_6_2 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_6_1 = {2'd0, _zz_when_ArraySlice_l166_6_2};
  assign _zz_when_ArraySlice_l166_6_3 = (_zz_when_ArraySlice_l166_6_4 + _zz_when_ArraySlice_l166_6_8);
  assign _zz_when_ArraySlice_l166_6_4 = (realValue_0_6 - _zz_when_ArraySlice_l166_6_5);
  assign _zz_when_ArraySlice_l166_6_5 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_6_6);
  assign _zz_when_ArraySlice_l166_6_7 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_6_6 = {1'd0, _zz_when_ArraySlice_l166_6_7};
  assign _zz_when_ArraySlice_l166_6_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_7_1);
  assign _zz_when_ArraySlice_l158_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_7_1 = {1'd0, _zz_when_ArraySlice_l158_7_2};
  assign _zz_when_ArraySlice_l158_7_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_7_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_7 = {3'd0, _zz_when_ArraySlice_l159_7_1};
  assign _zz_when_ArraySlice_l159_7_2 = (_zz_when_ArraySlice_l159_7_3 - _zz_when_ArraySlice_l159_7_4);
  assign _zz_when_ArraySlice_l159_7_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_7_5);
  assign _zz_when_ArraySlice_l159_7_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_7_5 = {1'd0, _zz_when_ArraySlice_l159_7_6};
  assign _zz__zz_realValue_0_7 = {1'd0, wReg};
  assign _zz__zz_realValue_0_7_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_7_1 = (_zz_realValue_0_7_2 + _zz_realValue_0_7_3);
  assign _zz_realValue_0_7_2 = {1'd0, wReg};
  assign _zz_realValue_0_7_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_7_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_7 = {3'd0, _zz_when_ArraySlice_l166_7_1};
  assign _zz_when_ArraySlice_l166_7_2 = (_zz_when_ArraySlice_l166_7_3 + _zz_when_ArraySlice_l166_7_7);
  assign _zz_when_ArraySlice_l166_7_3 = (realValue_0_7 - _zz_when_ArraySlice_l166_7_4);
  assign _zz_when_ArraySlice_l166_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_7_5);
  assign _zz_when_ArraySlice_l166_7_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_7_5 = {1'd0, _zz_when_ArraySlice_l166_7_6};
  assign _zz_when_ArraySlice_l166_7_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l376 = (selectReadFifo_0 + _zz_when_ArraySlice_l376_1);
  assign _zz_when_ArraySlice_l376_2 = 4'b0000;
  assign _zz_when_ArraySlice_l376_1 = {4'd0, _zz_when_ArraySlice_l376_2};
  assign _zz_when_ArraySlice_l376_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l377_3);
  assign _zz_when_ArraySlice_l377_1 = _zz_when_ArraySlice_l377_2[6:0];
  assign _zz_when_ArraySlice_l377_4 = 4'b0000;
  assign _zz_when_ArraySlice_l377_3 = {4'd0, _zz_when_ArraySlice_l377_4};
  assign _zz__zz_outputStreamArrayData_0_valid_1 = 4'b0000;
  assign _zz__zz_outputStreamArrayData_0_valid = {4'd0, _zz__zz_outputStreamArrayData_0_valid_1};
  assign _zz__zz_3 = _zz_outputStreamArrayData_0_valid[6:0];
  assign _zz_outputStreamArrayData_0_valid_3 = _zz_outputStreamArrayData_0_valid[6:0];
  assign _zz_outputStreamArrayData_0_payload_1 = _zz_outputStreamArrayData_0_valid[6:0];
  assign _zz_when_ArraySlice_l383_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l383_3);
  assign _zz_when_ArraySlice_l383_1 = _zz_when_ArraySlice_l383_2[6:0];
  assign _zz_when_ArraySlice_l383_4 = 4'b0000;
  assign _zz_when_ArraySlice_l383_3 = {4'd0, _zz_when_ArraySlice_l383_4};
  assign _zz_when_ArraySlice_l384_1 = (_zz_when_ArraySlice_l384_2 - 8'h01);
  assign _zz_when_ArraySlice_l384 = {5'd0, _zz_when_ArraySlice_l384_1};
  assign _zz_when_ArraySlice_l384_2 = (bReg * aReg);
  assign _zz_selectReadFifo_0 = (selectReadFifo_0 - _zz_selectReadFifo_0_1);
  assign _zz_selectReadFifo_0_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387 = (_zz_when_ArraySlice_l387_1 % aReg);
  assign _zz_when_ArraySlice_l387_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l392_3);
  assign _zz_when_ArraySlice_l392_1 = _zz_when_ArraySlice_l392_2[6:0];
  assign _zz_when_ArraySlice_l392_4 = 4'b0000;
  assign _zz_when_ArraySlice_l392_3 = {4'd0, _zz_when_ArraySlice_l392_4};
  assign _zz_when_ArraySlice_l393_1 = (_zz_when_ArraySlice_l393_2 - 8'h01);
  assign _zz_when_ArraySlice_l393 = {5'd0, _zz_when_ArraySlice_l393_1};
  assign _zz_when_ArraySlice_l393_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_48 = (_zz_realValue1_0_49 + _zz_realValue1_0_50);
  assign _zz_realValue1_0_49 = {1'd0, hReg};
  assign _zz_realValue1_0_50 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l395 = {1'd0, _zz_when_ArraySlice_l395_1};
  assign _zz_when_ArraySlice_l395_2 = (realValue1_0 / aReg);
  assign _zz_selectReadFifo_0_2 = (selectReadFifo_0 - _zz_selectReadFifo_0_3);
  assign _zz_selectReadFifo_0_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_0_5 = 1'b1;
  assign _zz_selectReadFifo_0_4 = {7'd0, _zz_selectReadFifo_0_5};
  assign _zz_when_ArraySlice_l158_8 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_8_1);
  assign _zz_when_ArraySlice_l158_8_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_8_1 = {4'd0, _zz_when_ArraySlice_l158_8_2};
  assign _zz_when_ArraySlice_l158_8_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_8 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_8_1 = (_zz_when_ArraySlice_l159_8_2 - _zz_when_ArraySlice_l159_8_3);
  assign _zz_when_ArraySlice_l159_8_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_8_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_8_4);
  assign _zz_when_ArraySlice_l159_8_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_8_4 = {4'd0, _zz_when_ArraySlice_l159_8_5};
  assign _zz__zz_realValue_0_8 = {1'd0, wReg};
  assign _zz__zz_realValue_0_8_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_8_1 = (_zz_realValue_0_8_2 + _zz_realValue_0_8_3);
  assign _zz_realValue_0_8_2 = {1'd0, wReg};
  assign _zz_realValue_0_8_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_8 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_8_1 = (_zz_when_ArraySlice_l166_8_2 + _zz_when_ArraySlice_l166_8_6);
  assign _zz_when_ArraySlice_l166_8_2 = (realValue_0_8 - _zz_when_ArraySlice_l166_8_3);
  assign _zz_when_ArraySlice_l166_8_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_8_4);
  assign _zz_when_ArraySlice_l166_8_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_8_4 = {4'd0, _zz_when_ArraySlice_l166_8_5};
  assign _zz_when_ArraySlice_l166_8_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_9 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_9_1);
  assign _zz_when_ArraySlice_l158_9_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_9_1 = {3'd0, _zz_when_ArraySlice_l158_9_2};
  assign _zz_when_ArraySlice_l158_9_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_9_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_9 = {1'd0, _zz_when_ArraySlice_l159_9_1};
  assign _zz_when_ArraySlice_l159_9_2 = (_zz_when_ArraySlice_l159_9_3 - _zz_when_ArraySlice_l159_9_4);
  assign _zz_when_ArraySlice_l159_9_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_9_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_9_5);
  assign _zz_when_ArraySlice_l159_9_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_9_5 = {3'd0, _zz_when_ArraySlice_l159_9_6};
  assign _zz__zz_realValue_0_9 = {1'd0, wReg};
  assign _zz__zz_realValue_0_9_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_9_1 = (_zz_realValue_0_9_2 + _zz_realValue_0_9_3);
  assign _zz_realValue_0_9_2 = {1'd0, wReg};
  assign _zz_realValue_0_9_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_9_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_9 = {1'd0, _zz_when_ArraySlice_l166_9_1};
  assign _zz_when_ArraySlice_l166_9_2 = (_zz_when_ArraySlice_l166_9_3 + _zz_when_ArraySlice_l166_9_7);
  assign _zz_when_ArraySlice_l166_9_3 = (realValue_0_9 - _zz_when_ArraySlice_l166_9_4);
  assign _zz_when_ArraySlice_l166_9_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_9_5);
  assign _zz_when_ArraySlice_l166_9_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_9_5 = {3'd0, _zz_when_ArraySlice_l166_9_6};
  assign _zz_when_ArraySlice_l166_9_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_10 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_10_1);
  assign _zz_when_ArraySlice_l158_10_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_10_1 = {2'd0, _zz_when_ArraySlice_l158_10_2};
  assign _zz_when_ArraySlice_l158_10_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_10_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_10 = {1'd0, _zz_when_ArraySlice_l159_10_1};
  assign _zz_when_ArraySlice_l159_10_2 = (_zz_when_ArraySlice_l159_10_3 - _zz_when_ArraySlice_l159_10_4);
  assign _zz_when_ArraySlice_l159_10_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_10_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_10_5);
  assign _zz_when_ArraySlice_l159_10_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_10_5 = {2'd0, _zz_when_ArraySlice_l159_10_6};
  assign _zz__zz_realValue_0_10 = {1'd0, wReg};
  assign _zz__zz_realValue_0_10_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_10_1 = (_zz_realValue_0_10_2 + _zz_realValue_0_10_3);
  assign _zz_realValue_0_10_2 = {1'd0, wReg};
  assign _zz_realValue_0_10_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_10_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_10 = {1'd0, _zz_when_ArraySlice_l166_10_1};
  assign _zz_when_ArraySlice_l166_10_2 = (_zz_when_ArraySlice_l166_10_3 + _zz_when_ArraySlice_l166_10_7);
  assign _zz_when_ArraySlice_l166_10_3 = (realValue_0_10 - _zz_when_ArraySlice_l166_10_4);
  assign _zz_when_ArraySlice_l166_10_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_10_5);
  assign _zz_when_ArraySlice_l166_10_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_10_5 = {2'd0, _zz_when_ArraySlice_l166_10_6};
  assign _zz_when_ArraySlice_l166_10_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_11 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_11_1);
  assign _zz_when_ArraySlice_l158_11_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_11_1 = {2'd0, _zz_when_ArraySlice_l158_11_2};
  assign _zz_when_ArraySlice_l158_11_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_11_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_11 = {1'd0, _zz_when_ArraySlice_l159_11_1};
  assign _zz_when_ArraySlice_l159_11_2 = (_zz_when_ArraySlice_l159_11_3 - _zz_when_ArraySlice_l159_11_4);
  assign _zz_when_ArraySlice_l159_11_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_11_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_11_5);
  assign _zz_when_ArraySlice_l159_11_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_11_5 = {2'd0, _zz_when_ArraySlice_l159_11_6};
  assign _zz__zz_realValue_0_11 = {1'd0, wReg};
  assign _zz__zz_realValue_0_11_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_11_1 = (_zz_realValue_0_11_2 + _zz_realValue_0_11_3);
  assign _zz_realValue_0_11_2 = {1'd0, wReg};
  assign _zz_realValue_0_11_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_11_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_11 = {1'd0, _zz_when_ArraySlice_l166_11_1};
  assign _zz_when_ArraySlice_l166_11_2 = (_zz_when_ArraySlice_l166_11_3 + _zz_when_ArraySlice_l166_11_7);
  assign _zz_when_ArraySlice_l166_11_3 = (realValue_0_11 - _zz_when_ArraySlice_l166_11_4);
  assign _zz_when_ArraySlice_l166_11_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_11_5);
  assign _zz_when_ArraySlice_l166_11_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_11_5 = {2'd0, _zz_when_ArraySlice_l166_11_6};
  assign _zz_when_ArraySlice_l166_11_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_12 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_12_1);
  assign _zz_when_ArraySlice_l158_12_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_12_1 = {1'd0, _zz_when_ArraySlice_l158_12_2};
  assign _zz_when_ArraySlice_l158_12_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_12_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_12 = {1'd0, _zz_when_ArraySlice_l159_12_1};
  assign _zz_when_ArraySlice_l159_12_2 = (_zz_when_ArraySlice_l159_12_3 - _zz_when_ArraySlice_l159_12_4);
  assign _zz_when_ArraySlice_l159_12_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_12_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_12_5);
  assign _zz_when_ArraySlice_l159_12_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_12_5 = {1'd0, _zz_when_ArraySlice_l159_12_6};
  assign _zz__zz_realValue_0_12 = {1'd0, wReg};
  assign _zz__zz_realValue_0_12_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_12_1 = (_zz_realValue_0_12_2 + _zz_realValue_0_12_3);
  assign _zz_realValue_0_12_2 = {1'd0, wReg};
  assign _zz_realValue_0_12_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_12_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_12 = {1'd0, _zz_when_ArraySlice_l166_12_1};
  assign _zz_when_ArraySlice_l166_12_2 = (_zz_when_ArraySlice_l166_12_3 + _zz_when_ArraySlice_l166_12_7);
  assign _zz_when_ArraySlice_l166_12_3 = (realValue_0_12 - _zz_when_ArraySlice_l166_12_4);
  assign _zz_when_ArraySlice_l166_12_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_12_5);
  assign _zz_when_ArraySlice_l166_12_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_12_5 = {1'd0, _zz_when_ArraySlice_l166_12_6};
  assign _zz_when_ArraySlice_l166_12_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_13 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_13_1);
  assign _zz_when_ArraySlice_l158_13_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_13_1 = {1'd0, _zz_when_ArraySlice_l158_13_2};
  assign _zz_when_ArraySlice_l158_13_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_13_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_13 = {2'd0, _zz_when_ArraySlice_l159_13_1};
  assign _zz_when_ArraySlice_l159_13_2 = (_zz_when_ArraySlice_l159_13_3 - _zz_when_ArraySlice_l159_13_4);
  assign _zz_when_ArraySlice_l159_13_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_13_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_13_5);
  assign _zz_when_ArraySlice_l159_13_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_13_5 = {1'd0, _zz_when_ArraySlice_l159_13_6};
  assign _zz__zz_realValue_0_13 = {1'd0, wReg};
  assign _zz__zz_realValue_0_13_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_13_1 = (_zz_realValue_0_13_2 + _zz_realValue_0_13_3);
  assign _zz_realValue_0_13_2 = {1'd0, wReg};
  assign _zz_realValue_0_13_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_13_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_13 = {2'd0, _zz_when_ArraySlice_l166_13_1};
  assign _zz_when_ArraySlice_l166_13_2 = (_zz_when_ArraySlice_l166_13_3 + _zz_when_ArraySlice_l166_13_7);
  assign _zz_when_ArraySlice_l166_13_3 = (realValue_0_13 - _zz_when_ArraySlice_l166_13_4);
  assign _zz_when_ArraySlice_l166_13_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_13_5);
  assign _zz_when_ArraySlice_l166_13_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_13_5 = {1'd0, _zz_when_ArraySlice_l166_13_6};
  assign _zz_when_ArraySlice_l166_13_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_14 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_14_1);
  assign _zz_when_ArraySlice_l158_14_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_14_1 = {1'd0, _zz_when_ArraySlice_l158_14_2};
  assign _zz_when_ArraySlice_l158_14_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_14_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_14 = {2'd0, _zz_when_ArraySlice_l159_14_1};
  assign _zz_when_ArraySlice_l159_14_2 = (_zz_when_ArraySlice_l159_14_3 - _zz_when_ArraySlice_l159_14_4);
  assign _zz_when_ArraySlice_l159_14_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_14_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_14_5);
  assign _zz_when_ArraySlice_l159_14_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_14_5 = {1'd0, _zz_when_ArraySlice_l159_14_6};
  assign _zz__zz_realValue_0_14 = {1'd0, wReg};
  assign _zz__zz_realValue_0_14_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_14_1 = (_zz_realValue_0_14_2 + _zz_realValue_0_14_3);
  assign _zz_realValue_0_14_2 = {1'd0, wReg};
  assign _zz_realValue_0_14_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_14_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_14 = {2'd0, _zz_when_ArraySlice_l166_14_1};
  assign _zz_when_ArraySlice_l166_14_2 = (_zz_when_ArraySlice_l166_14_3 + _zz_when_ArraySlice_l166_14_7);
  assign _zz_when_ArraySlice_l166_14_3 = (realValue_0_14 - _zz_when_ArraySlice_l166_14_4);
  assign _zz_when_ArraySlice_l166_14_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_14_5);
  assign _zz_when_ArraySlice_l166_14_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_14_5 = {1'd0, _zz_when_ArraySlice_l166_14_6};
  assign _zz_when_ArraySlice_l166_14_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_15 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_15_1);
  assign _zz_when_ArraySlice_l158_15_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_15_1 = {1'd0, _zz_when_ArraySlice_l158_15_2};
  assign _zz_when_ArraySlice_l158_15_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_15_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_15 = {3'd0, _zz_when_ArraySlice_l159_15_1};
  assign _zz_when_ArraySlice_l159_15_2 = (_zz_when_ArraySlice_l159_15_3 - _zz_when_ArraySlice_l159_15_4);
  assign _zz_when_ArraySlice_l159_15_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_15_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_15_5);
  assign _zz_when_ArraySlice_l159_15_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_15_5 = {1'd0, _zz_when_ArraySlice_l159_15_6};
  assign _zz__zz_realValue_0_15 = {1'd0, wReg};
  assign _zz__zz_realValue_0_15_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_15_1 = (_zz_realValue_0_15_2 + _zz_realValue_0_15_3);
  assign _zz_realValue_0_15_2 = {1'd0, wReg};
  assign _zz_realValue_0_15_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_15_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_15 = {3'd0, _zz_when_ArraySlice_l166_15_1};
  assign _zz_when_ArraySlice_l166_15_2 = (_zz_when_ArraySlice_l166_15_3 + _zz_when_ArraySlice_l166_15_7);
  assign _zz_when_ArraySlice_l166_15_3 = (realValue_0_15 - _zz_when_ArraySlice_l166_15_4);
  assign _zz_when_ArraySlice_l166_15_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_15_5);
  assign _zz_when_ArraySlice_l166_15_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_15_5 = {1'd0, _zz_when_ArraySlice_l166_15_6};
  assign _zz_when_ArraySlice_l166_15_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_1 = (_zz_when_ArraySlice_l403_2 + _zz_when_ArraySlice_l403_6);
  assign _zz_when_ArraySlice_l403_2 = (_zz_when_ArraySlice_l403_3 + 8'h01);
  assign _zz_when_ArraySlice_l403_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l403_4);
  assign _zz_when_ArraySlice_l403_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_4 = {1'd0, _zz_when_ArraySlice_l403_5};
  assign _zz_when_ArraySlice_l403_7 = 4'b0000;
  assign _zz_when_ArraySlice_l403_6 = {4'd0, _zz_when_ArraySlice_l403_7};
  assign _zz_when_ArraySlice_l406 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_1 = (_zz_when_ArraySlice_l406_2 + 8'h01);
  assign _zz_when_ArraySlice_l406_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l406_3);
  assign _zz_when_ArraySlice_l406_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_3 = {1'd0, _zz_when_ArraySlice_l406_4};
  assign _zz_selectReadFifo_0_6 = (selectReadFifo_0 + _zz_selectReadFifo_0_7);
  assign _zz_selectReadFifo_0_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_7 = {1'd0, _zz_selectReadFifo_0_8};
  assign _zz_when_ArraySlice_l413 = (_zz_when_ArraySlice_l413_1 % aReg);
  assign _zz_when_ArraySlice_l413_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l417_3);
  assign _zz_when_ArraySlice_l417_1 = _zz_when_ArraySlice_l417_2[6:0];
  assign _zz_when_ArraySlice_l417_4 = 4'b0000;
  assign _zz_when_ArraySlice_l417_3 = {4'd0, _zz_when_ArraySlice_l417_4};
  assign _zz_when_ArraySlice_l418_1 = (_zz_when_ArraySlice_l418_2 - _zz_when_ArraySlice_l418_3);
  assign _zz_when_ArraySlice_l418 = {5'd0, _zz_when_ArraySlice_l418_1};
  assign _zz_when_ArraySlice_l418_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_4 = 1'b1;
  assign _zz_when_ArraySlice_l418_3 = {7'd0, _zz_when_ArraySlice_l418_4};
  assign _zz__zz_realValue1_0_1_1 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_1_2 = (aReg * 4'b1000);
  assign _zz_realValue1_0_1_1 = (_zz_realValue1_0_1_2 + _zz_realValue1_0_1_3);
  assign _zz_realValue1_0_1_2 = {1'd0, hReg};
  assign _zz_realValue1_0_1_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l420 = {1'd0, _zz_when_ArraySlice_l420_1};
  assign _zz_when_ArraySlice_l420_2 = (realValue1_0_1 / aReg);
  assign _zz_selectReadFifo_0_9 = (selectReadFifo_0 - _zz_selectReadFifo_0_10);
  assign _zz_selectReadFifo_0_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_16 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_16_1);
  assign _zz_when_ArraySlice_l158_16_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_16_1 = {4'd0, _zz_when_ArraySlice_l158_16_2};
  assign _zz_when_ArraySlice_l158_16_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_16 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_16_1 = (_zz_when_ArraySlice_l159_16_2 - _zz_when_ArraySlice_l159_16_3);
  assign _zz_when_ArraySlice_l159_16_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_16_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_16_4);
  assign _zz_when_ArraySlice_l159_16_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_16_4 = {4'd0, _zz_when_ArraySlice_l159_16_5};
  assign _zz__zz_realValue_0_16 = {1'd0, wReg};
  assign _zz__zz_realValue_0_16_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_16_1 = (_zz_realValue_0_16_2 + _zz_realValue_0_16_3);
  assign _zz_realValue_0_16_2 = {1'd0, wReg};
  assign _zz_realValue_0_16_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_16 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_16_1 = (_zz_when_ArraySlice_l166_16_2 + _zz_when_ArraySlice_l166_16_6);
  assign _zz_when_ArraySlice_l166_16_2 = (realValue_0_16 - _zz_when_ArraySlice_l166_16_3);
  assign _zz_when_ArraySlice_l166_16_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_16_4);
  assign _zz_when_ArraySlice_l166_16_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_16_4 = {4'd0, _zz_when_ArraySlice_l166_16_5};
  assign _zz_when_ArraySlice_l166_16_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_17 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_17_1);
  assign _zz_when_ArraySlice_l158_17_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_17_1 = {3'd0, _zz_when_ArraySlice_l158_17_2};
  assign _zz_when_ArraySlice_l158_17_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_17_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_17 = {1'd0, _zz_when_ArraySlice_l159_17_1};
  assign _zz_when_ArraySlice_l159_17_2 = (_zz_when_ArraySlice_l159_17_3 - _zz_when_ArraySlice_l159_17_4);
  assign _zz_when_ArraySlice_l159_17_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_17_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_17_5);
  assign _zz_when_ArraySlice_l159_17_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_17_5 = {3'd0, _zz_when_ArraySlice_l159_17_6};
  assign _zz__zz_realValue_0_17 = {1'd0, wReg};
  assign _zz__zz_realValue_0_17_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_17_1 = (_zz_realValue_0_17_2 + _zz_realValue_0_17_3);
  assign _zz_realValue_0_17_2 = {1'd0, wReg};
  assign _zz_realValue_0_17_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_17_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_17 = {1'd0, _zz_when_ArraySlice_l166_17_1};
  assign _zz_when_ArraySlice_l166_17_2 = (_zz_when_ArraySlice_l166_17_3 + _zz_when_ArraySlice_l166_17_7);
  assign _zz_when_ArraySlice_l166_17_3 = (realValue_0_17 - _zz_when_ArraySlice_l166_17_4);
  assign _zz_when_ArraySlice_l166_17_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_17_5);
  assign _zz_when_ArraySlice_l166_17_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_17_5 = {3'd0, _zz_when_ArraySlice_l166_17_6};
  assign _zz_when_ArraySlice_l166_17_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_18 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_18_1);
  assign _zz_when_ArraySlice_l158_18_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_18_1 = {2'd0, _zz_when_ArraySlice_l158_18_2};
  assign _zz_when_ArraySlice_l158_18_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_18_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_18 = {1'd0, _zz_when_ArraySlice_l159_18_1};
  assign _zz_when_ArraySlice_l159_18_2 = (_zz_when_ArraySlice_l159_18_3 - _zz_when_ArraySlice_l159_18_4);
  assign _zz_when_ArraySlice_l159_18_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_18_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_18_5);
  assign _zz_when_ArraySlice_l159_18_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_18_5 = {2'd0, _zz_when_ArraySlice_l159_18_6};
  assign _zz__zz_realValue_0_18 = {1'd0, wReg};
  assign _zz__zz_realValue_0_18_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_18_1 = (_zz_realValue_0_18_2 + _zz_realValue_0_18_3);
  assign _zz_realValue_0_18_2 = {1'd0, wReg};
  assign _zz_realValue_0_18_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_18_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_18 = {1'd0, _zz_when_ArraySlice_l166_18_1};
  assign _zz_when_ArraySlice_l166_18_2 = (_zz_when_ArraySlice_l166_18_3 + _zz_when_ArraySlice_l166_18_7);
  assign _zz_when_ArraySlice_l166_18_3 = (realValue_0_18 - _zz_when_ArraySlice_l166_18_4);
  assign _zz_when_ArraySlice_l166_18_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_18_5);
  assign _zz_when_ArraySlice_l166_18_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_18_5 = {2'd0, _zz_when_ArraySlice_l166_18_6};
  assign _zz_when_ArraySlice_l166_18_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_19 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_19_1);
  assign _zz_when_ArraySlice_l158_19_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_19_1 = {2'd0, _zz_when_ArraySlice_l158_19_2};
  assign _zz_when_ArraySlice_l158_19_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_19_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_19 = {1'd0, _zz_when_ArraySlice_l159_19_1};
  assign _zz_when_ArraySlice_l159_19_2 = (_zz_when_ArraySlice_l159_19_3 - _zz_when_ArraySlice_l159_19_4);
  assign _zz_when_ArraySlice_l159_19_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_19_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_19_5);
  assign _zz_when_ArraySlice_l159_19_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_19_5 = {2'd0, _zz_when_ArraySlice_l159_19_6};
  assign _zz__zz_realValue_0_19 = {1'd0, wReg};
  assign _zz__zz_realValue_0_19_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_19_1 = (_zz_realValue_0_19_2 + _zz_realValue_0_19_3);
  assign _zz_realValue_0_19_2 = {1'd0, wReg};
  assign _zz_realValue_0_19_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_19_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_19 = {1'd0, _zz_when_ArraySlice_l166_19_1};
  assign _zz_when_ArraySlice_l166_19_2 = (_zz_when_ArraySlice_l166_19_3 + _zz_when_ArraySlice_l166_19_7);
  assign _zz_when_ArraySlice_l166_19_3 = (realValue_0_19 - _zz_when_ArraySlice_l166_19_4);
  assign _zz_when_ArraySlice_l166_19_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_19_5);
  assign _zz_when_ArraySlice_l166_19_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_19_5 = {2'd0, _zz_when_ArraySlice_l166_19_6};
  assign _zz_when_ArraySlice_l166_19_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_20 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_20_1);
  assign _zz_when_ArraySlice_l158_20_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_20_1 = {1'd0, _zz_when_ArraySlice_l158_20_2};
  assign _zz_when_ArraySlice_l158_20_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_20_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_20 = {1'd0, _zz_when_ArraySlice_l159_20_1};
  assign _zz_when_ArraySlice_l159_20_2 = (_zz_when_ArraySlice_l159_20_3 - _zz_when_ArraySlice_l159_20_4);
  assign _zz_when_ArraySlice_l159_20_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_20_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_20_5);
  assign _zz_when_ArraySlice_l159_20_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_20_5 = {1'd0, _zz_when_ArraySlice_l159_20_6};
  assign _zz__zz_realValue_0_20 = {1'd0, wReg};
  assign _zz__zz_realValue_0_20_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_20_1 = (_zz_realValue_0_20_2 + _zz_realValue_0_20_3);
  assign _zz_realValue_0_20_2 = {1'd0, wReg};
  assign _zz_realValue_0_20_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_20_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_20 = {1'd0, _zz_when_ArraySlice_l166_20_1};
  assign _zz_when_ArraySlice_l166_20_2 = (_zz_when_ArraySlice_l166_20_3 + _zz_when_ArraySlice_l166_20_7);
  assign _zz_when_ArraySlice_l166_20_3 = (realValue_0_20 - _zz_when_ArraySlice_l166_20_4);
  assign _zz_when_ArraySlice_l166_20_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_20_5);
  assign _zz_when_ArraySlice_l166_20_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_20_5 = {1'd0, _zz_when_ArraySlice_l166_20_6};
  assign _zz_when_ArraySlice_l166_20_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_21 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_21_1);
  assign _zz_when_ArraySlice_l158_21_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_21_1 = {1'd0, _zz_when_ArraySlice_l158_21_2};
  assign _zz_when_ArraySlice_l158_21_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_21_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_21 = {2'd0, _zz_when_ArraySlice_l159_21_1};
  assign _zz_when_ArraySlice_l159_21_2 = (_zz_when_ArraySlice_l159_21_3 - _zz_when_ArraySlice_l159_21_4);
  assign _zz_when_ArraySlice_l159_21_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_21_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_21_5);
  assign _zz_when_ArraySlice_l159_21_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_21_5 = {1'd0, _zz_when_ArraySlice_l159_21_6};
  assign _zz__zz_realValue_0_21 = {1'd0, wReg};
  assign _zz__zz_realValue_0_21_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_21_1 = (_zz_realValue_0_21_2 + _zz_realValue_0_21_3);
  assign _zz_realValue_0_21_2 = {1'd0, wReg};
  assign _zz_realValue_0_21_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_21_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_21 = {2'd0, _zz_when_ArraySlice_l166_21_1};
  assign _zz_when_ArraySlice_l166_21_2 = (_zz_when_ArraySlice_l166_21_3 + _zz_when_ArraySlice_l166_21_7);
  assign _zz_when_ArraySlice_l166_21_3 = (realValue_0_21 - _zz_when_ArraySlice_l166_21_4);
  assign _zz_when_ArraySlice_l166_21_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_21_5);
  assign _zz_when_ArraySlice_l166_21_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_21_5 = {1'd0, _zz_when_ArraySlice_l166_21_6};
  assign _zz_when_ArraySlice_l166_21_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_22 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_22_1);
  assign _zz_when_ArraySlice_l158_22_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_22_1 = {1'd0, _zz_when_ArraySlice_l158_22_2};
  assign _zz_when_ArraySlice_l158_22_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_22_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_22 = {2'd0, _zz_when_ArraySlice_l159_22_1};
  assign _zz_when_ArraySlice_l159_22_2 = (_zz_when_ArraySlice_l159_22_3 - _zz_when_ArraySlice_l159_22_4);
  assign _zz_when_ArraySlice_l159_22_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_22_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_22_5);
  assign _zz_when_ArraySlice_l159_22_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_22_5 = {1'd0, _zz_when_ArraySlice_l159_22_6};
  assign _zz__zz_realValue_0_22 = {1'd0, wReg};
  assign _zz__zz_realValue_0_22_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_22_1 = (_zz_realValue_0_22_2 + _zz_realValue_0_22_3);
  assign _zz_realValue_0_22_2 = {1'd0, wReg};
  assign _zz_realValue_0_22_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_22_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_22 = {2'd0, _zz_when_ArraySlice_l166_22_1};
  assign _zz_when_ArraySlice_l166_22_2 = (_zz_when_ArraySlice_l166_22_3 + _zz_when_ArraySlice_l166_22_7);
  assign _zz_when_ArraySlice_l166_22_3 = (realValue_0_22 - _zz_when_ArraySlice_l166_22_4);
  assign _zz_when_ArraySlice_l166_22_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_22_5);
  assign _zz_when_ArraySlice_l166_22_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_22_5 = {1'd0, _zz_when_ArraySlice_l166_22_6};
  assign _zz_when_ArraySlice_l166_22_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_23 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_23_1);
  assign _zz_when_ArraySlice_l158_23_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_23_1 = {1'd0, _zz_when_ArraySlice_l158_23_2};
  assign _zz_when_ArraySlice_l158_23_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_23_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_23 = {3'd0, _zz_when_ArraySlice_l159_23_1};
  assign _zz_when_ArraySlice_l159_23_2 = (_zz_when_ArraySlice_l159_23_3 - _zz_when_ArraySlice_l159_23_4);
  assign _zz_when_ArraySlice_l159_23_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_23_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_23_5);
  assign _zz_when_ArraySlice_l159_23_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_23_5 = {1'd0, _zz_when_ArraySlice_l159_23_6};
  assign _zz__zz_realValue_0_23 = {1'd0, wReg};
  assign _zz__zz_realValue_0_23_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_23_1 = (_zz_realValue_0_23_2 + _zz_realValue_0_23_3);
  assign _zz_realValue_0_23_2 = {1'd0, wReg};
  assign _zz_realValue_0_23_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_23_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_23 = {3'd0, _zz_when_ArraySlice_l166_23_1};
  assign _zz_when_ArraySlice_l166_23_2 = (_zz_when_ArraySlice_l166_23_3 + _zz_when_ArraySlice_l166_23_7);
  assign _zz_when_ArraySlice_l166_23_3 = (realValue_0_23 - _zz_when_ArraySlice_l166_23_4);
  assign _zz_when_ArraySlice_l166_23_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_23_5);
  assign _zz_when_ArraySlice_l166_23_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_23_5 = {1'd0, _zz_when_ArraySlice_l166_23_6};
  assign _zz_when_ArraySlice_l166_23_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_1 = (_zz_when_ArraySlice_l428_2 + _zz_when_ArraySlice_l428_6);
  assign _zz_when_ArraySlice_l428_2 = (_zz_when_ArraySlice_l428_3 + 8'h01);
  assign _zz_when_ArraySlice_l428_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l428_4);
  assign _zz_when_ArraySlice_l428_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_4 = {1'd0, _zz_when_ArraySlice_l428_5};
  assign _zz_when_ArraySlice_l428_7 = 4'b0000;
  assign _zz_when_ArraySlice_l428_6 = {4'd0, _zz_when_ArraySlice_l428_7};
  assign _zz_when_ArraySlice_l431 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_1 = (_zz_when_ArraySlice_l431_2 + 8'h01);
  assign _zz_when_ArraySlice_l431_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l431_3);
  assign _zz_when_ArraySlice_l431_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_3 = {1'd0, _zz_when_ArraySlice_l431_4};
  assign _zz_selectReadFifo_0_11 = (selectReadFifo_0 + _zz_selectReadFifo_0_12);
  assign _zz_selectReadFifo_0_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_12 = {1'd0, _zz_selectReadFifo_0_13};
  assign _zz_when_ArraySlice_l438 = (_zz_when_ArraySlice_l438_1 % aReg);
  assign _zz_when_ArraySlice_l438_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_1 = (_zz_when_ArraySlice_l449_2 - 8'h01);
  assign _zz_when_ArraySlice_l449 = {5'd0, _zz_when_ArraySlice_l449_1};
  assign _zz_when_ArraySlice_l449_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_2 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_2_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_2_1 = (_zz_realValue1_0_2_2 + _zz_realValue1_0_2_3);
  assign _zz_realValue1_0_2_2 = {1'd0, hReg};
  assign _zz_realValue1_0_2_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l450 = {1'd0, _zz_when_ArraySlice_l450_1};
  assign _zz_when_ArraySlice_l450_2 = (realValue1_0_2 / aReg);
  assign _zz_selectReadFifo_0_14 = (selectReadFifo_0 - _zz_selectReadFifo_0_15);
  assign _zz_selectReadFifo_0_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_24 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_24_1);
  assign _zz_when_ArraySlice_l158_24_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_24_1 = {4'd0, _zz_when_ArraySlice_l158_24_2};
  assign _zz_when_ArraySlice_l158_24_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_24 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_24_1 = (_zz_when_ArraySlice_l159_24_2 - _zz_when_ArraySlice_l159_24_3);
  assign _zz_when_ArraySlice_l159_24_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_24_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_24_4);
  assign _zz_when_ArraySlice_l159_24_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_24_4 = {4'd0, _zz_when_ArraySlice_l159_24_5};
  assign _zz__zz_realValue_0_24 = {1'd0, wReg};
  assign _zz__zz_realValue_0_24_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_24_1 = (_zz_realValue_0_24_2 + _zz_realValue_0_24_3);
  assign _zz_realValue_0_24_2 = {1'd0, wReg};
  assign _zz_realValue_0_24_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_24 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_24_1 = (_zz_when_ArraySlice_l166_24_2 + _zz_when_ArraySlice_l166_24_6);
  assign _zz_when_ArraySlice_l166_24_2 = (realValue_0_24 - _zz_when_ArraySlice_l166_24_3);
  assign _zz_when_ArraySlice_l166_24_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_24_4);
  assign _zz_when_ArraySlice_l166_24_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_24_4 = {4'd0, _zz_when_ArraySlice_l166_24_5};
  assign _zz_when_ArraySlice_l166_24_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_25 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_25_1);
  assign _zz_when_ArraySlice_l158_25_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_25_1 = {3'd0, _zz_when_ArraySlice_l158_25_2};
  assign _zz_when_ArraySlice_l158_25_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_25_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_25 = {1'd0, _zz_when_ArraySlice_l159_25_1};
  assign _zz_when_ArraySlice_l159_25_2 = (_zz_when_ArraySlice_l159_25_3 - _zz_when_ArraySlice_l159_25_4);
  assign _zz_when_ArraySlice_l159_25_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_25_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_25_5);
  assign _zz_when_ArraySlice_l159_25_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_25_5 = {3'd0, _zz_when_ArraySlice_l159_25_6};
  assign _zz__zz_realValue_0_25 = {1'd0, wReg};
  assign _zz__zz_realValue_0_25_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_25_1 = (_zz_realValue_0_25_2 + _zz_realValue_0_25_3);
  assign _zz_realValue_0_25_2 = {1'd0, wReg};
  assign _zz_realValue_0_25_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_25_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_25 = {1'd0, _zz_when_ArraySlice_l166_25_1};
  assign _zz_when_ArraySlice_l166_25_2 = (_zz_when_ArraySlice_l166_25_3 + _zz_when_ArraySlice_l166_25_7);
  assign _zz_when_ArraySlice_l166_25_3 = (realValue_0_25 - _zz_when_ArraySlice_l166_25_4);
  assign _zz_when_ArraySlice_l166_25_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_25_5);
  assign _zz_when_ArraySlice_l166_25_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_25_5 = {3'd0, _zz_when_ArraySlice_l166_25_6};
  assign _zz_when_ArraySlice_l166_25_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_26 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_26_1);
  assign _zz_when_ArraySlice_l158_26_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_26_1 = {2'd0, _zz_when_ArraySlice_l158_26_2};
  assign _zz_when_ArraySlice_l158_26_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_26_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_26 = {1'd0, _zz_when_ArraySlice_l159_26_1};
  assign _zz_when_ArraySlice_l159_26_2 = (_zz_when_ArraySlice_l159_26_3 - _zz_when_ArraySlice_l159_26_4);
  assign _zz_when_ArraySlice_l159_26_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_26_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_26_5);
  assign _zz_when_ArraySlice_l159_26_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_26_5 = {2'd0, _zz_when_ArraySlice_l159_26_6};
  assign _zz__zz_realValue_0_26 = {1'd0, wReg};
  assign _zz__zz_realValue_0_26_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_26_1 = (_zz_realValue_0_26_2 + _zz_realValue_0_26_3);
  assign _zz_realValue_0_26_2 = {1'd0, wReg};
  assign _zz_realValue_0_26_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_26_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_26 = {1'd0, _zz_when_ArraySlice_l166_26_1};
  assign _zz_when_ArraySlice_l166_26_2 = (_zz_when_ArraySlice_l166_26_3 + _zz_when_ArraySlice_l166_26_7);
  assign _zz_when_ArraySlice_l166_26_3 = (realValue_0_26 - _zz_when_ArraySlice_l166_26_4);
  assign _zz_when_ArraySlice_l166_26_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_26_5);
  assign _zz_when_ArraySlice_l166_26_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_26_5 = {2'd0, _zz_when_ArraySlice_l166_26_6};
  assign _zz_when_ArraySlice_l166_26_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_27 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_27_1);
  assign _zz_when_ArraySlice_l158_27_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_27_1 = {2'd0, _zz_when_ArraySlice_l158_27_2};
  assign _zz_when_ArraySlice_l158_27_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_27_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_27 = {1'd0, _zz_when_ArraySlice_l159_27_1};
  assign _zz_when_ArraySlice_l159_27_2 = (_zz_when_ArraySlice_l159_27_3 - _zz_when_ArraySlice_l159_27_4);
  assign _zz_when_ArraySlice_l159_27_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_27_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_27_5);
  assign _zz_when_ArraySlice_l159_27_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_27_5 = {2'd0, _zz_when_ArraySlice_l159_27_6};
  assign _zz__zz_realValue_0_27 = {1'd0, wReg};
  assign _zz__zz_realValue_0_27_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_27_1 = (_zz_realValue_0_27_2 + _zz_realValue_0_27_3);
  assign _zz_realValue_0_27_2 = {1'd0, wReg};
  assign _zz_realValue_0_27_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_27_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_27 = {1'd0, _zz_when_ArraySlice_l166_27_1};
  assign _zz_when_ArraySlice_l166_27_2 = (_zz_when_ArraySlice_l166_27_3 + _zz_when_ArraySlice_l166_27_7);
  assign _zz_when_ArraySlice_l166_27_3 = (realValue_0_27 - _zz_when_ArraySlice_l166_27_4);
  assign _zz_when_ArraySlice_l166_27_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_27_5);
  assign _zz_when_ArraySlice_l166_27_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_27_5 = {2'd0, _zz_when_ArraySlice_l166_27_6};
  assign _zz_when_ArraySlice_l166_27_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_28 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_28_1);
  assign _zz_when_ArraySlice_l158_28_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_28_1 = {1'd0, _zz_when_ArraySlice_l158_28_2};
  assign _zz_when_ArraySlice_l158_28_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_28_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_28 = {1'd0, _zz_when_ArraySlice_l159_28_1};
  assign _zz_when_ArraySlice_l159_28_2 = (_zz_when_ArraySlice_l159_28_3 - _zz_when_ArraySlice_l159_28_4);
  assign _zz_when_ArraySlice_l159_28_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_28_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_28_5);
  assign _zz_when_ArraySlice_l159_28_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_28_5 = {1'd0, _zz_when_ArraySlice_l159_28_6};
  assign _zz__zz_realValue_0_28 = {1'd0, wReg};
  assign _zz__zz_realValue_0_28_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_28_1 = (_zz_realValue_0_28_2 + _zz_realValue_0_28_3);
  assign _zz_realValue_0_28_2 = {1'd0, wReg};
  assign _zz_realValue_0_28_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_28_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_28 = {1'd0, _zz_when_ArraySlice_l166_28_1};
  assign _zz_when_ArraySlice_l166_28_2 = (_zz_when_ArraySlice_l166_28_3 + _zz_when_ArraySlice_l166_28_7);
  assign _zz_when_ArraySlice_l166_28_3 = (realValue_0_28 - _zz_when_ArraySlice_l166_28_4);
  assign _zz_when_ArraySlice_l166_28_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_28_5);
  assign _zz_when_ArraySlice_l166_28_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_28_5 = {1'd0, _zz_when_ArraySlice_l166_28_6};
  assign _zz_when_ArraySlice_l166_28_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_29 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_29_1);
  assign _zz_when_ArraySlice_l158_29_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_29_1 = {1'd0, _zz_when_ArraySlice_l158_29_2};
  assign _zz_when_ArraySlice_l158_29_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_29_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_29 = {2'd0, _zz_when_ArraySlice_l159_29_1};
  assign _zz_when_ArraySlice_l159_29_2 = (_zz_when_ArraySlice_l159_29_3 - _zz_when_ArraySlice_l159_29_4);
  assign _zz_when_ArraySlice_l159_29_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_29_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_29_5);
  assign _zz_when_ArraySlice_l159_29_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_29_5 = {1'd0, _zz_when_ArraySlice_l159_29_6};
  assign _zz__zz_realValue_0_29 = {1'd0, wReg};
  assign _zz__zz_realValue_0_29_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_29_1 = (_zz_realValue_0_29_2 + _zz_realValue_0_29_3);
  assign _zz_realValue_0_29_2 = {1'd0, wReg};
  assign _zz_realValue_0_29_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_29_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_29 = {2'd0, _zz_when_ArraySlice_l166_29_1};
  assign _zz_when_ArraySlice_l166_29_2 = (_zz_when_ArraySlice_l166_29_3 + _zz_when_ArraySlice_l166_29_7);
  assign _zz_when_ArraySlice_l166_29_3 = (realValue_0_29 - _zz_when_ArraySlice_l166_29_4);
  assign _zz_when_ArraySlice_l166_29_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_29_5);
  assign _zz_when_ArraySlice_l166_29_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_29_5 = {1'd0, _zz_when_ArraySlice_l166_29_6};
  assign _zz_when_ArraySlice_l166_29_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_30 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_30_1);
  assign _zz_when_ArraySlice_l158_30_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_30_1 = {1'd0, _zz_when_ArraySlice_l158_30_2};
  assign _zz_when_ArraySlice_l158_30_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_30_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_30 = {2'd0, _zz_when_ArraySlice_l159_30_1};
  assign _zz_when_ArraySlice_l159_30_2 = (_zz_when_ArraySlice_l159_30_3 - _zz_when_ArraySlice_l159_30_4);
  assign _zz_when_ArraySlice_l159_30_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_30_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_30_5);
  assign _zz_when_ArraySlice_l159_30_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_30_5 = {1'd0, _zz_when_ArraySlice_l159_30_6};
  assign _zz__zz_realValue_0_30 = {1'd0, wReg};
  assign _zz__zz_realValue_0_30_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_30_1 = (_zz_realValue_0_30_2 + _zz_realValue_0_30_3);
  assign _zz_realValue_0_30_2 = {1'd0, wReg};
  assign _zz_realValue_0_30_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_30_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_30 = {2'd0, _zz_when_ArraySlice_l166_30_1};
  assign _zz_when_ArraySlice_l166_30_2 = (_zz_when_ArraySlice_l166_30_3 + _zz_when_ArraySlice_l166_30_7);
  assign _zz_when_ArraySlice_l166_30_3 = (realValue_0_30 - _zz_when_ArraySlice_l166_30_4);
  assign _zz_when_ArraySlice_l166_30_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_30_5);
  assign _zz_when_ArraySlice_l166_30_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_30_5 = {1'd0, _zz_when_ArraySlice_l166_30_6};
  assign _zz_when_ArraySlice_l166_30_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_31 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_31_1);
  assign _zz_when_ArraySlice_l158_31_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_31_1 = {1'd0, _zz_when_ArraySlice_l158_31_2};
  assign _zz_when_ArraySlice_l158_31_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_31_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_31 = {3'd0, _zz_when_ArraySlice_l159_31_1};
  assign _zz_when_ArraySlice_l159_31_2 = (_zz_when_ArraySlice_l159_31_3 - _zz_when_ArraySlice_l159_31_4);
  assign _zz_when_ArraySlice_l159_31_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_31_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_31_5);
  assign _zz_when_ArraySlice_l159_31_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_31_5 = {1'd0, _zz_when_ArraySlice_l159_31_6};
  assign _zz__zz_realValue_0_31 = {1'd0, wReg};
  assign _zz__zz_realValue_0_31_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_31_1 = (_zz_realValue_0_31_2 + _zz_realValue_0_31_3);
  assign _zz_realValue_0_31_2 = {1'd0, wReg};
  assign _zz_realValue_0_31_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_31_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_31 = {3'd0, _zz_when_ArraySlice_l166_31_1};
  assign _zz_when_ArraySlice_l166_31_2 = (_zz_when_ArraySlice_l166_31_3 + _zz_when_ArraySlice_l166_31_7);
  assign _zz_when_ArraySlice_l166_31_3 = (realValue_0_31 - _zz_when_ArraySlice_l166_31_4);
  assign _zz_when_ArraySlice_l166_31_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_31_5);
  assign _zz_when_ArraySlice_l166_31_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_31_5 = {1'd0, _zz_when_ArraySlice_l166_31_6};
  assign _zz_when_ArraySlice_l166_31_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461 = (_zz_when_ArraySlice_l461_1 % aReg);
  assign _zz_when_ArraySlice_l461_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l447 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l447_2);
  assign _zz_when_ArraySlice_l447_3 = 4'b0000;
  assign _zz_when_ArraySlice_l447_2 = {4'd0, _zz_when_ArraySlice_l447_3};
  assign _zz_when_ArraySlice_l468_1 = (_zz_when_ArraySlice_l468_2 - 8'h01);
  assign _zz_when_ArraySlice_l468 = {5'd0, _zz_when_ArraySlice_l468_1};
  assign _zz_when_ArraySlice_l468_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l376_1_2);
  assign _zz_when_ArraySlice_l376_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l376_1_2 = {3'd0, _zz_when_ArraySlice_l376_1_3};
  assign _zz_when_ArraySlice_l376_1_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l377_1_4);
  assign _zz_when_ArraySlice_l377_1_2 = _zz_when_ArraySlice_l377_1_3[6:0];
  assign _zz_when_ArraySlice_l377_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l377_1_4 = {3'd0, _zz_when_ArraySlice_l377_1_5};
  assign _zz__zz_outputStreamArrayData_1_valid_1 = (bReg * 1'b1);
  assign _zz__zz_outputStreamArrayData_1_valid = {3'd0, _zz__zz_outputStreamArrayData_1_valid_1};
  assign _zz__zz_4 = _zz_outputStreamArrayData_1_valid[6:0];
  assign _zz_outputStreamArrayData_1_valid_3 = _zz_outputStreamArrayData_1_valid[6:0];
  assign _zz_outputStreamArrayData_1_payload_1 = _zz_outputStreamArrayData_1_valid[6:0];
  assign _zz_when_ArraySlice_l383_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l383_1_4);
  assign _zz_when_ArraySlice_l383_1_2 = _zz_when_ArraySlice_l383_1_3[6:0];
  assign _zz_when_ArraySlice_l383_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l383_1_4 = {3'd0, _zz_when_ArraySlice_l383_1_5};
  assign _zz_when_ArraySlice_l384_1_2 = (_zz_when_ArraySlice_l384_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l384_1_1 = {5'd0, _zz_when_ArraySlice_l384_1_2};
  assign _zz_when_ArraySlice_l384_1_3 = (bReg * aReg);
  assign _zz_selectReadFifo_1 = (selectReadFifo_1 - _zz_selectReadFifo_1_1);
  assign _zz_selectReadFifo_1_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_1_1 = (_zz_when_ArraySlice_l387_1_2 % aReg);
  assign _zz_when_ArraySlice_l387_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l392_1_4);
  assign _zz_when_ArraySlice_l392_1_2 = _zz_when_ArraySlice_l392_1_3[6:0];
  assign _zz_when_ArraySlice_l392_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l392_1_4 = {3'd0, _zz_when_ArraySlice_l392_1_5};
  assign _zz_when_ArraySlice_l393_1_2 = (_zz_when_ArraySlice_l393_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l393_1_1 = {5'd0, _zz_when_ArraySlice_l393_1_2};
  assign _zz_when_ArraySlice_l393_1_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_3 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_3_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_3_1 = (_zz_realValue1_0_3_2 + _zz_realValue1_0_3_3);
  assign _zz_realValue1_0_3_2 = {1'd0, hReg};
  assign _zz_realValue1_0_3_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l395_1_1 = {1'd0, _zz_when_ArraySlice_l395_1_2};
  assign _zz_when_ArraySlice_l395_1_3 = (realValue1_0_3 / aReg);
  assign _zz_selectReadFifo_1_2 = (selectReadFifo_1 - _zz_selectReadFifo_1_3);
  assign _zz_selectReadFifo_1_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_1_5 = 1'b1;
  assign _zz_selectReadFifo_1_4 = {7'd0, _zz_selectReadFifo_1_5};
  assign _zz_when_ArraySlice_l158_32 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_32_1);
  assign _zz_when_ArraySlice_l158_32_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_32_1 = {4'd0, _zz_when_ArraySlice_l158_32_2};
  assign _zz_when_ArraySlice_l158_32_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_32 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_32_1 = (_zz_when_ArraySlice_l159_32_2 - _zz_when_ArraySlice_l159_32_3);
  assign _zz_when_ArraySlice_l159_32_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_32_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_32_4);
  assign _zz_when_ArraySlice_l159_32_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_32_4 = {4'd0, _zz_when_ArraySlice_l159_32_5};
  assign _zz__zz_realValue_0_32 = {1'd0, wReg};
  assign _zz__zz_realValue_0_32_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_32_1 = (_zz_realValue_0_32_2 + _zz_realValue_0_32_3);
  assign _zz_realValue_0_32_2 = {1'd0, wReg};
  assign _zz_realValue_0_32_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_32 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_32_1 = (_zz_when_ArraySlice_l166_32_2 + _zz_when_ArraySlice_l166_32_6);
  assign _zz_when_ArraySlice_l166_32_2 = (realValue_0_32 - _zz_when_ArraySlice_l166_32_3);
  assign _zz_when_ArraySlice_l166_32_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_32_4);
  assign _zz_when_ArraySlice_l166_32_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_32_4 = {4'd0, _zz_when_ArraySlice_l166_32_5};
  assign _zz_when_ArraySlice_l166_32_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_33 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_33_1);
  assign _zz_when_ArraySlice_l158_33_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_33_1 = {3'd0, _zz_when_ArraySlice_l158_33_2};
  assign _zz_when_ArraySlice_l158_33_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_33_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_33 = {1'd0, _zz_when_ArraySlice_l159_33_1};
  assign _zz_when_ArraySlice_l159_33_2 = (_zz_when_ArraySlice_l159_33_3 - _zz_when_ArraySlice_l159_33_4);
  assign _zz_when_ArraySlice_l159_33_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_33_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_33_5);
  assign _zz_when_ArraySlice_l159_33_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_33_5 = {3'd0, _zz_when_ArraySlice_l159_33_6};
  assign _zz__zz_realValue_0_33 = {1'd0, wReg};
  assign _zz__zz_realValue_0_33_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_33_1 = (_zz_realValue_0_33_2 + _zz_realValue_0_33_3);
  assign _zz_realValue_0_33_2 = {1'd0, wReg};
  assign _zz_realValue_0_33_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_33_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_33 = {1'd0, _zz_when_ArraySlice_l166_33_1};
  assign _zz_when_ArraySlice_l166_33_2 = (_zz_when_ArraySlice_l166_33_3 + _zz_when_ArraySlice_l166_33_7);
  assign _zz_when_ArraySlice_l166_33_3 = (realValue_0_33 - _zz_when_ArraySlice_l166_33_4);
  assign _zz_when_ArraySlice_l166_33_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_33_5);
  assign _zz_when_ArraySlice_l166_33_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_33_5 = {3'd0, _zz_when_ArraySlice_l166_33_6};
  assign _zz_when_ArraySlice_l166_33_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_34 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_34_1);
  assign _zz_when_ArraySlice_l158_34_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_34_1 = {2'd0, _zz_when_ArraySlice_l158_34_2};
  assign _zz_when_ArraySlice_l158_34_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_34_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_34 = {1'd0, _zz_when_ArraySlice_l159_34_1};
  assign _zz_when_ArraySlice_l159_34_2 = (_zz_when_ArraySlice_l159_34_3 - _zz_when_ArraySlice_l159_34_4);
  assign _zz_when_ArraySlice_l159_34_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_34_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_34_5);
  assign _zz_when_ArraySlice_l159_34_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_34_5 = {2'd0, _zz_when_ArraySlice_l159_34_6};
  assign _zz__zz_realValue_0_34 = {1'd0, wReg};
  assign _zz__zz_realValue_0_34_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_34_1 = (_zz_realValue_0_34_2 + _zz_realValue_0_34_3);
  assign _zz_realValue_0_34_2 = {1'd0, wReg};
  assign _zz_realValue_0_34_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_34_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_34 = {1'd0, _zz_when_ArraySlice_l166_34_1};
  assign _zz_when_ArraySlice_l166_34_2 = (_zz_when_ArraySlice_l166_34_3 + _zz_when_ArraySlice_l166_34_7);
  assign _zz_when_ArraySlice_l166_34_3 = (realValue_0_34 - _zz_when_ArraySlice_l166_34_4);
  assign _zz_when_ArraySlice_l166_34_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_34_5);
  assign _zz_when_ArraySlice_l166_34_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_34_5 = {2'd0, _zz_when_ArraySlice_l166_34_6};
  assign _zz_when_ArraySlice_l166_34_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_35 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_35_1);
  assign _zz_when_ArraySlice_l158_35_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_35_1 = {2'd0, _zz_when_ArraySlice_l158_35_2};
  assign _zz_when_ArraySlice_l158_35_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_35_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_35 = {1'd0, _zz_when_ArraySlice_l159_35_1};
  assign _zz_when_ArraySlice_l159_35_2 = (_zz_when_ArraySlice_l159_35_3 - _zz_when_ArraySlice_l159_35_4);
  assign _zz_when_ArraySlice_l159_35_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_35_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_35_5);
  assign _zz_when_ArraySlice_l159_35_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_35_5 = {2'd0, _zz_when_ArraySlice_l159_35_6};
  assign _zz__zz_realValue_0_35 = {1'd0, wReg};
  assign _zz__zz_realValue_0_35_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_35_1 = (_zz_realValue_0_35_2 + _zz_realValue_0_35_3);
  assign _zz_realValue_0_35_2 = {1'd0, wReg};
  assign _zz_realValue_0_35_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_35_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_35 = {1'd0, _zz_when_ArraySlice_l166_35_1};
  assign _zz_when_ArraySlice_l166_35_2 = (_zz_when_ArraySlice_l166_35_3 + _zz_when_ArraySlice_l166_35_7);
  assign _zz_when_ArraySlice_l166_35_3 = (realValue_0_35 - _zz_when_ArraySlice_l166_35_4);
  assign _zz_when_ArraySlice_l166_35_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_35_5);
  assign _zz_when_ArraySlice_l166_35_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_35_5 = {2'd0, _zz_when_ArraySlice_l166_35_6};
  assign _zz_when_ArraySlice_l166_35_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_36 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_36_1);
  assign _zz_when_ArraySlice_l158_36_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_36_1 = {1'd0, _zz_when_ArraySlice_l158_36_2};
  assign _zz_when_ArraySlice_l158_36_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_36_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_36 = {1'd0, _zz_when_ArraySlice_l159_36_1};
  assign _zz_when_ArraySlice_l159_36_2 = (_zz_when_ArraySlice_l159_36_3 - _zz_when_ArraySlice_l159_36_4);
  assign _zz_when_ArraySlice_l159_36_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_36_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_36_5);
  assign _zz_when_ArraySlice_l159_36_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_36_5 = {1'd0, _zz_when_ArraySlice_l159_36_6};
  assign _zz__zz_realValue_0_36 = {1'd0, wReg};
  assign _zz__zz_realValue_0_36_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_36_1 = (_zz_realValue_0_36_2 + _zz_realValue_0_36_3);
  assign _zz_realValue_0_36_2 = {1'd0, wReg};
  assign _zz_realValue_0_36_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_36_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_36 = {1'd0, _zz_when_ArraySlice_l166_36_1};
  assign _zz_when_ArraySlice_l166_36_2 = (_zz_when_ArraySlice_l166_36_3 + _zz_when_ArraySlice_l166_36_7);
  assign _zz_when_ArraySlice_l166_36_3 = (realValue_0_36 - _zz_when_ArraySlice_l166_36_4);
  assign _zz_when_ArraySlice_l166_36_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_36_5);
  assign _zz_when_ArraySlice_l166_36_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_36_5 = {1'd0, _zz_when_ArraySlice_l166_36_6};
  assign _zz_when_ArraySlice_l166_36_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_37 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_37_1);
  assign _zz_when_ArraySlice_l158_37_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_37_1 = {1'd0, _zz_when_ArraySlice_l158_37_2};
  assign _zz_when_ArraySlice_l158_37_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_37_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_37 = {2'd0, _zz_when_ArraySlice_l159_37_1};
  assign _zz_when_ArraySlice_l159_37_2 = (_zz_when_ArraySlice_l159_37_3 - _zz_when_ArraySlice_l159_37_4);
  assign _zz_when_ArraySlice_l159_37_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_37_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_37_5);
  assign _zz_when_ArraySlice_l159_37_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_37_5 = {1'd0, _zz_when_ArraySlice_l159_37_6};
  assign _zz__zz_realValue_0_37 = {1'd0, wReg};
  assign _zz__zz_realValue_0_37_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_37_1 = (_zz_realValue_0_37_2 + _zz_realValue_0_37_3);
  assign _zz_realValue_0_37_2 = {1'd0, wReg};
  assign _zz_realValue_0_37_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_37_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_37 = {2'd0, _zz_when_ArraySlice_l166_37_1};
  assign _zz_when_ArraySlice_l166_37_2 = (_zz_when_ArraySlice_l166_37_3 + _zz_when_ArraySlice_l166_37_7);
  assign _zz_when_ArraySlice_l166_37_3 = (realValue_0_37 - _zz_when_ArraySlice_l166_37_4);
  assign _zz_when_ArraySlice_l166_37_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_37_5);
  assign _zz_when_ArraySlice_l166_37_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_37_5 = {1'd0, _zz_when_ArraySlice_l166_37_6};
  assign _zz_when_ArraySlice_l166_37_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_38 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_38_1);
  assign _zz_when_ArraySlice_l158_38_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_38_1 = {1'd0, _zz_when_ArraySlice_l158_38_2};
  assign _zz_when_ArraySlice_l158_38_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_38_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_38 = {2'd0, _zz_when_ArraySlice_l159_38_1};
  assign _zz_when_ArraySlice_l159_38_2 = (_zz_when_ArraySlice_l159_38_3 - _zz_when_ArraySlice_l159_38_4);
  assign _zz_when_ArraySlice_l159_38_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_38_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_38_5);
  assign _zz_when_ArraySlice_l159_38_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_38_5 = {1'd0, _zz_when_ArraySlice_l159_38_6};
  assign _zz__zz_realValue_0_38 = {1'd0, wReg};
  assign _zz__zz_realValue_0_38_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_38_1 = (_zz_realValue_0_38_2 + _zz_realValue_0_38_3);
  assign _zz_realValue_0_38_2 = {1'd0, wReg};
  assign _zz_realValue_0_38_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_38_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_38 = {2'd0, _zz_when_ArraySlice_l166_38_1};
  assign _zz_when_ArraySlice_l166_38_2 = (_zz_when_ArraySlice_l166_38_3 + _zz_when_ArraySlice_l166_38_7);
  assign _zz_when_ArraySlice_l166_38_3 = (realValue_0_38 - _zz_when_ArraySlice_l166_38_4);
  assign _zz_when_ArraySlice_l166_38_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_38_5);
  assign _zz_when_ArraySlice_l166_38_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_38_5 = {1'd0, _zz_when_ArraySlice_l166_38_6};
  assign _zz_when_ArraySlice_l166_38_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_39 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_39_1);
  assign _zz_when_ArraySlice_l158_39_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_39_1 = {1'd0, _zz_when_ArraySlice_l158_39_2};
  assign _zz_when_ArraySlice_l158_39_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_39_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_39 = {3'd0, _zz_when_ArraySlice_l159_39_1};
  assign _zz_when_ArraySlice_l159_39_2 = (_zz_when_ArraySlice_l159_39_3 - _zz_when_ArraySlice_l159_39_4);
  assign _zz_when_ArraySlice_l159_39_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_39_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_39_5);
  assign _zz_when_ArraySlice_l159_39_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_39_5 = {1'd0, _zz_when_ArraySlice_l159_39_6};
  assign _zz__zz_realValue_0_39 = {1'd0, wReg};
  assign _zz__zz_realValue_0_39_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_39_1 = (_zz_realValue_0_39_2 + _zz_realValue_0_39_3);
  assign _zz_realValue_0_39_2 = {1'd0, wReg};
  assign _zz_realValue_0_39_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_39_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_39 = {3'd0, _zz_when_ArraySlice_l166_39_1};
  assign _zz_when_ArraySlice_l166_39_2 = (_zz_when_ArraySlice_l166_39_3 + _zz_when_ArraySlice_l166_39_7);
  assign _zz_when_ArraySlice_l166_39_3 = (realValue_0_39 - _zz_when_ArraySlice_l166_39_4);
  assign _zz_when_ArraySlice_l166_39_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_39_5);
  assign _zz_when_ArraySlice_l166_39_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_39_5 = {1'd0, _zz_when_ArraySlice_l166_39_6};
  assign _zz_when_ArraySlice_l166_39_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_1_2 = (_zz_when_ArraySlice_l403_1_3 + _zz_when_ArraySlice_l403_1_7);
  assign _zz_when_ArraySlice_l403_1_3 = (_zz_when_ArraySlice_l403_1_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l403_1_5);
  assign _zz_when_ArraySlice_l403_1_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_1_5 = {1'd0, _zz_when_ArraySlice_l403_1_6};
  assign _zz_when_ArraySlice_l403_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l403_1_7 = {3'd0, _zz_when_ArraySlice_l403_1_8};
  assign _zz_when_ArraySlice_l406_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_1_2 = (_zz_when_ArraySlice_l406_1_3 + 8'h01);
  assign _zz_when_ArraySlice_l406_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l406_1_4);
  assign _zz_when_ArraySlice_l406_1_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_1_4 = {1'd0, _zz_when_ArraySlice_l406_1_5};
  assign _zz_selectReadFifo_1_6 = (selectReadFifo_1 + _zz_selectReadFifo_1_7);
  assign _zz_selectReadFifo_1_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_7 = {1'd0, _zz_selectReadFifo_1_8};
  assign _zz_when_ArraySlice_l413_1_1 = (_zz_when_ArraySlice_l413_1_2 % aReg);
  assign _zz_when_ArraySlice_l413_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l417_1_4);
  assign _zz_when_ArraySlice_l417_1_2 = _zz_when_ArraySlice_l417_1_3[6:0];
  assign _zz_when_ArraySlice_l417_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l417_1_4 = {3'd0, _zz_when_ArraySlice_l417_1_5};
  assign _zz_when_ArraySlice_l418_1_2 = (_zz_when_ArraySlice_l418_1_3 - _zz_when_ArraySlice_l418_1_4);
  assign _zz_when_ArraySlice_l418_1_1 = {5'd0, _zz_when_ArraySlice_l418_1_2};
  assign _zz_when_ArraySlice_l418_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l418_1_4 = {7'd0, _zz_when_ArraySlice_l418_1_5};
  assign _zz__zz_realValue1_0_4 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_4_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_4_1 = (_zz_realValue1_0_4_2 + _zz_realValue1_0_4_3);
  assign _zz_realValue1_0_4_2 = {1'd0, hReg};
  assign _zz_realValue1_0_4_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l420_1_1 = {1'd0, _zz_when_ArraySlice_l420_1_2};
  assign _zz_when_ArraySlice_l420_1_3 = (realValue1_0_4 / aReg);
  assign _zz_selectReadFifo_1_9 = (selectReadFifo_1 - _zz_selectReadFifo_1_10);
  assign _zz_selectReadFifo_1_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_40 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_40_1);
  assign _zz_when_ArraySlice_l158_40_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_40_1 = {4'd0, _zz_when_ArraySlice_l158_40_2};
  assign _zz_when_ArraySlice_l158_40_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_40 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_40_1 = (_zz_when_ArraySlice_l159_40_2 - _zz_when_ArraySlice_l159_40_3);
  assign _zz_when_ArraySlice_l159_40_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_40_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_40_4);
  assign _zz_when_ArraySlice_l159_40_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_40_4 = {4'd0, _zz_when_ArraySlice_l159_40_5};
  assign _zz__zz_realValue_0_40 = {1'd0, wReg};
  assign _zz__zz_realValue_0_40_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_40_1 = (_zz_realValue_0_40_2 + _zz_realValue_0_40_3);
  assign _zz_realValue_0_40_2 = {1'd0, wReg};
  assign _zz_realValue_0_40_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_40 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_40_1 = (_zz_when_ArraySlice_l166_40_2 + _zz_when_ArraySlice_l166_40_6);
  assign _zz_when_ArraySlice_l166_40_2 = (realValue_0_40 - _zz_when_ArraySlice_l166_40_3);
  assign _zz_when_ArraySlice_l166_40_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_40_4);
  assign _zz_when_ArraySlice_l166_40_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_40_4 = {4'd0, _zz_when_ArraySlice_l166_40_5};
  assign _zz_when_ArraySlice_l166_40_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_41 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_41_1);
  assign _zz_when_ArraySlice_l158_41_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_41_1 = {3'd0, _zz_when_ArraySlice_l158_41_2};
  assign _zz_when_ArraySlice_l158_41_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_41_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_41 = {1'd0, _zz_when_ArraySlice_l159_41_1};
  assign _zz_when_ArraySlice_l159_41_2 = (_zz_when_ArraySlice_l159_41_3 - _zz_when_ArraySlice_l159_41_4);
  assign _zz_when_ArraySlice_l159_41_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_41_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_41_5);
  assign _zz_when_ArraySlice_l159_41_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_41_5 = {3'd0, _zz_when_ArraySlice_l159_41_6};
  assign _zz__zz_realValue_0_41 = {1'd0, wReg};
  assign _zz__zz_realValue_0_41_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_41_1 = (_zz_realValue_0_41_2 + _zz_realValue_0_41_3);
  assign _zz_realValue_0_41_2 = {1'd0, wReg};
  assign _zz_realValue_0_41_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_41_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_41 = {1'd0, _zz_when_ArraySlice_l166_41_1};
  assign _zz_when_ArraySlice_l166_41_2 = (_zz_when_ArraySlice_l166_41_3 + _zz_when_ArraySlice_l166_41_7);
  assign _zz_when_ArraySlice_l166_41_3 = (realValue_0_41 - _zz_when_ArraySlice_l166_41_4);
  assign _zz_when_ArraySlice_l166_41_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_41_5);
  assign _zz_when_ArraySlice_l166_41_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_41_5 = {3'd0, _zz_when_ArraySlice_l166_41_6};
  assign _zz_when_ArraySlice_l166_41_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_42 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_42_1);
  assign _zz_when_ArraySlice_l158_42_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_42_1 = {2'd0, _zz_when_ArraySlice_l158_42_2};
  assign _zz_when_ArraySlice_l158_42_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_42_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_42 = {1'd0, _zz_when_ArraySlice_l159_42_1};
  assign _zz_when_ArraySlice_l159_42_2 = (_zz_when_ArraySlice_l159_42_3 - _zz_when_ArraySlice_l159_42_4);
  assign _zz_when_ArraySlice_l159_42_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_42_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_42_5);
  assign _zz_when_ArraySlice_l159_42_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_42_5 = {2'd0, _zz_when_ArraySlice_l159_42_6};
  assign _zz__zz_realValue_0_42 = {1'd0, wReg};
  assign _zz__zz_realValue_0_42_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_42_1 = (_zz_realValue_0_42_2 + _zz_realValue_0_42_3);
  assign _zz_realValue_0_42_2 = {1'd0, wReg};
  assign _zz_realValue_0_42_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_42_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_42 = {1'd0, _zz_when_ArraySlice_l166_42_1};
  assign _zz_when_ArraySlice_l166_42_2 = (_zz_when_ArraySlice_l166_42_3 + _zz_when_ArraySlice_l166_42_7);
  assign _zz_when_ArraySlice_l166_42_3 = (realValue_0_42 - _zz_when_ArraySlice_l166_42_4);
  assign _zz_when_ArraySlice_l166_42_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_42_5);
  assign _zz_when_ArraySlice_l166_42_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_42_5 = {2'd0, _zz_when_ArraySlice_l166_42_6};
  assign _zz_when_ArraySlice_l166_42_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_43 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_43_1);
  assign _zz_when_ArraySlice_l158_43_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_43_1 = {2'd0, _zz_when_ArraySlice_l158_43_2};
  assign _zz_when_ArraySlice_l158_43_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_43_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_43 = {1'd0, _zz_when_ArraySlice_l159_43_1};
  assign _zz_when_ArraySlice_l159_43_2 = (_zz_when_ArraySlice_l159_43_3 - _zz_when_ArraySlice_l159_43_4);
  assign _zz_when_ArraySlice_l159_43_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_43_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_43_5);
  assign _zz_when_ArraySlice_l159_43_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_43_5 = {2'd0, _zz_when_ArraySlice_l159_43_6};
  assign _zz__zz_realValue_0_43 = {1'd0, wReg};
  assign _zz__zz_realValue_0_43_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_43_1 = (_zz_realValue_0_43_2 + _zz_realValue_0_43_3);
  assign _zz_realValue_0_43_2 = {1'd0, wReg};
  assign _zz_realValue_0_43_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_43_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_43 = {1'd0, _zz_when_ArraySlice_l166_43_1};
  assign _zz_when_ArraySlice_l166_43_2 = (_zz_when_ArraySlice_l166_43_3 + _zz_when_ArraySlice_l166_43_7);
  assign _zz_when_ArraySlice_l166_43_3 = (realValue_0_43 - _zz_when_ArraySlice_l166_43_4);
  assign _zz_when_ArraySlice_l166_43_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_43_5);
  assign _zz_when_ArraySlice_l166_43_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_43_5 = {2'd0, _zz_when_ArraySlice_l166_43_6};
  assign _zz_when_ArraySlice_l166_43_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_44 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_44_1);
  assign _zz_when_ArraySlice_l158_44_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_44_1 = {1'd0, _zz_when_ArraySlice_l158_44_2};
  assign _zz_when_ArraySlice_l158_44_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_44_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_44 = {1'd0, _zz_when_ArraySlice_l159_44_1};
  assign _zz_when_ArraySlice_l159_44_2 = (_zz_when_ArraySlice_l159_44_3 - _zz_when_ArraySlice_l159_44_4);
  assign _zz_when_ArraySlice_l159_44_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_44_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_44_5);
  assign _zz_when_ArraySlice_l159_44_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_44_5 = {1'd0, _zz_when_ArraySlice_l159_44_6};
  assign _zz__zz_realValue_0_44 = {1'd0, wReg};
  assign _zz__zz_realValue_0_44_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_44_1 = (_zz_realValue_0_44_2 + _zz_realValue_0_44_3);
  assign _zz_realValue_0_44_2 = {1'd0, wReg};
  assign _zz_realValue_0_44_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_44_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_44 = {1'd0, _zz_when_ArraySlice_l166_44_1};
  assign _zz_when_ArraySlice_l166_44_2 = (_zz_when_ArraySlice_l166_44_3 + _zz_when_ArraySlice_l166_44_7);
  assign _zz_when_ArraySlice_l166_44_3 = (realValue_0_44 - _zz_when_ArraySlice_l166_44_4);
  assign _zz_when_ArraySlice_l166_44_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_44_5);
  assign _zz_when_ArraySlice_l166_44_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_44_5 = {1'd0, _zz_when_ArraySlice_l166_44_6};
  assign _zz_when_ArraySlice_l166_44_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_45 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_45_1);
  assign _zz_when_ArraySlice_l158_45_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_45_1 = {1'd0, _zz_when_ArraySlice_l158_45_2};
  assign _zz_when_ArraySlice_l158_45_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_45_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_45 = {2'd0, _zz_when_ArraySlice_l159_45_1};
  assign _zz_when_ArraySlice_l159_45_2 = (_zz_when_ArraySlice_l159_45_3 - _zz_when_ArraySlice_l159_45_4);
  assign _zz_when_ArraySlice_l159_45_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_45_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_45_5);
  assign _zz_when_ArraySlice_l159_45_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_45_5 = {1'd0, _zz_when_ArraySlice_l159_45_6};
  assign _zz__zz_realValue_0_45 = {1'd0, wReg};
  assign _zz__zz_realValue_0_45_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_45_1 = (_zz_realValue_0_45_2 + _zz_realValue_0_45_3);
  assign _zz_realValue_0_45_2 = {1'd0, wReg};
  assign _zz_realValue_0_45_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_45_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_45 = {2'd0, _zz_when_ArraySlice_l166_45_1};
  assign _zz_when_ArraySlice_l166_45_2 = (_zz_when_ArraySlice_l166_45_3 + _zz_when_ArraySlice_l166_45_7);
  assign _zz_when_ArraySlice_l166_45_3 = (realValue_0_45 - _zz_when_ArraySlice_l166_45_4);
  assign _zz_when_ArraySlice_l166_45_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_45_5);
  assign _zz_when_ArraySlice_l166_45_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_45_5 = {1'd0, _zz_when_ArraySlice_l166_45_6};
  assign _zz_when_ArraySlice_l166_45_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_46 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_46_1);
  assign _zz_when_ArraySlice_l158_46_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_46_1 = {1'd0, _zz_when_ArraySlice_l158_46_2};
  assign _zz_when_ArraySlice_l158_46_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_46_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_46 = {2'd0, _zz_when_ArraySlice_l159_46_1};
  assign _zz_when_ArraySlice_l159_46_2 = (_zz_when_ArraySlice_l159_46_3 - _zz_when_ArraySlice_l159_46_4);
  assign _zz_when_ArraySlice_l159_46_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_46_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_46_5);
  assign _zz_when_ArraySlice_l159_46_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_46_5 = {1'd0, _zz_when_ArraySlice_l159_46_6};
  assign _zz__zz_realValue_0_46 = {1'd0, wReg};
  assign _zz__zz_realValue_0_46_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_46_1 = (_zz_realValue_0_46_2 + _zz_realValue_0_46_3);
  assign _zz_realValue_0_46_2 = {1'd0, wReg};
  assign _zz_realValue_0_46_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_46_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_46 = {2'd0, _zz_when_ArraySlice_l166_46_1};
  assign _zz_when_ArraySlice_l166_46_2 = (_zz_when_ArraySlice_l166_46_3 + _zz_when_ArraySlice_l166_46_7);
  assign _zz_when_ArraySlice_l166_46_3 = (realValue_0_46 - _zz_when_ArraySlice_l166_46_4);
  assign _zz_when_ArraySlice_l166_46_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_46_5);
  assign _zz_when_ArraySlice_l166_46_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_46_5 = {1'd0, _zz_when_ArraySlice_l166_46_6};
  assign _zz_when_ArraySlice_l166_46_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_47 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_47_1);
  assign _zz_when_ArraySlice_l158_47_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_47_1 = {1'd0, _zz_when_ArraySlice_l158_47_2};
  assign _zz_when_ArraySlice_l158_47_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_47_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_47 = {3'd0, _zz_when_ArraySlice_l159_47_1};
  assign _zz_when_ArraySlice_l159_47_2 = (_zz_when_ArraySlice_l159_47_3 - _zz_when_ArraySlice_l159_47_4);
  assign _zz_when_ArraySlice_l159_47_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_47_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_47_5);
  assign _zz_when_ArraySlice_l159_47_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_47_5 = {1'd0, _zz_when_ArraySlice_l159_47_6};
  assign _zz__zz_realValue_0_47 = {1'd0, wReg};
  assign _zz__zz_realValue_0_47_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_47_1 = (_zz_realValue_0_47_2 + _zz_realValue_0_47_3);
  assign _zz_realValue_0_47_2 = {1'd0, wReg};
  assign _zz_realValue_0_47_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_47_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_47 = {3'd0, _zz_when_ArraySlice_l166_47_1};
  assign _zz_when_ArraySlice_l166_47_2 = (_zz_when_ArraySlice_l166_47_3 + _zz_when_ArraySlice_l166_47_7);
  assign _zz_when_ArraySlice_l166_47_3 = (realValue_0_47 - _zz_when_ArraySlice_l166_47_4);
  assign _zz_when_ArraySlice_l166_47_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_47_5);
  assign _zz_when_ArraySlice_l166_47_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_47_5 = {1'd0, _zz_when_ArraySlice_l166_47_6};
  assign _zz_when_ArraySlice_l166_47_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_1_2 = (_zz_when_ArraySlice_l428_1_3 + _zz_when_ArraySlice_l428_1_7);
  assign _zz_when_ArraySlice_l428_1_3 = (_zz_when_ArraySlice_l428_1_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l428_1_5);
  assign _zz_when_ArraySlice_l428_1_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_1_5 = {1'd0, _zz_when_ArraySlice_l428_1_6};
  assign _zz_when_ArraySlice_l428_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l428_1_7 = {3'd0, _zz_when_ArraySlice_l428_1_8};
  assign _zz_when_ArraySlice_l431_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_1_2 = (_zz_when_ArraySlice_l431_1_3 + 8'h01);
  assign _zz_when_ArraySlice_l431_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l431_1_4);
  assign _zz_when_ArraySlice_l431_1_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_1_4 = {1'd0, _zz_when_ArraySlice_l431_1_5};
  assign _zz_selectReadFifo_1_11 = (selectReadFifo_1 + _zz_selectReadFifo_1_12);
  assign _zz_selectReadFifo_1_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_12 = {1'd0, _zz_selectReadFifo_1_13};
  assign _zz_when_ArraySlice_l438_1_1 = (_zz_when_ArraySlice_l438_1_2 % aReg);
  assign _zz_when_ArraySlice_l438_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_1_2 = (_zz_when_ArraySlice_l449_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l449_1_1 = {5'd0, _zz_when_ArraySlice_l449_1_2};
  assign _zz_when_ArraySlice_l449_1_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_5 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_5_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_5_1 = (_zz_realValue1_0_5_2 + _zz_realValue1_0_5_3);
  assign _zz_realValue1_0_5_2 = {1'd0, hReg};
  assign _zz_realValue1_0_5_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l450_1_1 = {1'd0, _zz_when_ArraySlice_l450_1_2};
  assign _zz_when_ArraySlice_l450_1_3 = (realValue1_0_5 / aReg);
  assign _zz_selectReadFifo_1_14 = (selectReadFifo_1 - _zz_selectReadFifo_1_15);
  assign _zz_selectReadFifo_1_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_48 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_48_1);
  assign _zz_when_ArraySlice_l158_48_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_48_1 = {4'd0, _zz_when_ArraySlice_l158_48_2};
  assign _zz_when_ArraySlice_l158_48_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_48 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_48_1 = (_zz_when_ArraySlice_l159_48_2 - _zz_when_ArraySlice_l159_48_3);
  assign _zz_when_ArraySlice_l159_48_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_48_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_48_4);
  assign _zz_when_ArraySlice_l159_48_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_48_4 = {4'd0, _zz_when_ArraySlice_l159_48_5};
  assign _zz__zz_realValue_0_48 = {1'd0, wReg};
  assign _zz__zz_realValue_0_48_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_48_1 = (_zz_realValue_0_48_2 + _zz_realValue_0_48_3);
  assign _zz_realValue_0_48_2 = {1'd0, wReg};
  assign _zz_realValue_0_48_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_48 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_48_1 = (_zz_when_ArraySlice_l166_48_2 + _zz_when_ArraySlice_l166_48_6);
  assign _zz_when_ArraySlice_l166_48_2 = (realValue_0_48 - _zz_when_ArraySlice_l166_48_3);
  assign _zz_when_ArraySlice_l166_48_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_48_4);
  assign _zz_when_ArraySlice_l166_48_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_48_4 = {4'd0, _zz_when_ArraySlice_l166_48_5};
  assign _zz_when_ArraySlice_l166_48_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_49 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_49_1);
  assign _zz_when_ArraySlice_l158_49_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_49_1 = {3'd0, _zz_when_ArraySlice_l158_49_2};
  assign _zz_when_ArraySlice_l158_49_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_49_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_49 = {1'd0, _zz_when_ArraySlice_l159_49_1};
  assign _zz_when_ArraySlice_l159_49_2 = (_zz_when_ArraySlice_l159_49_3 - _zz_when_ArraySlice_l159_49_4);
  assign _zz_when_ArraySlice_l159_49_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_49_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_49_5);
  assign _zz_when_ArraySlice_l159_49_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_49_5 = {3'd0, _zz_when_ArraySlice_l159_49_6};
  assign _zz__zz_realValue_0_49 = {1'd0, wReg};
  assign _zz__zz_realValue_0_49_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_49_1 = (_zz_realValue_0_49_2 + _zz_realValue_0_49_3);
  assign _zz_realValue_0_49_2 = {1'd0, wReg};
  assign _zz_realValue_0_49_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_49_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_49 = {1'd0, _zz_when_ArraySlice_l166_49_1};
  assign _zz_when_ArraySlice_l166_49_2 = (_zz_when_ArraySlice_l166_49_3 + _zz_when_ArraySlice_l166_49_7);
  assign _zz_when_ArraySlice_l166_49_3 = (realValue_0_49 - _zz_when_ArraySlice_l166_49_4);
  assign _zz_when_ArraySlice_l166_49_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_49_5);
  assign _zz_when_ArraySlice_l166_49_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_49_5 = {3'd0, _zz_when_ArraySlice_l166_49_6};
  assign _zz_when_ArraySlice_l166_49_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_50 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_50_1);
  assign _zz_when_ArraySlice_l158_50_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_50_1 = {2'd0, _zz_when_ArraySlice_l158_50_2};
  assign _zz_when_ArraySlice_l158_50_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_50_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_50 = {1'd0, _zz_when_ArraySlice_l159_50_1};
  assign _zz_when_ArraySlice_l159_50_2 = (_zz_when_ArraySlice_l159_50_3 - _zz_when_ArraySlice_l159_50_4);
  assign _zz_when_ArraySlice_l159_50_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_50_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_50_5);
  assign _zz_when_ArraySlice_l159_50_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_50_5 = {2'd0, _zz_when_ArraySlice_l159_50_6};
  assign _zz__zz_realValue_0_50 = {1'd0, wReg};
  assign _zz__zz_realValue_0_50_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_50_1 = (_zz_realValue_0_50_2 + _zz_realValue_0_50_3);
  assign _zz_realValue_0_50_2 = {1'd0, wReg};
  assign _zz_realValue_0_50_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_50_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_50 = {1'd0, _zz_when_ArraySlice_l166_50_1};
  assign _zz_when_ArraySlice_l166_50_2 = (_zz_when_ArraySlice_l166_50_3 + _zz_when_ArraySlice_l166_50_7);
  assign _zz_when_ArraySlice_l166_50_3 = (realValue_0_50 - _zz_when_ArraySlice_l166_50_4);
  assign _zz_when_ArraySlice_l166_50_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_50_5);
  assign _zz_when_ArraySlice_l166_50_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_50_5 = {2'd0, _zz_when_ArraySlice_l166_50_6};
  assign _zz_when_ArraySlice_l166_50_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_51 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_51_1);
  assign _zz_when_ArraySlice_l158_51_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_51_1 = {2'd0, _zz_when_ArraySlice_l158_51_2};
  assign _zz_when_ArraySlice_l158_51_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_51_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_51 = {1'd0, _zz_when_ArraySlice_l159_51_1};
  assign _zz_when_ArraySlice_l159_51_2 = (_zz_when_ArraySlice_l159_51_3 - _zz_when_ArraySlice_l159_51_4);
  assign _zz_when_ArraySlice_l159_51_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_51_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_51_5);
  assign _zz_when_ArraySlice_l159_51_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_51_5 = {2'd0, _zz_when_ArraySlice_l159_51_6};
  assign _zz__zz_realValue_0_51 = {1'd0, wReg};
  assign _zz__zz_realValue_0_51_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_51_1 = (_zz_realValue_0_51_2 + _zz_realValue_0_51_3);
  assign _zz_realValue_0_51_2 = {1'd0, wReg};
  assign _zz_realValue_0_51_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_51_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_51 = {1'd0, _zz_when_ArraySlice_l166_51_1};
  assign _zz_when_ArraySlice_l166_51_2 = (_zz_when_ArraySlice_l166_51_3 + _zz_when_ArraySlice_l166_51_7);
  assign _zz_when_ArraySlice_l166_51_3 = (realValue_0_51 - _zz_when_ArraySlice_l166_51_4);
  assign _zz_when_ArraySlice_l166_51_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_51_5);
  assign _zz_when_ArraySlice_l166_51_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_51_5 = {2'd0, _zz_when_ArraySlice_l166_51_6};
  assign _zz_when_ArraySlice_l166_51_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_52 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_52_1);
  assign _zz_when_ArraySlice_l158_52_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_52_1 = {1'd0, _zz_when_ArraySlice_l158_52_2};
  assign _zz_when_ArraySlice_l158_52_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_52_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_52 = {1'd0, _zz_when_ArraySlice_l159_52_1};
  assign _zz_when_ArraySlice_l159_52_2 = (_zz_when_ArraySlice_l159_52_3 - _zz_when_ArraySlice_l159_52_4);
  assign _zz_when_ArraySlice_l159_52_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_52_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_52_5);
  assign _zz_when_ArraySlice_l159_52_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_52_5 = {1'd0, _zz_when_ArraySlice_l159_52_6};
  assign _zz__zz_realValue_0_52 = {1'd0, wReg};
  assign _zz__zz_realValue_0_52_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_52_1 = (_zz_realValue_0_52_2 + _zz_realValue_0_52_3);
  assign _zz_realValue_0_52_2 = {1'd0, wReg};
  assign _zz_realValue_0_52_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_52_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_52 = {1'd0, _zz_when_ArraySlice_l166_52_1};
  assign _zz_when_ArraySlice_l166_52_2 = (_zz_when_ArraySlice_l166_52_3 + _zz_when_ArraySlice_l166_52_7);
  assign _zz_when_ArraySlice_l166_52_3 = (realValue_0_52 - _zz_when_ArraySlice_l166_52_4);
  assign _zz_when_ArraySlice_l166_52_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_52_5);
  assign _zz_when_ArraySlice_l166_52_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_52_5 = {1'd0, _zz_when_ArraySlice_l166_52_6};
  assign _zz_when_ArraySlice_l166_52_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_53 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_53_1);
  assign _zz_when_ArraySlice_l158_53_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_53_1 = {1'd0, _zz_when_ArraySlice_l158_53_2};
  assign _zz_when_ArraySlice_l158_53_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_53_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_53 = {2'd0, _zz_when_ArraySlice_l159_53_1};
  assign _zz_when_ArraySlice_l159_53_2 = (_zz_when_ArraySlice_l159_53_3 - _zz_when_ArraySlice_l159_53_4);
  assign _zz_when_ArraySlice_l159_53_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_53_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_53_5);
  assign _zz_when_ArraySlice_l159_53_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_53_5 = {1'd0, _zz_when_ArraySlice_l159_53_6};
  assign _zz__zz_realValue_0_53 = {1'd0, wReg};
  assign _zz__zz_realValue_0_53_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_53_1 = (_zz_realValue_0_53_2 + _zz_realValue_0_53_3);
  assign _zz_realValue_0_53_2 = {1'd0, wReg};
  assign _zz_realValue_0_53_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_53_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_53 = {2'd0, _zz_when_ArraySlice_l166_53_1};
  assign _zz_when_ArraySlice_l166_53_2 = (_zz_when_ArraySlice_l166_53_3 + _zz_when_ArraySlice_l166_53_7);
  assign _zz_when_ArraySlice_l166_53_3 = (realValue_0_53 - _zz_when_ArraySlice_l166_53_4);
  assign _zz_when_ArraySlice_l166_53_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_53_5);
  assign _zz_when_ArraySlice_l166_53_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_53_5 = {1'd0, _zz_when_ArraySlice_l166_53_6};
  assign _zz_when_ArraySlice_l166_53_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_54 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_54_1);
  assign _zz_when_ArraySlice_l158_54_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_54_1 = {1'd0, _zz_when_ArraySlice_l158_54_2};
  assign _zz_when_ArraySlice_l158_54_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_54_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_54 = {2'd0, _zz_when_ArraySlice_l159_54_1};
  assign _zz_when_ArraySlice_l159_54_2 = (_zz_when_ArraySlice_l159_54_3 - _zz_when_ArraySlice_l159_54_4);
  assign _zz_when_ArraySlice_l159_54_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_54_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_54_5);
  assign _zz_when_ArraySlice_l159_54_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_54_5 = {1'd0, _zz_when_ArraySlice_l159_54_6};
  assign _zz__zz_realValue_0_54 = {1'd0, wReg};
  assign _zz__zz_realValue_0_54_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_54_1 = (_zz_realValue_0_54_2 + _zz_realValue_0_54_3);
  assign _zz_realValue_0_54_2 = {1'd0, wReg};
  assign _zz_realValue_0_54_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_54_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_54 = {2'd0, _zz_when_ArraySlice_l166_54_1};
  assign _zz_when_ArraySlice_l166_54_2 = (_zz_when_ArraySlice_l166_54_3 + _zz_when_ArraySlice_l166_54_7);
  assign _zz_when_ArraySlice_l166_54_3 = (realValue_0_54 - _zz_when_ArraySlice_l166_54_4);
  assign _zz_when_ArraySlice_l166_54_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_54_5);
  assign _zz_when_ArraySlice_l166_54_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_54_5 = {1'd0, _zz_when_ArraySlice_l166_54_6};
  assign _zz_when_ArraySlice_l166_54_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_55 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_55_1);
  assign _zz_when_ArraySlice_l158_55_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_55_1 = {1'd0, _zz_when_ArraySlice_l158_55_2};
  assign _zz_when_ArraySlice_l158_55_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_55_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_55 = {3'd0, _zz_when_ArraySlice_l159_55_1};
  assign _zz_when_ArraySlice_l159_55_2 = (_zz_when_ArraySlice_l159_55_3 - _zz_when_ArraySlice_l159_55_4);
  assign _zz_when_ArraySlice_l159_55_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_55_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_55_5);
  assign _zz_when_ArraySlice_l159_55_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_55_5 = {1'd0, _zz_when_ArraySlice_l159_55_6};
  assign _zz__zz_realValue_0_55 = {1'd0, wReg};
  assign _zz__zz_realValue_0_55_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_55_1 = (_zz_realValue_0_55_2 + _zz_realValue_0_55_3);
  assign _zz_realValue_0_55_2 = {1'd0, wReg};
  assign _zz_realValue_0_55_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_55_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_55 = {3'd0, _zz_when_ArraySlice_l166_55_1};
  assign _zz_when_ArraySlice_l166_55_2 = (_zz_when_ArraySlice_l166_55_3 + _zz_when_ArraySlice_l166_55_7);
  assign _zz_when_ArraySlice_l166_55_3 = (realValue_0_55 - _zz_when_ArraySlice_l166_55_4);
  assign _zz_when_ArraySlice_l166_55_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_55_5);
  assign _zz_when_ArraySlice_l166_55_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_55_5 = {1'd0, _zz_when_ArraySlice_l166_55_6};
  assign _zz_when_ArraySlice_l166_55_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_1_1 = (_zz_when_ArraySlice_l461_1_2 % aReg);
  assign _zz_when_ArraySlice_l461_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l447_1_3);
  assign _zz_when_ArraySlice_l447_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l447_1_3 = {3'd0, _zz_when_ArraySlice_l447_1_4};
  assign _zz_when_ArraySlice_l468_1_2 = (_zz_when_ArraySlice_l468_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l468_1_1 = {5'd0, _zz_when_ArraySlice_l468_1_2};
  assign _zz_when_ArraySlice_l468_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l376_2_2);
  assign _zz_when_ArraySlice_l376_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l376_2_2 = {2'd0, _zz_when_ArraySlice_l376_2_3};
  assign _zz_when_ArraySlice_l376_2_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l377_2_4);
  assign _zz_when_ArraySlice_l377_2_2 = _zz_when_ArraySlice_l377_2_3[6:0];
  assign _zz_when_ArraySlice_l377_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l377_2_4 = {2'd0, _zz_when_ArraySlice_l377_2_5};
  assign _zz__zz_outputStreamArrayData_2_valid_1 = (bReg * 2'b10);
  assign _zz__zz_outputStreamArrayData_2_valid = {2'd0, _zz__zz_outputStreamArrayData_2_valid_1};
  assign _zz__zz_5 = _zz_outputStreamArrayData_2_valid[6:0];
  assign _zz_outputStreamArrayData_2_valid_3 = _zz_outputStreamArrayData_2_valid[6:0];
  assign _zz_outputStreamArrayData_2_payload_1 = _zz_outputStreamArrayData_2_valid[6:0];
  assign _zz_when_ArraySlice_l383_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l383_2_4);
  assign _zz_when_ArraySlice_l383_2_2 = _zz_when_ArraySlice_l383_2_3[6:0];
  assign _zz_when_ArraySlice_l383_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l383_2_4 = {2'd0, _zz_when_ArraySlice_l383_2_5};
  assign _zz_when_ArraySlice_l384_2_2 = (_zz_when_ArraySlice_l384_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l384_2_1 = {5'd0, _zz_when_ArraySlice_l384_2_2};
  assign _zz_when_ArraySlice_l384_2_3 = (bReg * aReg);
  assign _zz_selectReadFifo_2 = (selectReadFifo_2 - _zz_selectReadFifo_2_1);
  assign _zz_selectReadFifo_2_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_2 = (_zz_when_ArraySlice_l387_2_1 % aReg);
  assign _zz_when_ArraySlice_l387_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l392_2_4);
  assign _zz_when_ArraySlice_l392_2_2 = _zz_when_ArraySlice_l392_2_3[6:0];
  assign _zz_when_ArraySlice_l392_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l392_2_4 = {2'd0, _zz_when_ArraySlice_l392_2_5};
  assign _zz_when_ArraySlice_l393_2_2 = (_zz_when_ArraySlice_l393_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l393_2_1 = {5'd0, _zz_when_ArraySlice_l393_2_2};
  assign _zz_when_ArraySlice_l393_2_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_6 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_6_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_6_1 = (_zz_realValue1_0_6_2 + _zz_realValue1_0_6_3);
  assign _zz_realValue1_0_6_2 = {1'd0, hReg};
  assign _zz_realValue1_0_6_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l395_2_1 = {1'd0, _zz_when_ArraySlice_l395_2_2};
  assign _zz_when_ArraySlice_l395_2_3 = (realValue1_0_6 / aReg);
  assign _zz_selectReadFifo_2_2 = (selectReadFifo_2 - _zz_selectReadFifo_2_3);
  assign _zz_selectReadFifo_2_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_2_5 = 1'b1;
  assign _zz_selectReadFifo_2_4 = {7'd0, _zz_selectReadFifo_2_5};
  assign _zz_when_ArraySlice_l158_56 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_56_1);
  assign _zz_when_ArraySlice_l158_56_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_56_1 = {4'd0, _zz_when_ArraySlice_l158_56_2};
  assign _zz_when_ArraySlice_l158_56_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_56 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_56_1 = (_zz_when_ArraySlice_l159_56_2 - _zz_when_ArraySlice_l159_56_3);
  assign _zz_when_ArraySlice_l159_56_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_56_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_56_4);
  assign _zz_when_ArraySlice_l159_56_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_56_4 = {4'd0, _zz_when_ArraySlice_l159_56_5};
  assign _zz__zz_realValue_0_56 = {1'd0, wReg};
  assign _zz__zz_realValue_0_56_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_56_1 = (_zz_realValue_0_56_2 + _zz_realValue_0_56_3);
  assign _zz_realValue_0_56_2 = {1'd0, wReg};
  assign _zz_realValue_0_56_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_56 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_56_1 = (_zz_when_ArraySlice_l166_56_2 + _zz_when_ArraySlice_l166_56_6);
  assign _zz_when_ArraySlice_l166_56_2 = (realValue_0_56 - _zz_when_ArraySlice_l166_56_3);
  assign _zz_when_ArraySlice_l166_56_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_56_4);
  assign _zz_when_ArraySlice_l166_56_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_56_4 = {4'd0, _zz_when_ArraySlice_l166_56_5};
  assign _zz_when_ArraySlice_l166_56_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_57 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_57_1);
  assign _zz_when_ArraySlice_l158_57_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_57_1 = {3'd0, _zz_when_ArraySlice_l158_57_2};
  assign _zz_when_ArraySlice_l158_57_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_57_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_57 = {1'd0, _zz_when_ArraySlice_l159_57_1};
  assign _zz_when_ArraySlice_l159_57_2 = (_zz_when_ArraySlice_l159_57_3 - _zz_when_ArraySlice_l159_57_4);
  assign _zz_when_ArraySlice_l159_57_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_57_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_57_5);
  assign _zz_when_ArraySlice_l159_57_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_57_5 = {3'd0, _zz_when_ArraySlice_l159_57_6};
  assign _zz__zz_realValue_0_57 = {1'd0, wReg};
  assign _zz__zz_realValue_0_57_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_57_1 = (_zz_realValue_0_57_2 + _zz_realValue_0_57_3);
  assign _zz_realValue_0_57_2 = {1'd0, wReg};
  assign _zz_realValue_0_57_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_57_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_57 = {1'd0, _zz_when_ArraySlice_l166_57_1};
  assign _zz_when_ArraySlice_l166_57_2 = (_zz_when_ArraySlice_l166_57_3 + _zz_when_ArraySlice_l166_57_7);
  assign _zz_when_ArraySlice_l166_57_3 = (realValue_0_57 - _zz_when_ArraySlice_l166_57_4);
  assign _zz_when_ArraySlice_l166_57_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_57_5);
  assign _zz_when_ArraySlice_l166_57_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_57_5 = {3'd0, _zz_when_ArraySlice_l166_57_6};
  assign _zz_when_ArraySlice_l166_57_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_58 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_58_1);
  assign _zz_when_ArraySlice_l158_58_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_58_1 = {2'd0, _zz_when_ArraySlice_l158_58_2};
  assign _zz_when_ArraySlice_l158_58_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_58_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_58 = {1'd0, _zz_when_ArraySlice_l159_58_1};
  assign _zz_when_ArraySlice_l159_58_2 = (_zz_when_ArraySlice_l159_58_3 - _zz_when_ArraySlice_l159_58_4);
  assign _zz_when_ArraySlice_l159_58_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_58_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_58_5);
  assign _zz_when_ArraySlice_l159_58_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_58_5 = {2'd0, _zz_when_ArraySlice_l159_58_6};
  assign _zz__zz_realValue_0_58 = {1'd0, wReg};
  assign _zz__zz_realValue_0_58_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_58_1 = (_zz_realValue_0_58_2 + _zz_realValue_0_58_3);
  assign _zz_realValue_0_58_2 = {1'd0, wReg};
  assign _zz_realValue_0_58_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_58_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_58 = {1'd0, _zz_when_ArraySlice_l166_58_1};
  assign _zz_when_ArraySlice_l166_58_2 = (_zz_when_ArraySlice_l166_58_3 + _zz_when_ArraySlice_l166_58_7);
  assign _zz_when_ArraySlice_l166_58_3 = (realValue_0_58 - _zz_when_ArraySlice_l166_58_4);
  assign _zz_when_ArraySlice_l166_58_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_58_5);
  assign _zz_when_ArraySlice_l166_58_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_58_5 = {2'd0, _zz_when_ArraySlice_l166_58_6};
  assign _zz_when_ArraySlice_l166_58_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_59 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_59_1);
  assign _zz_when_ArraySlice_l158_59_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_59_1 = {2'd0, _zz_when_ArraySlice_l158_59_2};
  assign _zz_when_ArraySlice_l158_59_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_59_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_59 = {1'd0, _zz_when_ArraySlice_l159_59_1};
  assign _zz_when_ArraySlice_l159_59_2 = (_zz_when_ArraySlice_l159_59_3 - _zz_when_ArraySlice_l159_59_4);
  assign _zz_when_ArraySlice_l159_59_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_59_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_59_5);
  assign _zz_when_ArraySlice_l159_59_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_59_5 = {2'd0, _zz_when_ArraySlice_l159_59_6};
  assign _zz__zz_realValue_0_59 = {1'd0, wReg};
  assign _zz__zz_realValue_0_59_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_59_1 = (_zz_realValue_0_59_2 + _zz_realValue_0_59_3);
  assign _zz_realValue_0_59_2 = {1'd0, wReg};
  assign _zz_realValue_0_59_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_59_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_59 = {1'd0, _zz_when_ArraySlice_l166_59_1};
  assign _zz_when_ArraySlice_l166_59_2 = (_zz_when_ArraySlice_l166_59_3 + _zz_when_ArraySlice_l166_59_7);
  assign _zz_when_ArraySlice_l166_59_3 = (realValue_0_59 - _zz_when_ArraySlice_l166_59_4);
  assign _zz_when_ArraySlice_l166_59_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_59_5);
  assign _zz_when_ArraySlice_l166_59_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_59_5 = {2'd0, _zz_when_ArraySlice_l166_59_6};
  assign _zz_when_ArraySlice_l166_59_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_60 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_60_1);
  assign _zz_when_ArraySlice_l158_60_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_60_1 = {1'd0, _zz_when_ArraySlice_l158_60_2};
  assign _zz_when_ArraySlice_l158_60_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_60_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_60 = {1'd0, _zz_when_ArraySlice_l159_60_1};
  assign _zz_when_ArraySlice_l159_60_2 = (_zz_when_ArraySlice_l159_60_3 - _zz_when_ArraySlice_l159_60_4);
  assign _zz_when_ArraySlice_l159_60_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_60_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_60_5);
  assign _zz_when_ArraySlice_l159_60_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_60_5 = {1'd0, _zz_when_ArraySlice_l159_60_6};
  assign _zz__zz_realValue_0_60 = {1'd0, wReg};
  assign _zz__zz_realValue_0_60_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_60_1 = (_zz_realValue_0_60_2 + _zz_realValue_0_60_3);
  assign _zz_realValue_0_60_2 = {1'd0, wReg};
  assign _zz_realValue_0_60_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_60_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_60 = {1'd0, _zz_when_ArraySlice_l166_60_1};
  assign _zz_when_ArraySlice_l166_60_2 = (_zz_when_ArraySlice_l166_60_3 + _zz_when_ArraySlice_l166_60_7);
  assign _zz_when_ArraySlice_l166_60_3 = (realValue_0_60 - _zz_when_ArraySlice_l166_60_4);
  assign _zz_when_ArraySlice_l166_60_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_60_5);
  assign _zz_when_ArraySlice_l166_60_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_60_5 = {1'd0, _zz_when_ArraySlice_l166_60_6};
  assign _zz_when_ArraySlice_l166_60_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_61 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_61_1);
  assign _zz_when_ArraySlice_l158_61_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_61_1 = {1'd0, _zz_when_ArraySlice_l158_61_2};
  assign _zz_when_ArraySlice_l158_61_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_61_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_61 = {2'd0, _zz_when_ArraySlice_l159_61_1};
  assign _zz_when_ArraySlice_l159_61_2 = (_zz_when_ArraySlice_l159_61_3 - _zz_when_ArraySlice_l159_61_4);
  assign _zz_when_ArraySlice_l159_61_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_61_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_61_5);
  assign _zz_when_ArraySlice_l159_61_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_61_5 = {1'd0, _zz_when_ArraySlice_l159_61_6};
  assign _zz__zz_realValue_0_61 = {1'd0, wReg};
  assign _zz__zz_realValue_0_61_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_61_1 = (_zz_realValue_0_61_2 + _zz_realValue_0_61_3);
  assign _zz_realValue_0_61_2 = {1'd0, wReg};
  assign _zz_realValue_0_61_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_61_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_61 = {2'd0, _zz_when_ArraySlice_l166_61_1};
  assign _zz_when_ArraySlice_l166_61_2 = (_zz_when_ArraySlice_l166_61_3 + _zz_when_ArraySlice_l166_61_7);
  assign _zz_when_ArraySlice_l166_61_3 = (realValue_0_61 - _zz_when_ArraySlice_l166_61_4);
  assign _zz_when_ArraySlice_l166_61_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_61_5);
  assign _zz_when_ArraySlice_l166_61_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_61_5 = {1'd0, _zz_when_ArraySlice_l166_61_6};
  assign _zz_when_ArraySlice_l166_61_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_62 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_62_1);
  assign _zz_when_ArraySlice_l158_62_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_62_1 = {1'd0, _zz_when_ArraySlice_l158_62_2};
  assign _zz_when_ArraySlice_l158_62_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_62_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_62 = {2'd0, _zz_when_ArraySlice_l159_62_1};
  assign _zz_when_ArraySlice_l159_62_2 = (_zz_when_ArraySlice_l159_62_3 - _zz_when_ArraySlice_l159_62_4);
  assign _zz_when_ArraySlice_l159_62_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_62_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_62_5);
  assign _zz_when_ArraySlice_l159_62_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_62_5 = {1'd0, _zz_when_ArraySlice_l159_62_6};
  assign _zz__zz_realValue_0_62 = {1'd0, wReg};
  assign _zz__zz_realValue_0_62_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_62_1 = (_zz_realValue_0_62_2 + _zz_realValue_0_62_3);
  assign _zz_realValue_0_62_2 = {1'd0, wReg};
  assign _zz_realValue_0_62_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_62_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_62 = {2'd0, _zz_when_ArraySlice_l166_62_1};
  assign _zz_when_ArraySlice_l166_62_2 = (_zz_when_ArraySlice_l166_62_3 + _zz_when_ArraySlice_l166_62_7);
  assign _zz_when_ArraySlice_l166_62_3 = (realValue_0_62 - _zz_when_ArraySlice_l166_62_4);
  assign _zz_when_ArraySlice_l166_62_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_62_5);
  assign _zz_when_ArraySlice_l166_62_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_62_5 = {1'd0, _zz_when_ArraySlice_l166_62_6};
  assign _zz_when_ArraySlice_l166_62_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_63 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_63_1);
  assign _zz_when_ArraySlice_l158_63_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_63_1 = {1'd0, _zz_when_ArraySlice_l158_63_2};
  assign _zz_when_ArraySlice_l158_63_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_63_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_63 = {3'd0, _zz_when_ArraySlice_l159_63_1};
  assign _zz_when_ArraySlice_l159_63_2 = (_zz_when_ArraySlice_l159_63_3 - _zz_when_ArraySlice_l159_63_4);
  assign _zz_when_ArraySlice_l159_63_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_63_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_63_5);
  assign _zz_when_ArraySlice_l159_63_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_63_5 = {1'd0, _zz_when_ArraySlice_l159_63_6};
  assign _zz__zz_realValue_0_63 = {1'd0, wReg};
  assign _zz__zz_realValue_0_63_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_63_1 = (_zz_realValue_0_63_2 + _zz_realValue_0_63_3);
  assign _zz_realValue_0_63_2 = {1'd0, wReg};
  assign _zz_realValue_0_63_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_63_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_63 = {3'd0, _zz_when_ArraySlice_l166_63_1};
  assign _zz_when_ArraySlice_l166_63_2 = (_zz_when_ArraySlice_l166_63_3 + _zz_when_ArraySlice_l166_63_7);
  assign _zz_when_ArraySlice_l166_63_3 = (realValue_0_63 - _zz_when_ArraySlice_l166_63_4);
  assign _zz_when_ArraySlice_l166_63_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_63_5);
  assign _zz_when_ArraySlice_l166_63_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_63_5 = {1'd0, _zz_when_ArraySlice_l166_63_6};
  assign _zz_when_ArraySlice_l166_63_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_2_2 = (_zz_when_ArraySlice_l403_2_3 + _zz_when_ArraySlice_l403_2_7);
  assign _zz_when_ArraySlice_l403_2_3 = (_zz_when_ArraySlice_l403_2_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l403_2_5);
  assign _zz_when_ArraySlice_l403_2_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_2_5 = {1'd0, _zz_when_ArraySlice_l403_2_6};
  assign _zz_when_ArraySlice_l403_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l403_2_7 = {2'd0, _zz_when_ArraySlice_l403_2_8};
  assign _zz_when_ArraySlice_l406_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_2_2 = (_zz_when_ArraySlice_l406_2_3 + 8'h01);
  assign _zz_when_ArraySlice_l406_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l406_2_4);
  assign _zz_when_ArraySlice_l406_2_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_2_4 = {1'd0, _zz_when_ArraySlice_l406_2_5};
  assign _zz_selectReadFifo_2_6 = (selectReadFifo_2 + _zz_selectReadFifo_2_7);
  assign _zz_selectReadFifo_2_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_7 = {1'd0, _zz_selectReadFifo_2_8};
  assign _zz_when_ArraySlice_l413_2 = (_zz_when_ArraySlice_l413_2_1 % aReg);
  assign _zz_when_ArraySlice_l413_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l417_2_4);
  assign _zz_when_ArraySlice_l417_2_2 = _zz_when_ArraySlice_l417_2_3[6:0];
  assign _zz_when_ArraySlice_l417_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l417_2_4 = {2'd0, _zz_when_ArraySlice_l417_2_5};
  assign _zz_when_ArraySlice_l418_2_2 = (_zz_when_ArraySlice_l418_2_3 - _zz_when_ArraySlice_l418_2_4);
  assign _zz_when_ArraySlice_l418_2_1 = {5'd0, _zz_when_ArraySlice_l418_2_2};
  assign _zz_when_ArraySlice_l418_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l418_2_4 = {7'd0, _zz_when_ArraySlice_l418_2_5};
  assign _zz__zz_realValue1_0_7 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_7_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_7_1 = (_zz_realValue1_0_7_2 + _zz_realValue1_0_7_3);
  assign _zz_realValue1_0_7_2 = {1'd0, hReg};
  assign _zz_realValue1_0_7_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l420_2_1 = {1'd0, _zz_when_ArraySlice_l420_2_2};
  assign _zz_when_ArraySlice_l420_2_3 = (realValue1_0_7 / aReg);
  assign _zz_selectReadFifo_2_9 = (selectReadFifo_2 - _zz_selectReadFifo_2_10);
  assign _zz_selectReadFifo_2_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_64 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_64_1);
  assign _zz_when_ArraySlice_l158_64_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_64_1 = {4'd0, _zz_when_ArraySlice_l158_64_2};
  assign _zz_when_ArraySlice_l158_64_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_64 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_64_1 = (_zz_when_ArraySlice_l159_64_2 - _zz_when_ArraySlice_l159_64_3);
  assign _zz_when_ArraySlice_l159_64_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_64_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_64_4);
  assign _zz_when_ArraySlice_l159_64_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_64_4 = {4'd0, _zz_when_ArraySlice_l159_64_5};
  assign _zz__zz_realValue_0_64 = {1'd0, wReg};
  assign _zz__zz_realValue_0_64_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_64_1 = (_zz_realValue_0_64_2 + _zz_realValue_0_64_3);
  assign _zz_realValue_0_64_2 = {1'd0, wReg};
  assign _zz_realValue_0_64_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_64 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_64_1 = (_zz_when_ArraySlice_l166_64_2 + _zz_when_ArraySlice_l166_64_6);
  assign _zz_when_ArraySlice_l166_64_2 = (realValue_0_64 - _zz_when_ArraySlice_l166_64_3);
  assign _zz_when_ArraySlice_l166_64_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_64_4);
  assign _zz_when_ArraySlice_l166_64_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_64_4 = {4'd0, _zz_when_ArraySlice_l166_64_5};
  assign _zz_when_ArraySlice_l166_64_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_65 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_65_1);
  assign _zz_when_ArraySlice_l158_65_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_65_1 = {3'd0, _zz_when_ArraySlice_l158_65_2};
  assign _zz_when_ArraySlice_l158_65_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_65_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_65 = {1'd0, _zz_when_ArraySlice_l159_65_1};
  assign _zz_when_ArraySlice_l159_65_2 = (_zz_when_ArraySlice_l159_65_3 - _zz_when_ArraySlice_l159_65_4);
  assign _zz_when_ArraySlice_l159_65_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_65_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_65_5);
  assign _zz_when_ArraySlice_l159_65_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_65_5 = {3'd0, _zz_when_ArraySlice_l159_65_6};
  assign _zz__zz_realValue_0_65 = {1'd0, wReg};
  assign _zz__zz_realValue_0_65_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_65_1 = (_zz_realValue_0_65_2 + _zz_realValue_0_65_3);
  assign _zz_realValue_0_65_2 = {1'd0, wReg};
  assign _zz_realValue_0_65_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_65_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_65 = {1'd0, _zz_when_ArraySlice_l166_65_1};
  assign _zz_when_ArraySlice_l166_65_2 = (_zz_when_ArraySlice_l166_65_3 + _zz_when_ArraySlice_l166_65_7);
  assign _zz_when_ArraySlice_l166_65_3 = (realValue_0_65 - _zz_when_ArraySlice_l166_65_4);
  assign _zz_when_ArraySlice_l166_65_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_65_5);
  assign _zz_when_ArraySlice_l166_65_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_65_5 = {3'd0, _zz_when_ArraySlice_l166_65_6};
  assign _zz_when_ArraySlice_l166_65_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_66 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_66_1);
  assign _zz_when_ArraySlice_l158_66_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_66_1 = {2'd0, _zz_when_ArraySlice_l158_66_2};
  assign _zz_when_ArraySlice_l158_66_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_66_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_66 = {1'd0, _zz_when_ArraySlice_l159_66_1};
  assign _zz_when_ArraySlice_l159_66_2 = (_zz_when_ArraySlice_l159_66_3 - _zz_when_ArraySlice_l159_66_4);
  assign _zz_when_ArraySlice_l159_66_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_66_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_66_5);
  assign _zz_when_ArraySlice_l159_66_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_66_5 = {2'd0, _zz_when_ArraySlice_l159_66_6};
  assign _zz__zz_realValue_0_66 = {1'd0, wReg};
  assign _zz__zz_realValue_0_66_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_66_1 = (_zz_realValue_0_66_2 + _zz_realValue_0_66_3);
  assign _zz_realValue_0_66_2 = {1'd0, wReg};
  assign _zz_realValue_0_66_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_66_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_66 = {1'd0, _zz_when_ArraySlice_l166_66_1};
  assign _zz_when_ArraySlice_l166_66_2 = (_zz_when_ArraySlice_l166_66_3 + _zz_when_ArraySlice_l166_66_7);
  assign _zz_when_ArraySlice_l166_66_3 = (realValue_0_66 - _zz_when_ArraySlice_l166_66_4);
  assign _zz_when_ArraySlice_l166_66_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_66_5);
  assign _zz_when_ArraySlice_l166_66_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_66_5 = {2'd0, _zz_when_ArraySlice_l166_66_6};
  assign _zz_when_ArraySlice_l166_66_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_67 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_67_1);
  assign _zz_when_ArraySlice_l158_67_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_67_1 = {2'd0, _zz_when_ArraySlice_l158_67_2};
  assign _zz_when_ArraySlice_l158_67_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_67_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_67 = {1'd0, _zz_when_ArraySlice_l159_67_1};
  assign _zz_when_ArraySlice_l159_67_2 = (_zz_when_ArraySlice_l159_67_3 - _zz_when_ArraySlice_l159_67_4);
  assign _zz_when_ArraySlice_l159_67_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_67_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_67_5);
  assign _zz_when_ArraySlice_l159_67_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_67_5 = {2'd0, _zz_when_ArraySlice_l159_67_6};
  assign _zz__zz_realValue_0_67 = {1'd0, wReg};
  assign _zz__zz_realValue_0_67_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_67_1 = (_zz_realValue_0_67_2 + _zz_realValue_0_67_3);
  assign _zz_realValue_0_67_2 = {1'd0, wReg};
  assign _zz_realValue_0_67_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_67_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_67 = {1'd0, _zz_when_ArraySlice_l166_67_1};
  assign _zz_when_ArraySlice_l166_67_2 = (_zz_when_ArraySlice_l166_67_3 + _zz_when_ArraySlice_l166_67_7);
  assign _zz_when_ArraySlice_l166_67_3 = (realValue_0_67 - _zz_when_ArraySlice_l166_67_4);
  assign _zz_when_ArraySlice_l166_67_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_67_5);
  assign _zz_when_ArraySlice_l166_67_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_67_5 = {2'd0, _zz_when_ArraySlice_l166_67_6};
  assign _zz_when_ArraySlice_l166_67_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_68 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_68_1);
  assign _zz_when_ArraySlice_l158_68_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_68_1 = {1'd0, _zz_when_ArraySlice_l158_68_2};
  assign _zz_when_ArraySlice_l158_68_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_68_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_68 = {1'd0, _zz_when_ArraySlice_l159_68_1};
  assign _zz_when_ArraySlice_l159_68_2 = (_zz_when_ArraySlice_l159_68_3 - _zz_when_ArraySlice_l159_68_4);
  assign _zz_when_ArraySlice_l159_68_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_68_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_68_5);
  assign _zz_when_ArraySlice_l159_68_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_68_5 = {1'd0, _zz_when_ArraySlice_l159_68_6};
  assign _zz__zz_realValue_0_68 = {1'd0, wReg};
  assign _zz__zz_realValue_0_68_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_68_1 = (_zz_realValue_0_68_2 + _zz_realValue_0_68_3);
  assign _zz_realValue_0_68_2 = {1'd0, wReg};
  assign _zz_realValue_0_68_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_68_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_68 = {1'd0, _zz_when_ArraySlice_l166_68_1};
  assign _zz_when_ArraySlice_l166_68_2 = (_zz_when_ArraySlice_l166_68_3 + _zz_when_ArraySlice_l166_68_7);
  assign _zz_when_ArraySlice_l166_68_3 = (realValue_0_68 - _zz_when_ArraySlice_l166_68_4);
  assign _zz_when_ArraySlice_l166_68_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_68_5);
  assign _zz_when_ArraySlice_l166_68_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_68_5 = {1'd0, _zz_when_ArraySlice_l166_68_6};
  assign _zz_when_ArraySlice_l166_68_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_69 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_69_1);
  assign _zz_when_ArraySlice_l158_69_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_69_1 = {1'd0, _zz_when_ArraySlice_l158_69_2};
  assign _zz_when_ArraySlice_l158_69_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_69_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_69 = {2'd0, _zz_when_ArraySlice_l159_69_1};
  assign _zz_when_ArraySlice_l159_69_2 = (_zz_when_ArraySlice_l159_69_3 - _zz_when_ArraySlice_l159_69_4);
  assign _zz_when_ArraySlice_l159_69_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_69_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_69_5);
  assign _zz_when_ArraySlice_l159_69_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_69_5 = {1'd0, _zz_when_ArraySlice_l159_69_6};
  assign _zz__zz_realValue_0_69 = {1'd0, wReg};
  assign _zz__zz_realValue_0_69_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_69_1 = (_zz_realValue_0_69_2 + _zz_realValue_0_69_3);
  assign _zz_realValue_0_69_2 = {1'd0, wReg};
  assign _zz_realValue_0_69_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_69_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_69 = {2'd0, _zz_when_ArraySlice_l166_69_1};
  assign _zz_when_ArraySlice_l166_69_2 = (_zz_when_ArraySlice_l166_69_3 + _zz_when_ArraySlice_l166_69_7);
  assign _zz_when_ArraySlice_l166_69_3 = (realValue_0_69 - _zz_when_ArraySlice_l166_69_4);
  assign _zz_when_ArraySlice_l166_69_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_69_5);
  assign _zz_when_ArraySlice_l166_69_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_69_5 = {1'd0, _zz_when_ArraySlice_l166_69_6};
  assign _zz_when_ArraySlice_l166_69_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_70 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_70_1);
  assign _zz_when_ArraySlice_l158_70_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_70_1 = {1'd0, _zz_when_ArraySlice_l158_70_2};
  assign _zz_when_ArraySlice_l158_70_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_70_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_70 = {2'd0, _zz_when_ArraySlice_l159_70_1};
  assign _zz_when_ArraySlice_l159_70_2 = (_zz_when_ArraySlice_l159_70_3 - _zz_when_ArraySlice_l159_70_4);
  assign _zz_when_ArraySlice_l159_70_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_70_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_70_5);
  assign _zz_when_ArraySlice_l159_70_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_70_5 = {1'd0, _zz_when_ArraySlice_l159_70_6};
  assign _zz__zz_realValue_0_70 = {1'd0, wReg};
  assign _zz__zz_realValue_0_70_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_70_1 = (_zz_realValue_0_70_2 + _zz_realValue_0_70_3);
  assign _zz_realValue_0_70_2 = {1'd0, wReg};
  assign _zz_realValue_0_70_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_70_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_70 = {2'd0, _zz_when_ArraySlice_l166_70_1};
  assign _zz_when_ArraySlice_l166_70_2 = (_zz_when_ArraySlice_l166_70_3 + _zz_when_ArraySlice_l166_70_7);
  assign _zz_when_ArraySlice_l166_70_3 = (realValue_0_70 - _zz_when_ArraySlice_l166_70_4);
  assign _zz_when_ArraySlice_l166_70_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_70_5);
  assign _zz_when_ArraySlice_l166_70_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_70_5 = {1'd0, _zz_when_ArraySlice_l166_70_6};
  assign _zz_when_ArraySlice_l166_70_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_71 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_71_1);
  assign _zz_when_ArraySlice_l158_71_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_71_1 = {1'd0, _zz_when_ArraySlice_l158_71_2};
  assign _zz_when_ArraySlice_l158_71_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_71_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_71 = {3'd0, _zz_when_ArraySlice_l159_71_1};
  assign _zz_when_ArraySlice_l159_71_2 = (_zz_when_ArraySlice_l159_71_3 - _zz_when_ArraySlice_l159_71_4);
  assign _zz_when_ArraySlice_l159_71_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_71_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_71_5);
  assign _zz_when_ArraySlice_l159_71_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_71_5 = {1'd0, _zz_when_ArraySlice_l159_71_6};
  assign _zz__zz_realValue_0_71 = {1'd0, wReg};
  assign _zz__zz_realValue_0_71_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_71_1 = (_zz_realValue_0_71_2 + _zz_realValue_0_71_3);
  assign _zz_realValue_0_71_2 = {1'd0, wReg};
  assign _zz_realValue_0_71_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_71_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_71 = {3'd0, _zz_when_ArraySlice_l166_71_1};
  assign _zz_when_ArraySlice_l166_71_2 = (_zz_when_ArraySlice_l166_71_3 + _zz_when_ArraySlice_l166_71_7);
  assign _zz_when_ArraySlice_l166_71_3 = (realValue_0_71 - _zz_when_ArraySlice_l166_71_4);
  assign _zz_when_ArraySlice_l166_71_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_71_5);
  assign _zz_when_ArraySlice_l166_71_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_71_5 = {1'd0, _zz_when_ArraySlice_l166_71_6};
  assign _zz_when_ArraySlice_l166_71_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_2_2 = (_zz_when_ArraySlice_l428_2_3 + _zz_when_ArraySlice_l428_2_7);
  assign _zz_when_ArraySlice_l428_2_3 = (_zz_when_ArraySlice_l428_2_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l428_2_5);
  assign _zz_when_ArraySlice_l428_2_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_2_5 = {1'd0, _zz_when_ArraySlice_l428_2_6};
  assign _zz_when_ArraySlice_l428_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l428_2_7 = {2'd0, _zz_when_ArraySlice_l428_2_8};
  assign _zz_when_ArraySlice_l431_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_2_2 = (_zz_when_ArraySlice_l431_2_3 + 8'h01);
  assign _zz_when_ArraySlice_l431_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l431_2_4);
  assign _zz_when_ArraySlice_l431_2_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_2_4 = {1'd0, _zz_when_ArraySlice_l431_2_5};
  assign _zz_selectReadFifo_2_11 = (selectReadFifo_2 + _zz_selectReadFifo_2_12);
  assign _zz_selectReadFifo_2_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_12 = {1'd0, _zz_selectReadFifo_2_13};
  assign _zz_when_ArraySlice_l438_2 = (_zz_when_ArraySlice_l438_2_1 % aReg);
  assign _zz_when_ArraySlice_l438_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_2_2 = (_zz_when_ArraySlice_l449_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l449_2_1 = {5'd0, _zz_when_ArraySlice_l449_2_2};
  assign _zz_when_ArraySlice_l449_2_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_8 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_8_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_8_1 = (_zz_realValue1_0_8_2 + _zz_realValue1_0_8_3);
  assign _zz_realValue1_0_8_2 = {1'd0, hReg};
  assign _zz_realValue1_0_8_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l450_2_1 = {1'd0, _zz_when_ArraySlice_l450_2_2};
  assign _zz_when_ArraySlice_l450_2_3 = (realValue1_0_8 / aReg);
  assign _zz_selectReadFifo_2_14 = (selectReadFifo_2 - _zz_selectReadFifo_2_15);
  assign _zz_selectReadFifo_2_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_72 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_72_1);
  assign _zz_when_ArraySlice_l158_72_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_72_1 = {4'd0, _zz_when_ArraySlice_l158_72_2};
  assign _zz_when_ArraySlice_l158_72_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_72 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_72_1 = (_zz_when_ArraySlice_l159_72_2 - _zz_when_ArraySlice_l159_72_3);
  assign _zz_when_ArraySlice_l159_72_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_72_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_72_4);
  assign _zz_when_ArraySlice_l159_72_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_72_4 = {4'd0, _zz_when_ArraySlice_l159_72_5};
  assign _zz__zz_realValue_0_72 = {1'd0, wReg};
  assign _zz__zz_realValue_0_72_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_72_1 = (_zz_realValue_0_72_2 + _zz_realValue_0_72_3);
  assign _zz_realValue_0_72_2 = {1'd0, wReg};
  assign _zz_realValue_0_72_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_72 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_72_1 = (_zz_when_ArraySlice_l166_72_2 + _zz_when_ArraySlice_l166_72_6);
  assign _zz_when_ArraySlice_l166_72_2 = (realValue_0_72 - _zz_when_ArraySlice_l166_72_3);
  assign _zz_when_ArraySlice_l166_72_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_72_4);
  assign _zz_when_ArraySlice_l166_72_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_72_4 = {4'd0, _zz_when_ArraySlice_l166_72_5};
  assign _zz_when_ArraySlice_l166_72_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_73 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_73_1);
  assign _zz_when_ArraySlice_l158_73_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_73_1 = {3'd0, _zz_when_ArraySlice_l158_73_2};
  assign _zz_when_ArraySlice_l158_73_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_73_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_73 = {1'd0, _zz_when_ArraySlice_l159_73_1};
  assign _zz_when_ArraySlice_l159_73_2 = (_zz_when_ArraySlice_l159_73_3 - _zz_when_ArraySlice_l159_73_4);
  assign _zz_when_ArraySlice_l159_73_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_73_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_73_5);
  assign _zz_when_ArraySlice_l159_73_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_73_5 = {3'd0, _zz_when_ArraySlice_l159_73_6};
  assign _zz__zz_realValue_0_73 = {1'd0, wReg};
  assign _zz__zz_realValue_0_73_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_73_1 = (_zz_realValue_0_73_2 + _zz_realValue_0_73_3);
  assign _zz_realValue_0_73_2 = {1'd0, wReg};
  assign _zz_realValue_0_73_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_73_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_73 = {1'd0, _zz_when_ArraySlice_l166_73_1};
  assign _zz_when_ArraySlice_l166_73_2 = (_zz_when_ArraySlice_l166_73_3 + _zz_when_ArraySlice_l166_73_7);
  assign _zz_when_ArraySlice_l166_73_3 = (realValue_0_73 - _zz_when_ArraySlice_l166_73_4);
  assign _zz_when_ArraySlice_l166_73_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_73_5);
  assign _zz_when_ArraySlice_l166_73_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_73_5 = {3'd0, _zz_when_ArraySlice_l166_73_6};
  assign _zz_when_ArraySlice_l166_73_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_74 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_74_1);
  assign _zz_when_ArraySlice_l158_74_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_74_1 = {2'd0, _zz_when_ArraySlice_l158_74_2};
  assign _zz_when_ArraySlice_l158_74_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_74_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_74 = {1'd0, _zz_when_ArraySlice_l159_74_1};
  assign _zz_when_ArraySlice_l159_74_2 = (_zz_when_ArraySlice_l159_74_3 - _zz_when_ArraySlice_l159_74_4);
  assign _zz_when_ArraySlice_l159_74_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_74_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_74_5);
  assign _zz_when_ArraySlice_l159_74_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_74_5 = {2'd0, _zz_when_ArraySlice_l159_74_6};
  assign _zz__zz_realValue_0_74 = {1'd0, wReg};
  assign _zz__zz_realValue_0_74_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_74_1 = (_zz_realValue_0_74_2 + _zz_realValue_0_74_3);
  assign _zz_realValue_0_74_2 = {1'd0, wReg};
  assign _zz_realValue_0_74_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_74_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_74 = {1'd0, _zz_when_ArraySlice_l166_74_1};
  assign _zz_when_ArraySlice_l166_74_2 = (_zz_when_ArraySlice_l166_74_3 + _zz_when_ArraySlice_l166_74_7);
  assign _zz_when_ArraySlice_l166_74_3 = (realValue_0_74 - _zz_when_ArraySlice_l166_74_4);
  assign _zz_when_ArraySlice_l166_74_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_74_5);
  assign _zz_when_ArraySlice_l166_74_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_74_5 = {2'd0, _zz_when_ArraySlice_l166_74_6};
  assign _zz_when_ArraySlice_l166_74_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_75 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_75_1);
  assign _zz_when_ArraySlice_l158_75_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_75_1 = {2'd0, _zz_when_ArraySlice_l158_75_2};
  assign _zz_when_ArraySlice_l158_75_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_75_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_75 = {1'd0, _zz_when_ArraySlice_l159_75_1};
  assign _zz_when_ArraySlice_l159_75_2 = (_zz_when_ArraySlice_l159_75_3 - _zz_when_ArraySlice_l159_75_4);
  assign _zz_when_ArraySlice_l159_75_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_75_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_75_5);
  assign _zz_when_ArraySlice_l159_75_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_75_5 = {2'd0, _zz_when_ArraySlice_l159_75_6};
  assign _zz__zz_realValue_0_75 = {1'd0, wReg};
  assign _zz__zz_realValue_0_75_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_75_1 = (_zz_realValue_0_75_2 + _zz_realValue_0_75_3);
  assign _zz_realValue_0_75_2 = {1'd0, wReg};
  assign _zz_realValue_0_75_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_75_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_75 = {1'd0, _zz_when_ArraySlice_l166_75_1};
  assign _zz_when_ArraySlice_l166_75_2 = (_zz_when_ArraySlice_l166_75_3 + _zz_when_ArraySlice_l166_75_7);
  assign _zz_when_ArraySlice_l166_75_3 = (realValue_0_75 - _zz_when_ArraySlice_l166_75_4);
  assign _zz_when_ArraySlice_l166_75_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_75_5);
  assign _zz_when_ArraySlice_l166_75_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_75_5 = {2'd0, _zz_when_ArraySlice_l166_75_6};
  assign _zz_when_ArraySlice_l166_75_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_76 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_76_1);
  assign _zz_when_ArraySlice_l158_76_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_76_1 = {1'd0, _zz_when_ArraySlice_l158_76_2};
  assign _zz_when_ArraySlice_l158_76_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_76_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_76 = {1'd0, _zz_when_ArraySlice_l159_76_1};
  assign _zz_when_ArraySlice_l159_76_2 = (_zz_when_ArraySlice_l159_76_3 - _zz_when_ArraySlice_l159_76_4);
  assign _zz_when_ArraySlice_l159_76_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_76_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_76_5);
  assign _zz_when_ArraySlice_l159_76_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_76_5 = {1'd0, _zz_when_ArraySlice_l159_76_6};
  assign _zz__zz_realValue_0_76 = {1'd0, wReg};
  assign _zz__zz_realValue_0_76_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_76_1 = (_zz_realValue_0_76_2 + _zz_realValue_0_76_3);
  assign _zz_realValue_0_76_2 = {1'd0, wReg};
  assign _zz_realValue_0_76_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_76_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_76 = {1'd0, _zz_when_ArraySlice_l166_76_1};
  assign _zz_when_ArraySlice_l166_76_2 = (_zz_when_ArraySlice_l166_76_3 + _zz_when_ArraySlice_l166_76_7);
  assign _zz_when_ArraySlice_l166_76_3 = (realValue_0_76 - _zz_when_ArraySlice_l166_76_4);
  assign _zz_when_ArraySlice_l166_76_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_76_5);
  assign _zz_when_ArraySlice_l166_76_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_76_5 = {1'd0, _zz_when_ArraySlice_l166_76_6};
  assign _zz_when_ArraySlice_l166_76_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_77 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_77_1);
  assign _zz_when_ArraySlice_l158_77_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_77_1 = {1'd0, _zz_when_ArraySlice_l158_77_2};
  assign _zz_when_ArraySlice_l158_77_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_77_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_77 = {2'd0, _zz_when_ArraySlice_l159_77_1};
  assign _zz_when_ArraySlice_l159_77_2 = (_zz_when_ArraySlice_l159_77_3 - _zz_when_ArraySlice_l159_77_4);
  assign _zz_when_ArraySlice_l159_77_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_77_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_77_5);
  assign _zz_when_ArraySlice_l159_77_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_77_5 = {1'd0, _zz_when_ArraySlice_l159_77_6};
  assign _zz__zz_realValue_0_77 = {1'd0, wReg};
  assign _zz__zz_realValue_0_77_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_77_1 = (_zz_realValue_0_77_2 + _zz_realValue_0_77_3);
  assign _zz_realValue_0_77_2 = {1'd0, wReg};
  assign _zz_realValue_0_77_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_77_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_77 = {2'd0, _zz_when_ArraySlice_l166_77_1};
  assign _zz_when_ArraySlice_l166_77_2 = (_zz_when_ArraySlice_l166_77_3 + _zz_when_ArraySlice_l166_77_7);
  assign _zz_when_ArraySlice_l166_77_3 = (realValue_0_77 - _zz_when_ArraySlice_l166_77_4);
  assign _zz_when_ArraySlice_l166_77_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_77_5);
  assign _zz_when_ArraySlice_l166_77_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_77_5 = {1'd0, _zz_when_ArraySlice_l166_77_6};
  assign _zz_when_ArraySlice_l166_77_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_78 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_78_1);
  assign _zz_when_ArraySlice_l158_78_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_78_1 = {1'd0, _zz_when_ArraySlice_l158_78_2};
  assign _zz_when_ArraySlice_l158_78_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_78_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_78 = {2'd0, _zz_when_ArraySlice_l159_78_1};
  assign _zz_when_ArraySlice_l159_78_2 = (_zz_when_ArraySlice_l159_78_3 - _zz_when_ArraySlice_l159_78_4);
  assign _zz_when_ArraySlice_l159_78_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_78_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_78_5);
  assign _zz_when_ArraySlice_l159_78_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_78_5 = {1'd0, _zz_when_ArraySlice_l159_78_6};
  assign _zz__zz_realValue_0_78 = {1'd0, wReg};
  assign _zz__zz_realValue_0_78_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_78_1 = (_zz_realValue_0_78_2 + _zz_realValue_0_78_3);
  assign _zz_realValue_0_78_2 = {1'd0, wReg};
  assign _zz_realValue_0_78_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_78_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_78 = {2'd0, _zz_when_ArraySlice_l166_78_1};
  assign _zz_when_ArraySlice_l166_78_2 = (_zz_when_ArraySlice_l166_78_3 + _zz_when_ArraySlice_l166_78_7);
  assign _zz_when_ArraySlice_l166_78_3 = (realValue_0_78 - _zz_when_ArraySlice_l166_78_4);
  assign _zz_when_ArraySlice_l166_78_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_78_5);
  assign _zz_when_ArraySlice_l166_78_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_78_5 = {1'd0, _zz_when_ArraySlice_l166_78_6};
  assign _zz_when_ArraySlice_l166_78_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_79 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_79_1);
  assign _zz_when_ArraySlice_l158_79_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_79_1 = {1'd0, _zz_when_ArraySlice_l158_79_2};
  assign _zz_when_ArraySlice_l158_79_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_79_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_79 = {3'd0, _zz_when_ArraySlice_l159_79_1};
  assign _zz_when_ArraySlice_l159_79_2 = (_zz_when_ArraySlice_l159_79_3 - _zz_when_ArraySlice_l159_79_4);
  assign _zz_when_ArraySlice_l159_79_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_79_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_79_5);
  assign _zz_when_ArraySlice_l159_79_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_79_5 = {1'd0, _zz_when_ArraySlice_l159_79_6};
  assign _zz__zz_realValue_0_79 = {1'd0, wReg};
  assign _zz__zz_realValue_0_79_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_79_1 = (_zz_realValue_0_79_2 + _zz_realValue_0_79_3);
  assign _zz_realValue_0_79_2 = {1'd0, wReg};
  assign _zz_realValue_0_79_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_79_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_79 = {3'd0, _zz_when_ArraySlice_l166_79_1};
  assign _zz_when_ArraySlice_l166_79_2 = (_zz_when_ArraySlice_l166_79_3 + _zz_when_ArraySlice_l166_79_7);
  assign _zz_when_ArraySlice_l166_79_3 = (realValue_0_79 - _zz_when_ArraySlice_l166_79_4);
  assign _zz_when_ArraySlice_l166_79_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_79_5);
  assign _zz_when_ArraySlice_l166_79_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_79_5 = {1'd0, _zz_when_ArraySlice_l166_79_6};
  assign _zz_when_ArraySlice_l166_79_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_2 = (_zz_when_ArraySlice_l461_2_1 % aReg);
  assign _zz_when_ArraySlice_l461_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l447_2_3);
  assign _zz_when_ArraySlice_l447_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l447_2_3 = {2'd0, _zz_when_ArraySlice_l447_2_4};
  assign _zz_when_ArraySlice_l468_2_2 = (_zz_when_ArraySlice_l468_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l468_2_1 = {5'd0, _zz_when_ArraySlice_l468_2_2};
  assign _zz_when_ArraySlice_l468_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_3_1 = (selectReadFifo_3 + _zz_when_ArraySlice_l376_3_2);
  assign _zz_when_ArraySlice_l376_3_3 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l376_3_2 = {2'd0, _zz_when_ArraySlice_l376_3_3};
  assign _zz_when_ArraySlice_l376_3_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l377_3_4);
  assign _zz_when_ArraySlice_l377_3_2 = _zz_when_ArraySlice_l377_3_3[6:0];
  assign _zz_when_ArraySlice_l377_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l377_3_4 = {2'd0, _zz_when_ArraySlice_l377_3_5};
  assign _zz__zz_outputStreamArrayData_3_valid_1 = (bReg * 2'b11);
  assign _zz__zz_outputStreamArrayData_3_valid = {2'd0, _zz__zz_outputStreamArrayData_3_valid_1};
  assign _zz__zz_6 = _zz_outputStreamArrayData_3_valid[6:0];
  assign _zz_outputStreamArrayData_3_valid_3 = _zz_outputStreamArrayData_3_valid[6:0];
  assign _zz_outputStreamArrayData_3_payload_1 = _zz_outputStreamArrayData_3_valid[6:0];
  assign _zz_when_ArraySlice_l383_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l383_3_4);
  assign _zz_when_ArraySlice_l383_3_2 = _zz_when_ArraySlice_l383_3_3[6:0];
  assign _zz_when_ArraySlice_l383_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l383_3_4 = {2'd0, _zz_when_ArraySlice_l383_3_5};
  assign _zz_when_ArraySlice_l384_3_1 = (_zz_when_ArraySlice_l384_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l384_3 = {5'd0, _zz_when_ArraySlice_l384_3_1};
  assign _zz_when_ArraySlice_l384_3_2 = (bReg * aReg);
  assign _zz_selectReadFifo_3 = (selectReadFifo_3 - _zz_selectReadFifo_3_1);
  assign _zz_selectReadFifo_3_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_3 = (_zz_when_ArraySlice_l387_3_1 % aReg);
  assign _zz_when_ArraySlice_l387_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l392_3_4);
  assign _zz_when_ArraySlice_l392_3_2 = _zz_when_ArraySlice_l392_3_3[6:0];
  assign _zz_when_ArraySlice_l392_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l392_3_4 = {2'd0, _zz_when_ArraySlice_l392_3_5};
  assign _zz_when_ArraySlice_l393_3_1 = (_zz_when_ArraySlice_l393_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l393_3 = {5'd0, _zz_when_ArraySlice_l393_3_1};
  assign _zz_when_ArraySlice_l393_3_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_9 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_9_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_9_1 = (_zz_realValue1_0_9_2 + _zz_realValue1_0_9_3);
  assign _zz_realValue1_0_9_2 = {1'd0, hReg};
  assign _zz_realValue1_0_9_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l395_3 = {1'd0, _zz_when_ArraySlice_l395_3_1};
  assign _zz_when_ArraySlice_l395_3_2 = (realValue1_0_9 / aReg);
  assign _zz_selectReadFifo_3_2 = (selectReadFifo_3 - _zz_selectReadFifo_3_3);
  assign _zz_selectReadFifo_3_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_3_5 = 1'b1;
  assign _zz_selectReadFifo_3_4 = {7'd0, _zz_selectReadFifo_3_5};
  assign _zz_when_ArraySlice_l158_80 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_80_1);
  assign _zz_when_ArraySlice_l158_80_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_80_1 = {4'd0, _zz_when_ArraySlice_l158_80_2};
  assign _zz_when_ArraySlice_l158_80_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_80 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_80_1 = (_zz_when_ArraySlice_l159_80_2 - _zz_when_ArraySlice_l159_80_3);
  assign _zz_when_ArraySlice_l159_80_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_80_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_80_4);
  assign _zz_when_ArraySlice_l159_80_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_80_4 = {4'd0, _zz_when_ArraySlice_l159_80_5};
  assign _zz__zz_realValue_0_80 = {1'd0, wReg};
  assign _zz__zz_realValue_0_80_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_80_1 = (_zz_realValue_0_80_2 + _zz_realValue_0_80_3);
  assign _zz_realValue_0_80_2 = {1'd0, wReg};
  assign _zz_realValue_0_80_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_80 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_80_1 = (_zz_when_ArraySlice_l166_80_2 + _zz_when_ArraySlice_l166_80_6);
  assign _zz_when_ArraySlice_l166_80_2 = (realValue_0_80 - _zz_when_ArraySlice_l166_80_3);
  assign _zz_when_ArraySlice_l166_80_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_80_4);
  assign _zz_when_ArraySlice_l166_80_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_80_4 = {4'd0, _zz_when_ArraySlice_l166_80_5};
  assign _zz_when_ArraySlice_l166_80_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_81 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_81_1);
  assign _zz_when_ArraySlice_l158_81_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_81_1 = {3'd0, _zz_when_ArraySlice_l158_81_2};
  assign _zz_when_ArraySlice_l158_81_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_81_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_81 = {1'd0, _zz_when_ArraySlice_l159_81_1};
  assign _zz_when_ArraySlice_l159_81_2 = (_zz_when_ArraySlice_l159_81_3 - _zz_when_ArraySlice_l159_81_4);
  assign _zz_when_ArraySlice_l159_81_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_81_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_81_5);
  assign _zz_when_ArraySlice_l159_81_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_81_5 = {3'd0, _zz_when_ArraySlice_l159_81_6};
  assign _zz__zz_realValue_0_81 = {1'd0, wReg};
  assign _zz__zz_realValue_0_81_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_81_1 = (_zz_realValue_0_81_2 + _zz_realValue_0_81_3);
  assign _zz_realValue_0_81_2 = {1'd0, wReg};
  assign _zz_realValue_0_81_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_81_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_81 = {1'd0, _zz_when_ArraySlice_l166_81_1};
  assign _zz_when_ArraySlice_l166_81_2 = (_zz_when_ArraySlice_l166_81_3 + _zz_when_ArraySlice_l166_81_7);
  assign _zz_when_ArraySlice_l166_81_3 = (realValue_0_81 - _zz_when_ArraySlice_l166_81_4);
  assign _zz_when_ArraySlice_l166_81_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_81_5);
  assign _zz_when_ArraySlice_l166_81_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_81_5 = {3'd0, _zz_when_ArraySlice_l166_81_6};
  assign _zz_when_ArraySlice_l166_81_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_82 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_82_1);
  assign _zz_when_ArraySlice_l158_82_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_82_1 = {2'd0, _zz_when_ArraySlice_l158_82_2};
  assign _zz_when_ArraySlice_l158_82_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_82_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_82 = {1'd0, _zz_when_ArraySlice_l159_82_1};
  assign _zz_when_ArraySlice_l159_82_2 = (_zz_when_ArraySlice_l159_82_3 - _zz_when_ArraySlice_l159_82_4);
  assign _zz_when_ArraySlice_l159_82_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_82_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_82_5);
  assign _zz_when_ArraySlice_l159_82_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_82_5 = {2'd0, _zz_when_ArraySlice_l159_82_6};
  assign _zz__zz_realValue_0_82 = {1'd0, wReg};
  assign _zz__zz_realValue_0_82_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_82_1 = (_zz_realValue_0_82_2 + _zz_realValue_0_82_3);
  assign _zz_realValue_0_82_2 = {1'd0, wReg};
  assign _zz_realValue_0_82_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_82_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_82 = {1'd0, _zz_when_ArraySlice_l166_82_1};
  assign _zz_when_ArraySlice_l166_82_2 = (_zz_when_ArraySlice_l166_82_3 + _zz_when_ArraySlice_l166_82_7);
  assign _zz_when_ArraySlice_l166_82_3 = (realValue_0_82 - _zz_when_ArraySlice_l166_82_4);
  assign _zz_when_ArraySlice_l166_82_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_82_5);
  assign _zz_when_ArraySlice_l166_82_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_82_5 = {2'd0, _zz_when_ArraySlice_l166_82_6};
  assign _zz_when_ArraySlice_l166_82_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_83 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_83_1);
  assign _zz_when_ArraySlice_l158_83_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_83_1 = {2'd0, _zz_when_ArraySlice_l158_83_2};
  assign _zz_when_ArraySlice_l158_83_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_83_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_83 = {1'd0, _zz_when_ArraySlice_l159_83_1};
  assign _zz_when_ArraySlice_l159_83_2 = (_zz_when_ArraySlice_l159_83_3 - _zz_when_ArraySlice_l159_83_4);
  assign _zz_when_ArraySlice_l159_83_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_83_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_83_5);
  assign _zz_when_ArraySlice_l159_83_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_83_5 = {2'd0, _zz_when_ArraySlice_l159_83_6};
  assign _zz__zz_realValue_0_83 = {1'd0, wReg};
  assign _zz__zz_realValue_0_83_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_83_1 = (_zz_realValue_0_83_2 + _zz_realValue_0_83_3);
  assign _zz_realValue_0_83_2 = {1'd0, wReg};
  assign _zz_realValue_0_83_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_83_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_83 = {1'd0, _zz_when_ArraySlice_l166_83_1};
  assign _zz_when_ArraySlice_l166_83_2 = (_zz_when_ArraySlice_l166_83_3 + _zz_when_ArraySlice_l166_83_7);
  assign _zz_when_ArraySlice_l166_83_3 = (realValue_0_83 - _zz_when_ArraySlice_l166_83_4);
  assign _zz_when_ArraySlice_l166_83_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_83_5);
  assign _zz_when_ArraySlice_l166_83_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_83_5 = {2'd0, _zz_when_ArraySlice_l166_83_6};
  assign _zz_when_ArraySlice_l166_83_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_84 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_84_1);
  assign _zz_when_ArraySlice_l158_84_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_84_1 = {1'd0, _zz_when_ArraySlice_l158_84_2};
  assign _zz_when_ArraySlice_l158_84_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_84_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_84 = {1'd0, _zz_when_ArraySlice_l159_84_1};
  assign _zz_when_ArraySlice_l159_84_2 = (_zz_when_ArraySlice_l159_84_3 - _zz_when_ArraySlice_l159_84_4);
  assign _zz_when_ArraySlice_l159_84_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_84_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_84_5);
  assign _zz_when_ArraySlice_l159_84_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_84_5 = {1'd0, _zz_when_ArraySlice_l159_84_6};
  assign _zz__zz_realValue_0_84 = {1'd0, wReg};
  assign _zz__zz_realValue_0_84_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_84_1 = (_zz_realValue_0_84_2 + _zz_realValue_0_84_3);
  assign _zz_realValue_0_84_2 = {1'd0, wReg};
  assign _zz_realValue_0_84_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_84_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_84 = {1'd0, _zz_when_ArraySlice_l166_84_1};
  assign _zz_when_ArraySlice_l166_84_2 = (_zz_when_ArraySlice_l166_84_3 + _zz_when_ArraySlice_l166_84_7);
  assign _zz_when_ArraySlice_l166_84_3 = (realValue_0_84 - _zz_when_ArraySlice_l166_84_4);
  assign _zz_when_ArraySlice_l166_84_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_84_5);
  assign _zz_when_ArraySlice_l166_84_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_84_5 = {1'd0, _zz_when_ArraySlice_l166_84_6};
  assign _zz_when_ArraySlice_l166_84_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_85 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_85_1);
  assign _zz_when_ArraySlice_l158_85_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_85_1 = {1'd0, _zz_when_ArraySlice_l158_85_2};
  assign _zz_when_ArraySlice_l158_85_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_85_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_85 = {2'd0, _zz_when_ArraySlice_l159_85_1};
  assign _zz_when_ArraySlice_l159_85_2 = (_zz_when_ArraySlice_l159_85_3 - _zz_when_ArraySlice_l159_85_4);
  assign _zz_when_ArraySlice_l159_85_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_85_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_85_5);
  assign _zz_when_ArraySlice_l159_85_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_85_5 = {1'd0, _zz_when_ArraySlice_l159_85_6};
  assign _zz__zz_realValue_0_85 = {1'd0, wReg};
  assign _zz__zz_realValue_0_85_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_85_1 = (_zz_realValue_0_85_2 + _zz_realValue_0_85_3);
  assign _zz_realValue_0_85_2 = {1'd0, wReg};
  assign _zz_realValue_0_85_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_85_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_85 = {2'd0, _zz_when_ArraySlice_l166_85_1};
  assign _zz_when_ArraySlice_l166_85_2 = (_zz_when_ArraySlice_l166_85_3 + _zz_when_ArraySlice_l166_85_7);
  assign _zz_when_ArraySlice_l166_85_3 = (realValue_0_85 - _zz_when_ArraySlice_l166_85_4);
  assign _zz_when_ArraySlice_l166_85_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_85_5);
  assign _zz_when_ArraySlice_l166_85_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_85_5 = {1'd0, _zz_when_ArraySlice_l166_85_6};
  assign _zz_when_ArraySlice_l166_85_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_86 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_86_1);
  assign _zz_when_ArraySlice_l158_86_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_86_1 = {1'd0, _zz_when_ArraySlice_l158_86_2};
  assign _zz_when_ArraySlice_l158_86_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_86_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_86 = {2'd0, _zz_when_ArraySlice_l159_86_1};
  assign _zz_when_ArraySlice_l159_86_2 = (_zz_when_ArraySlice_l159_86_3 - _zz_when_ArraySlice_l159_86_4);
  assign _zz_when_ArraySlice_l159_86_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_86_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_86_5);
  assign _zz_when_ArraySlice_l159_86_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_86_5 = {1'd0, _zz_when_ArraySlice_l159_86_6};
  assign _zz__zz_realValue_0_86 = {1'd0, wReg};
  assign _zz__zz_realValue_0_86_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_86_1 = (_zz_realValue_0_86_2 + _zz_realValue_0_86_3);
  assign _zz_realValue_0_86_2 = {1'd0, wReg};
  assign _zz_realValue_0_86_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_86_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_86 = {2'd0, _zz_when_ArraySlice_l166_86_1};
  assign _zz_when_ArraySlice_l166_86_2 = (_zz_when_ArraySlice_l166_86_3 + _zz_when_ArraySlice_l166_86_7);
  assign _zz_when_ArraySlice_l166_86_3 = (realValue_0_86 - _zz_when_ArraySlice_l166_86_4);
  assign _zz_when_ArraySlice_l166_86_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_86_5);
  assign _zz_when_ArraySlice_l166_86_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_86_5 = {1'd0, _zz_when_ArraySlice_l166_86_6};
  assign _zz_when_ArraySlice_l166_86_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_87 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_87_1);
  assign _zz_when_ArraySlice_l158_87_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_87_1 = {1'd0, _zz_when_ArraySlice_l158_87_2};
  assign _zz_when_ArraySlice_l158_87_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_87_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_87 = {3'd0, _zz_when_ArraySlice_l159_87_1};
  assign _zz_when_ArraySlice_l159_87_2 = (_zz_when_ArraySlice_l159_87_3 - _zz_when_ArraySlice_l159_87_4);
  assign _zz_when_ArraySlice_l159_87_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_87_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_87_5);
  assign _zz_when_ArraySlice_l159_87_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_87_5 = {1'd0, _zz_when_ArraySlice_l159_87_6};
  assign _zz__zz_realValue_0_87 = {1'd0, wReg};
  assign _zz__zz_realValue_0_87_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_87_1 = (_zz_realValue_0_87_2 + _zz_realValue_0_87_3);
  assign _zz_realValue_0_87_2 = {1'd0, wReg};
  assign _zz_realValue_0_87_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_87_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_87 = {3'd0, _zz_when_ArraySlice_l166_87_1};
  assign _zz_when_ArraySlice_l166_87_2 = (_zz_when_ArraySlice_l166_87_3 + _zz_when_ArraySlice_l166_87_7);
  assign _zz_when_ArraySlice_l166_87_3 = (realValue_0_87 - _zz_when_ArraySlice_l166_87_4);
  assign _zz_when_ArraySlice_l166_87_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_87_5);
  assign _zz_when_ArraySlice_l166_87_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_87_5 = {1'd0, _zz_when_ArraySlice_l166_87_6};
  assign _zz_when_ArraySlice_l166_87_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_3_2 = (_zz_when_ArraySlice_l403_3_3 + _zz_when_ArraySlice_l403_3_7);
  assign _zz_when_ArraySlice_l403_3_3 = (_zz_when_ArraySlice_l403_3_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l403_3_5);
  assign _zz_when_ArraySlice_l403_3_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_3_5 = {1'd0, _zz_when_ArraySlice_l403_3_6};
  assign _zz_when_ArraySlice_l403_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l403_3_7 = {2'd0, _zz_when_ArraySlice_l403_3_8};
  assign _zz_when_ArraySlice_l406_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_3_2 = (_zz_when_ArraySlice_l406_3_3 + 8'h01);
  assign _zz_when_ArraySlice_l406_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l406_3_4);
  assign _zz_when_ArraySlice_l406_3_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_3_4 = {1'd0, _zz_when_ArraySlice_l406_3_5};
  assign _zz_selectReadFifo_3_6 = (selectReadFifo_3 + _zz_selectReadFifo_3_7);
  assign _zz_selectReadFifo_3_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_7 = {1'd0, _zz_selectReadFifo_3_8};
  assign _zz_when_ArraySlice_l413_3 = (_zz_when_ArraySlice_l413_3_1 % aReg);
  assign _zz_when_ArraySlice_l413_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l417_3_4);
  assign _zz_when_ArraySlice_l417_3_2 = _zz_when_ArraySlice_l417_3_3[6:0];
  assign _zz_when_ArraySlice_l417_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l417_3_4 = {2'd0, _zz_when_ArraySlice_l417_3_5};
  assign _zz_when_ArraySlice_l418_3_2 = (_zz_when_ArraySlice_l418_3_3 - _zz_when_ArraySlice_l418_3_4);
  assign _zz_when_ArraySlice_l418_3_1 = {5'd0, _zz_when_ArraySlice_l418_3_2};
  assign _zz_when_ArraySlice_l418_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l418_3_4 = {7'd0, _zz_when_ArraySlice_l418_3_5};
  assign _zz__zz_realValue1_0_10 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_10_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_10_1 = (_zz_realValue1_0_10_2 + _zz_realValue1_0_10_3);
  assign _zz_realValue1_0_10_2 = {1'd0, hReg};
  assign _zz_realValue1_0_10_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l420_3 = {1'd0, _zz_when_ArraySlice_l420_3_1};
  assign _zz_when_ArraySlice_l420_3_2 = (realValue1_0_10 / aReg);
  assign _zz_selectReadFifo_3_9 = (selectReadFifo_3 - _zz_selectReadFifo_3_10);
  assign _zz_selectReadFifo_3_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_88 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_88_1);
  assign _zz_when_ArraySlice_l158_88_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_88_1 = {4'd0, _zz_when_ArraySlice_l158_88_2};
  assign _zz_when_ArraySlice_l158_88_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_88 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_88_1 = (_zz_when_ArraySlice_l159_88_2 - _zz_when_ArraySlice_l159_88_3);
  assign _zz_when_ArraySlice_l159_88_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_88_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_88_4);
  assign _zz_when_ArraySlice_l159_88_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_88_4 = {4'd0, _zz_when_ArraySlice_l159_88_5};
  assign _zz__zz_realValue_0_88 = {1'd0, wReg};
  assign _zz__zz_realValue_0_88_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_88_1 = (_zz_realValue_0_88_2 + _zz_realValue_0_88_3);
  assign _zz_realValue_0_88_2 = {1'd0, wReg};
  assign _zz_realValue_0_88_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_88 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_88_1 = (_zz_when_ArraySlice_l166_88_2 + _zz_when_ArraySlice_l166_88_6);
  assign _zz_when_ArraySlice_l166_88_2 = (realValue_0_88 - _zz_when_ArraySlice_l166_88_3);
  assign _zz_when_ArraySlice_l166_88_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_88_4);
  assign _zz_when_ArraySlice_l166_88_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_88_4 = {4'd0, _zz_when_ArraySlice_l166_88_5};
  assign _zz_when_ArraySlice_l166_88_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_89 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_89_1);
  assign _zz_when_ArraySlice_l158_89_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_89_1 = {3'd0, _zz_when_ArraySlice_l158_89_2};
  assign _zz_when_ArraySlice_l158_89_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_89_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_89 = {1'd0, _zz_when_ArraySlice_l159_89_1};
  assign _zz_when_ArraySlice_l159_89_2 = (_zz_when_ArraySlice_l159_89_3 - _zz_when_ArraySlice_l159_89_4);
  assign _zz_when_ArraySlice_l159_89_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_89_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_89_5);
  assign _zz_when_ArraySlice_l159_89_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_89_5 = {3'd0, _zz_when_ArraySlice_l159_89_6};
  assign _zz__zz_realValue_0_89 = {1'd0, wReg};
  assign _zz__zz_realValue_0_89_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_89_1 = (_zz_realValue_0_89_2 + _zz_realValue_0_89_3);
  assign _zz_realValue_0_89_2 = {1'd0, wReg};
  assign _zz_realValue_0_89_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_89_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_89 = {1'd0, _zz_when_ArraySlice_l166_89_1};
  assign _zz_when_ArraySlice_l166_89_2 = (_zz_when_ArraySlice_l166_89_3 + _zz_when_ArraySlice_l166_89_7);
  assign _zz_when_ArraySlice_l166_89_3 = (realValue_0_89 - _zz_when_ArraySlice_l166_89_4);
  assign _zz_when_ArraySlice_l166_89_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_89_5);
  assign _zz_when_ArraySlice_l166_89_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_89_5 = {3'd0, _zz_when_ArraySlice_l166_89_6};
  assign _zz_when_ArraySlice_l166_89_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_90 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_90_1);
  assign _zz_when_ArraySlice_l158_90_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_90_1 = {2'd0, _zz_when_ArraySlice_l158_90_2};
  assign _zz_when_ArraySlice_l158_90_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_90_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_90 = {1'd0, _zz_when_ArraySlice_l159_90_1};
  assign _zz_when_ArraySlice_l159_90_2 = (_zz_when_ArraySlice_l159_90_3 - _zz_when_ArraySlice_l159_90_4);
  assign _zz_when_ArraySlice_l159_90_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_90_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_90_5);
  assign _zz_when_ArraySlice_l159_90_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_90_5 = {2'd0, _zz_when_ArraySlice_l159_90_6};
  assign _zz__zz_realValue_0_90 = {1'd0, wReg};
  assign _zz__zz_realValue_0_90_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_90_1 = (_zz_realValue_0_90_2 + _zz_realValue_0_90_3);
  assign _zz_realValue_0_90_2 = {1'd0, wReg};
  assign _zz_realValue_0_90_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_90_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_90 = {1'd0, _zz_when_ArraySlice_l166_90_1};
  assign _zz_when_ArraySlice_l166_90_2 = (_zz_when_ArraySlice_l166_90_3 + _zz_when_ArraySlice_l166_90_7);
  assign _zz_when_ArraySlice_l166_90_3 = (realValue_0_90 - _zz_when_ArraySlice_l166_90_4);
  assign _zz_when_ArraySlice_l166_90_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_90_5);
  assign _zz_when_ArraySlice_l166_90_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_90_5 = {2'd0, _zz_when_ArraySlice_l166_90_6};
  assign _zz_when_ArraySlice_l166_90_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_91 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_91_1);
  assign _zz_when_ArraySlice_l158_91_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_91_1 = {2'd0, _zz_when_ArraySlice_l158_91_2};
  assign _zz_when_ArraySlice_l158_91_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_91_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_91 = {1'd0, _zz_when_ArraySlice_l159_91_1};
  assign _zz_when_ArraySlice_l159_91_2 = (_zz_when_ArraySlice_l159_91_3 - _zz_when_ArraySlice_l159_91_4);
  assign _zz_when_ArraySlice_l159_91_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_91_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_91_5);
  assign _zz_when_ArraySlice_l159_91_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_91_5 = {2'd0, _zz_when_ArraySlice_l159_91_6};
  assign _zz__zz_realValue_0_91 = {1'd0, wReg};
  assign _zz__zz_realValue_0_91_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_91_1 = (_zz_realValue_0_91_2 + _zz_realValue_0_91_3);
  assign _zz_realValue_0_91_2 = {1'd0, wReg};
  assign _zz_realValue_0_91_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_91_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_91 = {1'd0, _zz_when_ArraySlice_l166_91_1};
  assign _zz_when_ArraySlice_l166_91_2 = (_zz_when_ArraySlice_l166_91_3 + _zz_when_ArraySlice_l166_91_7);
  assign _zz_when_ArraySlice_l166_91_3 = (realValue_0_91 - _zz_when_ArraySlice_l166_91_4);
  assign _zz_when_ArraySlice_l166_91_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_91_5);
  assign _zz_when_ArraySlice_l166_91_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_91_5 = {2'd0, _zz_when_ArraySlice_l166_91_6};
  assign _zz_when_ArraySlice_l166_91_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_92 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_92_1);
  assign _zz_when_ArraySlice_l158_92_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_92_1 = {1'd0, _zz_when_ArraySlice_l158_92_2};
  assign _zz_when_ArraySlice_l158_92_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_92_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_92 = {1'd0, _zz_when_ArraySlice_l159_92_1};
  assign _zz_when_ArraySlice_l159_92_2 = (_zz_when_ArraySlice_l159_92_3 - _zz_when_ArraySlice_l159_92_4);
  assign _zz_when_ArraySlice_l159_92_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_92_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_92_5);
  assign _zz_when_ArraySlice_l159_92_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_92_5 = {1'd0, _zz_when_ArraySlice_l159_92_6};
  assign _zz__zz_realValue_0_92 = {1'd0, wReg};
  assign _zz__zz_realValue_0_92_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_92_1 = (_zz_realValue_0_92_2 + _zz_realValue_0_92_3);
  assign _zz_realValue_0_92_2 = {1'd0, wReg};
  assign _zz_realValue_0_92_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_92_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_92 = {1'd0, _zz_when_ArraySlice_l166_92_1};
  assign _zz_when_ArraySlice_l166_92_2 = (_zz_when_ArraySlice_l166_92_3 + _zz_when_ArraySlice_l166_92_7);
  assign _zz_when_ArraySlice_l166_92_3 = (realValue_0_92 - _zz_when_ArraySlice_l166_92_4);
  assign _zz_when_ArraySlice_l166_92_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_92_5);
  assign _zz_when_ArraySlice_l166_92_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_92_5 = {1'd0, _zz_when_ArraySlice_l166_92_6};
  assign _zz_when_ArraySlice_l166_92_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_93 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_93_1);
  assign _zz_when_ArraySlice_l158_93_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_93_1 = {1'd0, _zz_when_ArraySlice_l158_93_2};
  assign _zz_when_ArraySlice_l158_93_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_93_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_93 = {2'd0, _zz_when_ArraySlice_l159_93_1};
  assign _zz_when_ArraySlice_l159_93_2 = (_zz_when_ArraySlice_l159_93_3 - _zz_when_ArraySlice_l159_93_4);
  assign _zz_when_ArraySlice_l159_93_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_93_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_93_5);
  assign _zz_when_ArraySlice_l159_93_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_93_5 = {1'd0, _zz_when_ArraySlice_l159_93_6};
  assign _zz__zz_realValue_0_93 = {1'd0, wReg};
  assign _zz__zz_realValue_0_93_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_93_1 = (_zz_realValue_0_93_2 + _zz_realValue_0_93_3);
  assign _zz_realValue_0_93_2 = {1'd0, wReg};
  assign _zz_realValue_0_93_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_93_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_93 = {2'd0, _zz_when_ArraySlice_l166_93_1};
  assign _zz_when_ArraySlice_l166_93_2 = (_zz_when_ArraySlice_l166_93_3 + _zz_when_ArraySlice_l166_93_7);
  assign _zz_when_ArraySlice_l166_93_3 = (realValue_0_93 - _zz_when_ArraySlice_l166_93_4);
  assign _zz_when_ArraySlice_l166_93_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_93_5);
  assign _zz_when_ArraySlice_l166_93_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_93_5 = {1'd0, _zz_when_ArraySlice_l166_93_6};
  assign _zz_when_ArraySlice_l166_93_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_94 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_94_1);
  assign _zz_when_ArraySlice_l158_94_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_94_1 = {1'd0, _zz_when_ArraySlice_l158_94_2};
  assign _zz_when_ArraySlice_l158_94_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_94_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_94 = {2'd0, _zz_when_ArraySlice_l159_94_1};
  assign _zz_when_ArraySlice_l159_94_2 = (_zz_when_ArraySlice_l159_94_3 - _zz_when_ArraySlice_l159_94_4);
  assign _zz_when_ArraySlice_l159_94_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_94_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_94_5);
  assign _zz_when_ArraySlice_l159_94_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_94_5 = {1'd0, _zz_when_ArraySlice_l159_94_6};
  assign _zz__zz_realValue_0_94 = {1'd0, wReg};
  assign _zz__zz_realValue_0_94_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_94_1 = (_zz_realValue_0_94_2 + _zz_realValue_0_94_3);
  assign _zz_realValue_0_94_2 = {1'd0, wReg};
  assign _zz_realValue_0_94_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_94_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_94 = {2'd0, _zz_when_ArraySlice_l166_94_1};
  assign _zz_when_ArraySlice_l166_94_2 = (_zz_when_ArraySlice_l166_94_3 + _zz_when_ArraySlice_l166_94_7);
  assign _zz_when_ArraySlice_l166_94_3 = (realValue_0_94 - _zz_when_ArraySlice_l166_94_4);
  assign _zz_when_ArraySlice_l166_94_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_94_5);
  assign _zz_when_ArraySlice_l166_94_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_94_5 = {1'd0, _zz_when_ArraySlice_l166_94_6};
  assign _zz_when_ArraySlice_l166_94_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_95 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_95_1);
  assign _zz_when_ArraySlice_l158_95_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_95_1 = {1'd0, _zz_when_ArraySlice_l158_95_2};
  assign _zz_when_ArraySlice_l158_95_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_95_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_95 = {3'd0, _zz_when_ArraySlice_l159_95_1};
  assign _zz_when_ArraySlice_l159_95_2 = (_zz_when_ArraySlice_l159_95_3 - _zz_when_ArraySlice_l159_95_4);
  assign _zz_when_ArraySlice_l159_95_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_95_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_95_5);
  assign _zz_when_ArraySlice_l159_95_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_95_5 = {1'd0, _zz_when_ArraySlice_l159_95_6};
  assign _zz__zz_realValue_0_95 = {1'd0, wReg};
  assign _zz__zz_realValue_0_95_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_95_1 = (_zz_realValue_0_95_2 + _zz_realValue_0_95_3);
  assign _zz_realValue_0_95_2 = {1'd0, wReg};
  assign _zz_realValue_0_95_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_95_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_95 = {3'd0, _zz_when_ArraySlice_l166_95_1};
  assign _zz_when_ArraySlice_l166_95_2 = (_zz_when_ArraySlice_l166_95_3 + _zz_when_ArraySlice_l166_95_7);
  assign _zz_when_ArraySlice_l166_95_3 = (realValue_0_95 - _zz_when_ArraySlice_l166_95_4);
  assign _zz_when_ArraySlice_l166_95_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_95_5);
  assign _zz_when_ArraySlice_l166_95_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_95_5 = {1'd0, _zz_when_ArraySlice_l166_95_6};
  assign _zz_when_ArraySlice_l166_95_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_3_2 = (_zz_when_ArraySlice_l428_3_3 + _zz_when_ArraySlice_l428_3_7);
  assign _zz_when_ArraySlice_l428_3_3 = (_zz_when_ArraySlice_l428_3_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l428_3_5);
  assign _zz_when_ArraySlice_l428_3_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_3_5 = {1'd0, _zz_when_ArraySlice_l428_3_6};
  assign _zz_when_ArraySlice_l428_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l428_3_7 = {2'd0, _zz_when_ArraySlice_l428_3_8};
  assign _zz_when_ArraySlice_l431_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_3_2 = (_zz_when_ArraySlice_l431_3_3 + 8'h01);
  assign _zz_when_ArraySlice_l431_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l431_3_4);
  assign _zz_when_ArraySlice_l431_3_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_3_4 = {1'd0, _zz_when_ArraySlice_l431_3_5};
  assign _zz_selectReadFifo_3_11 = (selectReadFifo_3 + _zz_selectReadFifo_3_12);
  assign _zz_selectReadFifo_3_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_12 = {1'd0, _zz_selectReadFifo_3_13};
  assign _zz_when_ArraySlice_l438_3 = (_zz_when_ArraySlice_l438_3_1 % aReg);
  assign _zz_when_ArraySlice_l438_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_3_1 = (_zz_when_ArraySlice_l449_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l449_3 = {5'd0, _zz_when_ArraySlice_l449_3_1};
  assign _zz_when_ArraySlice_l449_3_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_11 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_11_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_11_1 = (_zz_realValue1_0_11_2 + _zz_realValue1_0_11_3);
  assign _zz_realValue1_0_11_2 = {1'd0, hReg};
  assign _zz_realValue1_0_11_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l450_3 = {1'd0, _zz_when_ArraySlice_l450_3_1};
  assign _zz_when_ArraySlice_l450_3_2 = (realValue1_0_11 / aReg);
  assign _zz_selectReadFifo_3_14 = (selectReadFifo_3 - _zz_selectReadFifo_3_15);
  assign _zz_selectReadFifo_3_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_96 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_96_1);
  assign _zz_when_ArraySlice_l158_96_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_96_1 = {4'd0, _zz_when_ArraySlice_l158_96_2};
  assign _zz_when_ArraySlice_l158_96_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_96 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_96_1 = (_zz_when_ArraySlice_l159_96_2 - _zz_when_ArraySlice_l159_96_3);
  assign _zz_when_ArraySlice_l159_96_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_96_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_96_4);
  assign _zz_when_ArraySlice_l159_96_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_96_4 = {4'd0, _zz_when_ArraySlice_l159_96_5};
  assign _zz__zz_realValue_0_96 = {1'd0, wReg};
  assign _zz__zz_realValue_0_96_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_96_1 = (_zz_realValue_0_96_2 + _zz_realValue_0_96_3);
  assign _zz_realValue_0_96_2 = {1'd0, wReg};
  assign _zz_realValue_0_96_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_96 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_96_1 = (_zz_when_ArraySlice_l166_96_2 + _zz_when_ArraySlice_l166_96_6);
  assign _zz_when_ArraySlice_l166_96_2 = (realValue_0_96 - _zz_when_ArraySlice_l166_96_3);
  assign _zz_when_ArraySlice_l166_96_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_96_4);
  assign _zz_when_ArraySlice_l166_96_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_96_4 = {4'd0, _zz_when_ArraySlice_l166_96_5};
  assign _zz_when_ArraySlice_l166_96_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_97 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_97_1);
  assign _zz_when_ArraySlice_l158_97_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_97_1 = {3'd0, _zz_when_ArraySlice_l158_97_2};
  assign _zz_when_ArraySlice_l158_97_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_97_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_97 = {1'd0, _zz_when_ArraySlice_l159_97_1};
  assign _zz_when_ArraySlice_l159_97_2 = (_zz_when_ArraySlice_l159_97_3 - _zz_when_ArraySlice_l159_97_4);
  assign _zz_when_ArraySlice_l159_97_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_97_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_97_5);
  assign _zz_when_ArraySlice_l159_97_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_97_5 = {3'd0, _zz_when_ArraySlice_l159_97_6};
  assign _zz__zz_realValue_0_97 = {1'd0, wReg};
  assign _zz__zz_realValue_0_97_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_97_1 = (_zz_realValue_0_97_2 + _zz_realValue_0_97_3);
  assign _zz_realValue_0_97_2 = {1'd0, wReg};
  assign _zz_realValue_0_97_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_97_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_97 = {1'd0, _zz_when_ArraySlice_l166_97_1};
  assign _zz_when_ArraySlice_l166_97_2 = (_zz_when_ArraySlice_l166_97_3 + _zz_when_ArraySlice_l166_97_7);
  assign _zz_when_ArraySlice_l166_97_3 = (realValue_0_97 - _zz_when_ArraySlice_l166_97_4);
  assign _zz_when_ArraySlice_l166_97_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_97_5);
  assign _zz_when_ArraySlice_l166_97_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_97_5 = {3'd0, _zz_when_ArraySlice_l166_97_6};
  assign _zz_when_ArraySlice_l166_97_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_98 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_98_1);
  assign _zz_when_ArraySlice_l158_98_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_98_1 = {2'd0, _zz_when_ArraySlice_l158_98_2};
  assign _zz_when_ArraySlice_l158_98_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_98_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_98 = {1'd0, _zz_when_ArraySlice_l159_98_1};
  assign _zz_when_ArraySlice_l159_98_2 = (_zz_when_ArraySlice_l159_98_3 - _zz_when_ArraySlice_l159_98_4);
  assign _zz_when_ArraySlice_l159_98_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_98_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_98_5);
  assign _zz_when_ArraySlice_l159_98_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_98_5 = {2'd0, _zz_when_ArraySlice_l159_98_6};
  assign _zz__zz_realValue_0_98 = {1'd0, wReg};
  assign _zz__zz_realValue_0_98_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_98_1 = (_zz_realValue_0_98_2 + _zz_realValue_0_98_3);
  assign _zz_realValue_0_98_2 = {1'd0, wReg};
  assign _zz_realValue_0_98_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_98_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_98 = {1'd0, _zz_when_ArraySlice_l166_98_1};
  assign _zz_when_ArraySlice_l166_98_2 = (_zz_when_ArraySlice_l166_98_3 + _zz_when_ArraySlice_l166_98_7);
  assign _zz_when_ArraySlice_l166_98_3 = (realValue_0_98 - _zz_when_ArraySlice_l166_98_4);
  assign _zz_when_ArraySlice_l166_98_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_98_5);
  assign _zz_when_ArraySlice_l166_98_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_98_5 = {2'd0, _zz_when_ArraySlice_l166_98_6};
  assign _zz_when_ArraySlice_l166_98_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_99 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_99_1);
  assign _zz_when_ArraySlice_l158_99_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_99_1 = {2'd0, _zz_when_ArraySlice_l158_99_2};
  assign _zz_when_ArraySlice_l158_99_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_99_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_99 = {1'd0, _zz_when_ArraySlice_l159_99_1};
  assign _zz_when_ArraySlice_l159_99_2 = (_zz_when_ArraySlice_l159_99_3 - _zz_when_ArraySlice_l159_99_4);
  assign _zz_when_ArraySlice_l159_99_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_99_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_99_5);
  assign _zz_when_ArraySlice_l159_99_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_99_5 = {2'd0, _zz_when_ArraySlice_l159_99_6};
  assign _zz__zz_realValue_0_99 = {1'd0, wReg};
  assign _zz__zz_realValue_0_99_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_99_1 = (_zz_realValue_0_99_2 + _zz_realValue_0_99_3);
  assign _zz_realValue_0_99_2 = {1'd0, wReg};
  assign _zz_realValue_0_99_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_99_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_99 = {1'd0, _zz_when_ArraySlice_l166_99_1};
  assign _zz_when_ArraySlice_l166_99_2 = (_zz_when_ArraySlice_l166_99_3 + _zz_when_ArraySlice_l166_99_7);
  assign _zz_when_ArraySlice_l166_99_3 = (realValue_0_99 - _zz_when_ArraySlice_l166_99_4);
  assign _zz_when_ArraySlice_l166_99_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_99_5);
  assign _zz_when_ArraySlice_l166_99_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_99_5 = {2'd0, _zz_when_ArraySlice_l166_99_6};
  assign _zz_when_ArraySlice_l166_99_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_100 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_100_1);
  assign _zz_when_ArraySlice_l158_100_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_100_1 = {1'd0, _zz_when_ArraySlice_l158_100_2};
  assign _zz_when_ArraySlice_l158_100_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_100_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_100 = {1'd0, _zz_when_ArraySlice_l159_100_1};
  assign _zz_when_ArraySlice_l159_100_2 = (_zz_when_ArraySlice_l159_100_3 - _zz_when_ArraySlice_l159_100_4);
  assign _zz_when_ArraySlice_l159_100_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_100_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_100_5);
  assign _zz_when_ArraySlice_l159_100_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_100_5 = {1'd0, _zz_when_ArraySlice_l159_100_6};
  assign _zz__zz_realValue_0_100 = {1'd0, wReg};
  assign _zz__zz_realValue_0_100_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_100_1 = (_zz_realValue_0_100_2 + _zz_realValue_0_100_3);
  assign _zz_realValue_0_100_2 = {1'd0, wReg};
  assign _zz_realValue_0_100_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_100_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_100 = {1'd0, _zz_when_ArraySlice_l166_100_1};
  assign _zz_when_ArraySlice_l166_100_2 = (_zz_when_ArraySlice_l166_100_3 + _zz_when_ArraySlice_l166_100_7);
  assign _zz_when_ArraySlice_l166_100_3 = (realValue_0_100 - _zz_when_ArraySlice_l166_100_4);
  assign _zz_when_ArraySlice_l166_100_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_100_5);
  assign _zz_when_ArraySlice_l166_100_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_100_5 = {1'd0, _zz_when_ArraySlice_l166_100_6};
  assign _zz_when_ArraySlice_l166_100_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_101 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_101_1);
  assign _zz_when_ArraySlice_l158_101_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_101_1 = {1'd0, _zz_when_ArraySlice_l158_101_2};
  assign _zz_when_ArraySlice_l158_101_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_101_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_101 = {2'd0, _zz_when_ArraySlice_l159_101_1};
  assign _zz_when_ArraySlice_l159_101_2 = (_zz_when_ArraySlice_l159_101_3 - _zz_when_ArraySlice_l159_101_4);
  assign _zz_when_ArraySlice_l159_101_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_101_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_101_5);
  assign _zz_when_ArraySlice_l159_101_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_101_5 = {1'd0, _zz_when_ArraySlice_l159_101_6};
  assign _zz__zz_realValue_0_101 = {1'd0, wReg};
  assign _zz__zz_realValue_0_101_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_101_1 = (_zz_realValue_0_101_2 + _zz_realValue_0_101_3);
  assign _zz_realValue_0_101_2 = {1'd0, wReg};
  assign _zz_realValue_0_101_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_101_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_101 = {2'd0, _zz_when_ArraySlice_l166_101_1};
  assign _zz_when_ArraySlice_l166_101_2 = (_zz_when_ArraySlice_l166_101_3 + _zz_when_ArraySlice_l166_101_7);
  assign _zz_when_ArraySlice_l166_101_3 = (realValue_0_101 - _zz_when_ArraySlice_l166_101_4);
  assign _zz_when_ArraySlice_l166_101_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_101_5);
  assign _zz_when_ArraySlice_l166_101_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_101_5 = {1'd0, _zz_when_ArraySlice_l166_101_6};
  assign _zz_when_ArraySlice_l166_101_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_102 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_102_1);
  assign _zz_when_ArraySlice_l158_102_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_102_1 = {1'd0, _zz_when_ArraySlice_l158_102_2};
  assign _zz_when_ArraySlice_l158_102_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_102_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_102 = {2'd0, _zz_when_ArraySlice_l159_102_1};
  assign _zz_when_ArraySlice_l159_102_2 = (_zz_when_ArraySlice_l159_102_3 - _zz_when_ArraySlice_l159_102_4);
  assign _zz_when_ArraySlice_l159_102_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_102_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_102_5);
  assign _zz_when_ArraySlice_l159_102_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_102_5 = {1'd0, _zz_when_ArraySlice_l159_102_6};
  assign _zz__zz_realValue_0_102 = {1'd0, wReg};
  assign _zz__zz_realValue_0_102_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_102_1 = (_zz_realValue_0_102_2 + _zz_realValue_0_102_3);
  assign _zz_realValue_0_102_2 = {1'd0, wReg};
  assign _zz_realValue_0_102_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_102_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_102 = {2'd0, _zz_when_ArraySlice_l166_102_1};
  assign _zz_when_ArraySlice_l166_102_2 = (_zz_when_ArraySlice_l166_102_3 + _zz_when_ArraySlice_l166_102_7);
  assign _zz_when_ArraySlice_l166_102_3 = (realValue_0_102 - _zz_when_ArraySlice_l166_102_4);
  assign _zz_when_ArraySlice_l166_102_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_102_5);
  assign _zz_when_ArraySlice_l166_102_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_102_5 = {1'd0, _zz_when_ArraySlice_l166_102_6};
  assign _zz_when_ArraySlice_l166_102_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_103 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_103_1);
  assign _zz_when_ArraySlice_l158_103_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_103_1 = {1'd0, _zz_when_ArraySlice_l158_103_2};
  assign _zz_when_ArraySlice_l158_103_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_103_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_103 = {3'd0, _zz_when_ArraySlice_l159_103_1};
  assign _zz_when_ArraySlice_l159_103_2 = (_zz_when_ArraySlice_l159_103_3 - _zz_when_ArraySlice_l159_103_4);
  assign _zz_when_ArraySlice_l159_103_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_103_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_103_5);
  assign _zz_when_ArraySlice_l159_103_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_103_5 = {1'd0, _zz_when_ArraySlice_l159_103_6};
  assign _zz__zz_realValue_0_103 = {1'd0, wReg};
  assign _zz__zz_realValue_0_103_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_103_1 = (_zz_realValue_0_103_2 + _zz_realValue_0_103_3);
  assign _zz_realValue_0_103_2 = {1'd0, wReg};
  assign _zz_realValue_0_103_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_103_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_103 = {3'd0, _zz_when_ArraySlice_l166_103_1};
  assign _zz_when_ArraySlice_l166_103_2 = (_zz_when_ArraySlice_l166_103_3 + _zz_when_ArraySlice_l166_103_7);
  assign _zz_when_ArraySlice_l166_103_3 = (realValue_0_103 - _zz_when_ArraySlice_l166_103_4);
  assign _zz_when_ArraySlice_l166_103_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_103_5);
  assign _zz_when_ArraySlice_l166_103_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_103_5 = {1'd0, _zz_when_ArraySlice_l166_103_6};
  assign _zz_when_ArraySlice_l166_103_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_3 = (_zz_when_ArraySlice_l461_3_1 % aReg);
  assign _zz_when_ArraySlice_l461_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l447_3_3);
  assign _zz_when_ArraySlice_l447_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l447_3_3 = {2'd0, _zz_when_ArraySlice_l447_3_4};
  assign _zz_when_ArraySlice_l468_3_1 = (_zz_when_ArraySlice_l468_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l468_3 = {5'd0, _zz_when_ArraySlice_l468_3_1};
  assign _zz_when_ArraySlice_l468_3_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l376_4_1);
  assign _zz_when_ArraySlice_l376_4_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l376_4_1 = {1'd0, _zz_when_ArraySlice_l376_4_2};
  assign _zz_when_ArraySlice_l376_4_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l377_4_4);
  assign _zz_when_ArraySlice_l377_4_2 = _zz_when_ArraySlice_l377_4_3[6:0];
  assign _zz_when_ArraySlice_l377_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l377_4_4 = {1'd0, _zz_when_ArraySlice_l377_4_5};
  assign _zz__zz_outputStreamArrayData_4_valid_1 = (bReg * 3'b100);
  assign _zz__zz_outputStreamArrayData_4_valid = {1'd0, _zz__zz_outputStreamArrayData_4_valid_1};
  assign _zz__zz_7 = _zz_outputStreamArrayData_4_valid[6:0];
  assign _zz_outputStreamArrayData_4_valid_3 = _zz_outputStreamArrayData_4_valid[6:0];
  assign _zz_outputStreamArrayData_4_payload_1 = _zz_outputStreamArrayData_4_valid[6:0];
  assign _zz_when_ArraySlice_l383_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l383_4_4);
  assign _zz_when_ArraySlice_l383_4_2 = _zz_when_ArraySlice_l383_4_3[6:0];
  assign _zz_when_ArraySlice_l383_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l383_4_4 = {1'd0, _zz_when_ArraySlice_l383_4_5};
  assign _zz_when_ArraySlice_l384_4_1 = (_zz_when_ArraySlice_l384_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l384_4 = {5'd0, _zz_when_ArraySlice_l384_4_1};
  assign _zz_when_ArraySlice_l384_4_2 = (bReg * aReg);
  assign _zz_selectReadFifo_4 = (selectReadFifo_4 - _zz_selectReadFifo_4_1);
  assign _zz_selectReadFifo_4_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_4 = (_zz_when_ArraySlice_l387_4_1 % aReg);
  assign _zz_when_ArraySlice_l387_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l392_4_4);
  assign _zz_when_ArraySlice_l392_4_2 = _zz_when_ArraySlice_l392_4_3[6:0];
  assign _zz_when_ArraySlice_l392_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l392_4_4 = {1'd0, _zz_when_ArraySlice_l392_4_5};
  assign _zz_when_ArraySlice_l393_4_1 = (_zz_when_ArraySlice_l393_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l393_4 = {5'd0, _zz_when_ArraySlice_l393_4_1};
  assign _zz_when_ArraySlice_l393_4_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_12 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_12_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_12_1 = (_zz_realValue1_0_12_2 + _zz_realValue1_0_12_3);
  assign _zz_realValue1_0_12_2 = {1'd0, hReg};
  assign _zz_realValue1_0_12_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l395_4 = {1'd0, _zz_when_ArraySlice_l395_4_1};
  assign _zz_when_ArraySlice_l395_4_2 = (realValue1_0_12 / aReg);
  assign _zz_selectReadFifo_4_2 = (selectReadFifo_4 - _zz_selectReadFifo_4_3);
  assign _zz_selectReadFifo_4_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_4_5 = 1'b1;
  assign _zz_selectReadFifo_4_4 = {7'd0, _zz_selectReadFifo_4_5};
  assign _zz_when_ArraySlice_l158_104 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_104_1);
  assign _zz_when_ArraySlice_l158_104_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_104_1 = {4'd0, _zz_when_ArraySlice_l158_104_2};
  assign _zz_when_ArraySlice_l158_104_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_104 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_104_1 = (_zz_when_ArraySlice_l159_104_2 - _zz_when_ArraySlice_l159_104_3);
  assign _zz_when_ArraySlice_l159_104_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_104_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_104_4);
  assign _zz_when_ArraySlice_l159_104_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_104_4 = {4'd0, _zz_when_ArraySlice_l159_104_5};
  assign _zz__zz_realValue_0_104 = {1'd0, wReg};
  assign _zz__zz_realValue_0_104_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_104_1 = (_zz_realValue_0_104_2 + _zz_realValue_0_104_3);
  assign _zz_realValue_0_104_2 = {1'd0, wReg};
  assign _zz_realValue_0_104_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_104 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_104_1 = (_zz_when_ArraySlice_l166_104_2 + _zz_when_ArraySlice_l166_104_6);
  assign _zz_when_ArraySlice_l166_104_2 = (realValue_0_104 - _zz_when_ArraySlice_l166_104_3);
  assign _zz_when_ArraySlice_l166_104_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_104_4);
  assign _zz_when_ArraySlice_l166_104_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_104_4 = {4'd0, _zz_when_ArraySlice_l166_104_5};
  assign _zz_when_ArraySlice_l166_104_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_105 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_105_1);
  assign _zz_when_ArraySlice_l158_105_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_105_1 = {3'd0, _zz_when_ArraySlice_l158_105_2};
  assign _zz_when_ArraySlice_l158_105_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_105_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_105 = {1'd0, _zz_when_ArraySlice_l159_105_1};
  assign _zz_when_ArraySlice_l159_105_2 = (_zz_when_ArraySlice_l159_105_3 - _zz_when_ArraySlice_l159_105_4);
  assign _zz_when_ArraySlice_l159_105_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_105_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_105_5);
  assign _zz_when_ArraySlice_l159_105_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_105_5 = {3'd0, _zz_when_ArraySlice_l159_105_6};
  assign _zz__zz_realValue_0_105 = {1'd0, wReg};
  assign _zz__zz_realValue_0_105_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_105_1 = (_zz_realValue_0_105_2 + _zz_realValue_0_105_3);
  assign _zz_realValue_0_105_2 = {1'd0, wReg};
  assign _zz_realValue_0_105_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_105_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_105 = {1'd0, _zz_when_ArraySlice_l166_105_1};
  assign _zz_when_ArraySlice_l166_105_2 = (_zz_when_ArraySlice_l166_105_3 + _zz_when_ArraySlice_l166_105_7);
  assign _zz_when_ArraySlice_l166_105_3 = (realValue_0_105 - _zz_when_ArraySlice_l166_105_4);
  assign _zz_when_ArraySlice_l166_105_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_105_5);
  assign _zz_when_ArraySlice_l166_105_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_105_5 = {3'd0, _zz_when_ArraySlice_l166_105_6};
  assign _zz_when_ArraySlice_l166_105_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_106 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_106_1);
  assign _zz_when_ArraySlice_l158_106_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_106_1 = {2'd0, _zz_when_ArraySlice_l158_106_2};
  assign _zz_when_ArraySlice_l158_106_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_106_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_106 = {1'd0, _zz_when_ArraySlice_l159_106_1};
  assign _zz_when_ArraySlice_l159_106_2 = (_zz_when_ArraySlice_l159_106_3 - _zz_when_ArraySlice_l159_106_4);
  assign _zz_when_ArraySlice_l159_106_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_106_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_106_5);
  assign _zz_when_ArraySlice_l159_106_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_106_5 = {2'd0, _zz_when_ArraySlice_l159_106_6};
  assign _zz__zz_realValue_0_106 = {1'd0, wReg};
  assign _zz__zz_realValue_0_106_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_106_1 = (_zz_realValue_0_106_2 + _zz_realValue_0_106_3);
  assign _zz_realValue_0_106_2 = {1'd0, wReg};
  assign _zz_realValue_0_106_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_106_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_106 = {1'd0, _zz_when_ArraySlice_l166_106_1};
  assign _zz_when_ArraySlice_l166_106_2 = (_zz_when_ArraySlice_l166_106_3 + _zz_when_ArraySlice_l166_106_7);
  assign _zz_when_ArraySlice_l166_106_3 = (realValue_0_106 - _zz_when_ArraySlice_l166_106_4);
  assign _zz_when_ArraySlice_l166_106_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_106_5);
  assign _zz_when_ArraySlice_l166_106_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_106_5 = {2'd0, _zz_when_ArraySlice_l166_106_6};
  assign _zz_when_ArraySlice_l166_106_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_107 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_107_1);
  assign _zz_when_ArraySlice_l158_107_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_107_1 = {2'd0, _zz_when_ArraySlice_l158_107_2};
  assign _zz_when_ArraySlice_l158_107_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_107_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_107 = {1'd0, _zz_when_ArraySlice_l159_107_1};
  assign _zz_when_ArraySlice_l159_107_2 = (_zz_when_ArraySlice_l159_107_3 - _zz_when_ArraySlice_l159_107_4);
  assign _zz_when_ArraySlice_l159_107_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_107_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_107_5);
  assign _zz_when_ArraySlice_l159_107_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_107_5 = {2'd0, _zz_when_ArraySlice_l159_107_6};
  assign _zz__zz_realValue_0_107 = {1'd0, wReg};
  assign _zz__zz_realValue_0_107_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_107_1 = (_zz_realValue_0_107_2 + _zz_realValue_0_107_3);
  assign _zz_realValue_0_107_2 = {1'd0, wReg};
  assign _zz_realValue_0_107_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_107_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_107 = {1'd0, _zz_when_ArraySlice_l166_107_1};
  assign _zz_when_ArraySlice_l166_107_2 = (_zz_when_ArraySlice_l166_107_3 + _zz_when_ArraySlice_l166_107_7);
  assign _zz_when_ArraySlice_l166_107_3 = (realValue_0_107 - _zz_when_ArraySlice_l166_107_4);
  assign _zz_when_ArraySlice_l166_107_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_107_5);
  assign _zz_when_ArraySlice_l166_107_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_107_5 = {2'd0, _zz_when_ArraySlice_l166_107_6};
  assign _zz_when_ArraySlice_l166_107_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_108 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_108_1);
  assign _zz_when_ArraySlice_l158_108_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_108_1 = {1'd0, _zz_when_ArraySlice_l158_108_2};
  assign _zz_when_ArraySlice_l158_108_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_108_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_108 = {1'd0, _zz_when_ArraySlice_l159_108_1};
  assign _zz_when_ArraySlice_l159_108_2 = (_zz_when_ArraySlice_l159_108_3 - _zz_when_ArraySlice_l159_108_4);
  assign _zz_when_ArraySlice_l159_108_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_108_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_108_5);
  assign _zz_when_ArraySlice_l159_108_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_108_5 = {1'd0, _zz_when_ArraySlice_l159_108_6};
  assign _zz__zz_realValue_0_108 = {1'd0, wReg};
  assign _zz__zz_realValue_0_108_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_108_1 = (_zz_realValue_0_108_2 + _zz_realValue_0_108_3);
  assign _zz_realValue_0_108_2 = {1'd0, wReg};
  assign _zz_realValue_0_108_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_108_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_108 = {1'd0, _zz_when_ArraySlice_l166_108_1};
  assign _zz_when_ArraySlice_l166_108_2 = (_zz_when_ArraySlice_l166_108_3 + _zz_when_ArraySlice_l166_108_7);
  assign _zz_when_ArraySlice_l166_108_3 = (realValue_0_108 - _zz_when_ArraySlice_l166_108_4);
  assign _zz_when_ArraySlice_l166_108_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_108_5);
  assign _zz_when_ArraySlice_l166_108_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_108_5 = {1'd0, _zz_when_ArraySlice_l166_108_6};
  assign _zz_when_ArraySlice_l166_108_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_109 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_109_1);
  assign _zz_when_ArraySlice_l158_109_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_109_1 = {1'd0, _zz_when_ArraySlice_l158_109_2};
  assign _zz_when_ArraySlice_l158_109_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_109_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_109 = {2'd0, _zz_when_ArraySlice_l159_109_1};
  assign _zz_when_ArraySlice_l159_109_2 = (_zz_when_ArraySlice_l159_109_3 - _zz_when_ArraySlice_l159_109_4);
  assign _zz_when_ArraySlice_l159_109_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_109_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_109_5);
  assign _zz_when_ArraySlice_l159_109_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_109_5 = {1'd0, _zz_when_ArraySlice_l159_109_6};
  assign _zz__zz_realValue_0_109 = {1'd0, wReg};
  assign _zz__zz_realValue_0_109_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_109_1 = (_zz_realValue_0_109_2 + _zz_realValue_0_109_3);
  assign _zz_realValue_0_109_2 = {1'd0, wReg};
  assign _zz_realValue_0_109_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_109_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_109 = {2'd0, _zz_when_ArraySlice_l166_109_1};
  assign _zz_when_ArraySlice_l166_109_2 = (_zz_when_ArraySlice_l166_109_3 + _zz_when_ArraySlice_l166_109_7);
  assign _zz_when_ArraySlice_l166_109_3 = (realValue_0_109 - _zz_when_ArraySlice_l166_109_4);
  assign _zz_when_ArraySlice_l166_109_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_109_5);
  assign _zz_when_ArraySlice_l166_109_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_109_5 = {1'd0, _zz_when_ArraySlice_l166_109_6};
  assign _zz_when_ArraySlice_l166_109_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_110 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_110_1);
  assign _zz_when_ArraySlice_l158_110_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_110_1 = {1'd0, _zz_when_ArraySlice_l158_110_2};
  assign _zz_when_ArraySlice_l158_110_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_110_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_110 = {2'd0, _zz_when_ArraySlice_l159_110_1};
  assign _zz_when_ArraySlice_l159_110_2 = (_zz_when_ArraySlice_l159_110_3 - _zz_when_ArraySlice_l159_110_4);
  assign _zz_when_ArraySlice_l159_110_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_110_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_110_5);
  assign _zz_when_ArraySlice_l159_110_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_110_5 = {1'd0, _zz_when_ArraySlice_l159_110_6};
  assign _zz__zz_realValue_0_110 = {1'd0, wReg};
  assign _zz__zz_realValue_0_110_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_110_1 = (_zz_realValue_0_110_2 + _zz_realValue_0_110_3);
  assign _zz_realValue_0_110_2 = {1'd0, wReg};
  assign _zz_realValue_0_110_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_110_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_110 = {2'd0, _zz_when_ArraySlice_l166_110_1};
  assign _zz_when_ArraySlice_l166_110_2 = (_zz_when_ArraySlice_l166_110_3 + _zz_when_ArraySlice_l166_110_7);
  assign _zz_when_ArraySlice_l166_110_3 = (realValue_0_110 - _zz_when_ArraySlice_l166_110_4);
  assign _zz_when_ArraySlice_l166_110_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_110_5);
  assign _zz_when_ArraySlice_l166_110_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_110_5 = {1'd0, _zz_when_ArraySlice_l166_110_6};
  assign _zz_when_ArraySlice_l166_110_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_111 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_111_1);
  assign _zz_when_ArraySlice_l158_111_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_111_1 = {1'd0, _zz_when_ArraySlice_l158_111_2};
  assign _zz_when_ArraySlice_l158_111_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_111_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_111 = {3'd0, _zz_when_ArraySlice_l159_111_1};
  assign _zz_when_ArraySlice_l159_111_2 = (_zz_when_ArraySlice_l159_111_3 - _zz_when_ArraySlice_l159_111_4);
  assign _zz_when_ArraySlice_l159_111_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_111_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_111_5);
  assign _zz_when_ArraySlice_l159_111_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_111_5 = {1'd0, _zz_when_ArraySlice_l159_111_6};
  assign _zz__zz_realValue_0_111 = {1'd0, wReg};
  assign _zz__zz_realValue_0_111_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_111_1 = (_zz_realValue_0_111_2 + _zz_realValue_0_111_3);
  assign _zz_realValue_0_111_2 = {1'd0, wReg};
  assign _zz_realValue_0_111_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_111_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_111 = {3'd0, _zz_when_ArraySlice_l166_111_1};
  assign _zz_when_ArraySlice_l166_111_2 = (_zz_when_ArraySlice_l166_111_3 + _zz_when_ArraySlice_l166_111_7);
  assign _zz_when_ArraySlice_l166_111_3 = (realValue_0_111 - _zz_when_ArraySlice_l166_111_4);
  assign _zz_when_ArraySlice_l166_111_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_111_5);
  assign _zz_when_ArraySlice_l166_111_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_111_5 = {1'd0, _zz_when_ArraySlice_l166_111_6};
  assign _zz_when_ArraySlice_l166_111_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_4_2 = (_zz_when_ArraySlice_l403_4_3 + _zz_when_ArraySlice_l403_4_7);
  assign _zz_when_ArraySlice_l403_4_3 = (_zz_when_ArraySlice_l403_4_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l403_4_5);
  assign _zz_when_ArraySlice_l403_4_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_4_5 = {1'd0, _zz_when_ArraySlice_l403_4_6};
  assign _zz_when_ArraySlice_l403_4_8 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l403_4_7 = {1'd0, _zz_when_ArraySlice_l403_4_8};
  assign _zz_when_ArraySlice_l406_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_4_2 = (_zz_when_ArraySlice_l406_4_3 + 8'h01);
  assign _zz_when_ArraySlice_l406_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l406_4_4);
  assign _zz_when_ArraySlice_l406_4_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_4_4 = {1'd0, _zz_when_ArraySlice_l406_4_5};
  assign _zz_selectReadFifo_4_6 = (selectReadFifo_4 + _zz_selectReadFifo_4_7);
  assign _zz_selectReadFifo_4_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_7 = {1'd0, _zz_selectReadFifo_4_8};
  assign _zz_when_ArraySlice_l413_4 = (_zz_when_ArraySlice_l413_4_1 % aReg);
  assign _zz_when_ArraySlice_l413_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l417_4_4);
  assign _zz_when_ArraySlice_l417_4_2 = _zz_when_ArraySlice_l417_4_3[6:0];
  assign _zz_when_ArraySlice_l417_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l417_4_4 = {1'd0, _zz_when_ArraySlice_l417_4_5};
  assign _zz_when_ArraySlice_l418_4_2 = (_zz_when_ArraySlice_l418_4_3 - _zz_when_ArraySlice_l418_4_4);
  assign _zz_when_ArraySlice_l418_4_1 = {5'd0, _zz_when_ArraySlice_l418_4_2};
  assign _zz_when_ArraySlice_l418_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l418_4_4 = {7'd0, _zz_when_ArraySlice_l418_4_5};
  assign _zz__zz_realValue1_0_13 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_13_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_13_1 = (_zz_realValue1_0_13_2 + _zz_realValue1_0_13_3);
  assign _zz_realValue1_0_13_2 = {1'd0, hReg};
  assign _zz_realValue1_0_13_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l420_4 = {1'd0, _zz_when_ArraySlice_l420_4_1};
  assign _zz_when_ArraySlice_l420_4_2 = (realValue1_0_13 / aReg);
  assign _zz_selectReadFifo_4_9 = (selectReadFifo_4 - _zz_selectReadFifo_4_10);
  assign _zz_selectReadFifo_4_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_112 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_112_1);
  assign _zz_when_ArraySlice_l158_112_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_112_1 = {4'd0, _zz_when_ArraySlice_l158_112_2};
  assign _zz_when_ArraySlice_l158_112_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_112 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_112_1 = (_zz_when_ArraySlice_l159_112_2 - _zz_when_ArraySlice_l159_112_3);
  assign _zz_when_ArraySlice_l159_112_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_112_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_112_4);
  assign _zz_when_ArraySlice_l159_112_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_112_4 = {4'd0, _zz_when_ArraySlice_l159_112_5};
  assign _zz__zz_realValue_0_112 = {1'd0, wReg};
  assign _zz__zz_realValue_0_112_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_112_1 = (_zz_realValue_0_112_2 + _zz_realValue_0_112_3);
  assign _zz_realValue_0_112_2 = {1'd0, wReg};
  assign _zz_realValue_0_112_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_112 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_112_1 = (_zz_when_ArraySlice_l166_112_2 + _zz_when_ArraySlice_l166_112_6);
  assign _zz_when_ArraySlice_l166_112_2 = (realValue_0_112 - _zz_when_ArraySlice_l166_112_3);
  assign _zz_when_ArraySlice_l166_112_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_112_4);
  assign _zz_when_ArraySlice_l166_112_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_112_4 = {4'd0, _zz_when_ArraySlice_l166_112_5};
  assign _zz_when_ArraySlice_l166_112_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_113 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_113_1);
  assign _zz_when_ArraySlice_l158_113_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_113_1 = {3'd0, _zz_when_ArraySlice_l158_113_2};
  assign _zz_when_ArraySlice_l158_113_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_113_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_113 = {1'd0, _zz_when_ArraySlice_l159_113_1};
  assign _zz_when_ArraySlice_l159_113_2 = (_zz_when_ArraySlice_l159_113_3 - _zz_when_ArraySlice_l159_113_4);
  assign _zz_when_ArraySlice_l159_113_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_113_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_113_5);
  assign _zz_when_ArraySlice_l159_113_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_113_5 = {3'd0, _zz_when_ArraySlice_l159_113_6};
  assign _zz__zz_realValue_0_113 = {1'd0, wReg};
  assign _zz__zz_realValue_0_113_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_113_1 = (_zz_realValue_0_113_2 + _zz_realValue_0_113_3);
  assign _zz_realValue_0_113_2 = {1'd0, wReg};
  assign _zz_realValue_0_113_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_113_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_113 = {1'd0, _zz_when_ArraySlice_l166_113_1};
  assign _zz_when_ArraySlice_l166_113_2 = (_zz_when_ArraySlice_l166_113_3 + _zz_when_ArraySlice_l166_113_7);
  assign _zz_when_ArraySlice_l166_113_3 = (realValue_0_113 - _zz_when_ArraySlice_l166_113_4);
  assign _zz_when_ArraySlice_l166_113_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_113_5);
  assign _zz_when_ArraySlice_l166_113_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_113_5 = {3'd0, _zz_when_ArraySlice_l166_113_6};
  assign _zz_when_ArraySlice_l166_113_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_114 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_114_1);
  assign _zz_when_ArraySlice_l158_114_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_114_1 = {2'd0, _zz_when_ArraySlice_l158_114_2};
  assign _zz_when_ArraySlice_l158_114_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_114_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_114 = {1'd0, _zz_when_ArraySlice_l159_114_1};
  assign _zz_when_ArraySlice_l159_114_2 = (_zz_when_ArraySlice_l159_114_3 - _zz_when_ArraySlice_l159_114_4);
  assign _zz_when_ArraySlice_l159_114_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_114_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_114_5);
  assign _zz_when_ArraySlice_l159_114_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_114_5 = {2'd0, _zz_when_ArraySlice_l159_114_6};
  assign _zz__zz_realValue_0_114 = {1'd0, wReg};
  assign _zz__zz_realValue_0_114_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_114_1 = (_zz_realValue_0_114_2 + _zz_realValue_0_114_3);
  assign _zz_realValue_0_114_2 = {1'd0, wReg};
  assign _zz_realValue_0_114_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_114_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_114 = {1'd0, _zz_when_ArraySlice_l166_114_1};
  assign _zz_when_ArraySlice_l166_114_2 = (_zz_when_ArraySlice_l166_114_3 + _zz_when_ArraySlice_l166_114_7);
  assign _zz_when_ArraySlice_l166_114_3 = (realValue_0_114 - _zz_when_ArraySlice_l166_114_4);
  assign _zz_when_ArraySlice_l166_114_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_114_5);
  assign _zz_when_ArraySlice_l166_114_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_114_5 = {2'd0, _zz_when_ArraySlice_l166_114_6};
  assign _zz_when_ArraySlice_l166_114_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_115 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_115_1);
  assign _zz_when_ArraySlice_l158_115_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_115_1 = {2'd0, _zz_when_ArraySlice_l158_115_2};
  assign _zz_when_ArraySlice_l158_115_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_115_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_115 = {1'd0, _zz_when_ArraySlice_l159_115_1};
  assign _zz_when_ArraySlice_l159_115_2 = (_zz_when_ArraySlice_l159_115_3 - _zz_when_ArraySlice_l159_115_4);
  assign _zz_when_ArraySlice_l159_115_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_115_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_115_5);
  assign _zz_when_ArraySlice_l159_115_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_115_5 = {2'd0, _zz_when_ArraySlice_l159_115_6};
  assign _zz__zz_realValue_0_115 = {1'd0, wReg};
  assign _zz__zz_realValue_0_115_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_115_1 = (_zz_realValue_0_115_2 + _zz_realValue_0_115_3);
  assign _zz_realValue_0_115_2 = {1'd0, wReg};
  assign _zz_realValue_0_115_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_115_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_115 = {1'd0, _zz_when_ArraySlice_l166_115_1};
  assign _zz_when_ArraySlice_l166_115_2 = (_zz_when_ArraySlice_l166_115_3 + _zz_when_ArraySlice_l166_115_7);
  assign _zz_when_ArraySlice_l166_115_3 = (realValue_0_115 - _zz_when_ArraySlice_l166_115_4);
  assign _zz_when_ArraySlice_l166_115_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_115_5);
  assign _zz_when_ArraySlice_l166_115_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_115_5 = {2'd0, _zz_when_ArraySlice_l166_115_6};
  assign _zz_when_ArraySlice_l166_115_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_116 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_116_1);
  assign _zz_when_ArraySlice_l158_116_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_116_1 = {1'd0, _zz_when_ArraySlice_l158_116_2};
  assign _zz_when_ArraySlice_l158_116_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_116_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_116 = {1'd0, _zz_when_ArraySlice_l159_116_1};
  assign _zz_when_ArraySlice_l159_116_2 = (_zz_when_ArraySlice_l159_116_3 - _zz_when_ArraySlice_l159_116_4);
  assign _zz_when_ArraySlice_l159_116_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_116_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_116_5);
  assign _zz_when_ArraySlice_l159_116_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_116_5 = {1'd0, _zz_when_ArraySlice_l159_116_6};
  assign _zz__zz_realValue_0_116 = {1'd0, wReg};
  assign _zz__zz_realValue_0_116_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_116_1 = (_zz_realValue_0_116_2 + _zz_realValue_0_116_3);
  assign _zz_realValue_0_116_2 = {1'd0, wReg};
  assign _zz_realValue_0_116_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_116_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_116 = {1'd0, _zz_when_ArraySlice_l166_116_1};
  assign _zz_when_ArraySlice_l166_116_2 = (_zz_when_ArraySlice_l166_116_3 + _zz_when_ArraySlice_l166_116_7);
  assign _zz_when_ArraySlice_l166_116_3 = (realValue_0_116 - _zz_when_ArraySlice_l166_116_4);
  assign _zz_when_ArraySlice_l166_116_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_116_5);
  assign _zz_when_ArraySlice_l166_116_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_116_5 = {1'd0, _zz_when_ArraySlice_l166_116_6};
  assign _zz_when_ArraySlice_l166_116_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_117 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_117_1);
  assign _zz_when_ArraySlice_l158_117_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_117_1 = {1'd0, _zz_when_ArraySlice_l158_117_2};
  assign _zz_when_ArraySlice_l158_117_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_117_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_117 = {2'd0, _zz_when_ArraySlice_l159_117_1};
  assign _zz_when_ArraySlice_l159_117_2 = (_zz_when_ArraySlice_l159_117_3 - _zz_when_ArraySlice_l159_117_4);
  assign _zz_when_ArraySlice_l159_117_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_117_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_117_5);
  assign _zz_when_ArraySlice_l159_117_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_117_5 = {1'd0, _zz_when_ArraySlice_l159_117_6};
  assign _zz__zz_realValue_0_117 = {1'd0, wReg};
  assign _zz__zz_realValue_0_117_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_117_1 = (_zz_realValue_0_117_2 + _zz_realValue_0_117_3);
  assign _zz_realValue_0_117_2 = {1'd0, wReg};
  assign _zz_realValue_0_117_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_117_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_117 = {2'd0, _zz_when_ArraySlice_l166_117_1};
  assign _zz_when_ArraySlice_l166_117_2 = (_zz_when_ArraySlice_l166_117_3 + _zz_when_ArraySlice_l166_117_7);
  assign _zz_when_ArraySlice_l166_117_3 = (realValue_0_117 - _zz_when_ArraySlice_l166_117_4);
  assign _zz_when_ArraySlice_l166_117_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_117_5);
  assign _zz_when_ArraySlice_l166_117_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_117_5 = {1'd0, _zz_when_ArraySlice_l166_117_6};
  assign _zz_when_ArraySlice_l166_117_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_118 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_118_1);
  assign _zz_when_ArraySlice_l158_118_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_118_1 = {1'd0, _zz_when_ArraySlice_l158_118_2};
  assign _zz_when_ArraySlice_l158_118_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_118_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_118 = {2'd0, _zz_when_ArraySlice_l159_118_1};
  assign _zz_when_ArraySlice_l159_118_2 = (_zz_when_ArraySlice_l159_118_3 - _zz_when_ArraySlice_l159_118_4);
  assign _zz_when_ArraySlice_l159_118_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_118_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_118_5);
  assign _zz_when_ArraySlice_l159_118_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_118_5 = {1'd0, _zz_when_ArraySlice_l159_118_6};
  assign _zz__zz_realValue_0_118 = {1'd0, wReg};
  assign _zz__zz_realValue_0_118_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_118_1 = (_zz_realValue_0_118_2 + _zz_realValue_0_118_3);
  assign _zz_realValue_0_118_2 = {1'd0, wReg};
  assign _zz_realValue_0_118_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_118_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_118 = {2'd0, _zz_when_ArraySlice_l166_118_1};
  assign _zz_when_ArraySlice_l166_118_2 = (_zz_when_ArraySlice_l166_118_3 + _zz_when_ArraySlice_l166_118_7);
  assign _zz_when_ArraySlice_l166_118_3 = (realValue_0_118 - _zz_when_ArraySlice_l166_118_4);
  assign _zz_when_ArraySlice_l166_118_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_118_5);
  assign _zz_when_ArraySlice_l166_118_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_118_5 = {1'd0, _zz_when_ArraySlice_l166_118_6};
  assign _zz_when_ArraySlice_l166_118_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_119 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_119_1);
  assign _zz_when_ArraySlice_l158_119_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_119_1 = {1'd0, _zz_when_ArraySlice_l158_119_2};
  assign _zz_when_ArraySlice_l158_119_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_119_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_119 = {3'd0, _zz_when_ArraySlice_l159_119_1};
  assign _zz_when_ArraySlice_l159_119_2 = (_zz_when_ArraySlice_l159_119_3 - _zz_when_ArraySlice_l159_119_4);
  assign _zz_when_ArraySlice_l159_119_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_119_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_119_5);
  assign _zz_when_ArraySlice_l159_119_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_119_5 = {1'd0, _zz_when_ArraySlice_l159_119_6};
  assign _zz__zz_realValue_0_119 = {1'd0, wReg};
  assign _zz__zz_realValue_0_119_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_119_1 = (_zz_realValue_0_119_2 + _zz_realValue_0_119_3);
  assign _zz_realValue_0_119_2 = {1'd0, wReg};
  assign _zz_realValue_0_119_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_119_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_119 = {3'd0, _zz_when_ArraySlice_l166_119_1};
  assign _zz_when_ArraySlice_l166_119_2 = (_zz_when_ArraySlice_l166_119_3 + _zz_when_ArraySlice_l166_119_7);
  assign _zz_when_ArraySlice_l166_119_3 = (realValue_0_119 - _zz_when_ArraySlice_l166_119_4);
  assign _zz_when_ArraySlice_l166_119_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_119_5);
  assign _zz_when_ArraySlice_l166_119_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_119_5 = {1'd0, _zz_when_ArraySlice_l166_119_6};
  assign _zz_when_ArraySlice_l166_119_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_4_2 = (_zz_when_ArraySlice_l428_4_3 + _zz_when_ArraySlice_l428_4_7);
  assign _zz_when_ArraySlice_l428_4_3 = (_zz_when_ArraySlice_l428_4_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l428_4_5);
  assign _zz_when_ArraySlice_l428_4_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_4_5 = {1'd0, _zz_when_ArraySlice_l428_4_6};
  assign _zz_when_ArraySlice_l428_4_8 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l428_4_7 = {1'd0, _zz_when_ArraySlice_l428_4_8};
  assign _zz_when_ArraySlice_l431_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_4_2 = (_zz_when_ArraySlice_l431_4_3 + 8'h01);
  assign _zz_when_ArraySlice_l431_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l431_4_4);
  assign _zz_when_ArraySlice_l431_4_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_4_4 = {1'd0, _zz_when_ArraySlice_l431_4_5};
  assign _zz_selectReadFifo_4_11 = (selectReadFifo_4 + _zz_selectReadFifo_4_12);
  assign _zz_selectReadFifo_4_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_12 = {1'd0, _zz_selectReadFifo_4_13};
  assign _zz_when_ArraySlice_l438_4 = (_zz_when_ArraySlice_l438_4_1 % aReg);
  assign _zz_when_ArraySlice_l438_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_4_1 = (_zz_when_ArraySlice_l449_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l449_4 = {5'd0, _zz_when_ArraySlice_l449_4_1};
  assign _zz_when_ArraySlice_l449_4_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_14 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_14_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_14_1 = (_zz_realValue1_0_14_2 + _zz_realValue1_0_14_3);
  assign _zz_realValue1_0_14_2 = {1'd0, hReg};
  assign _zz_realValue1_0_14_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l450_4 = {1'd0, _zz_when_ArraySlice_l450_4_1};
  assign _zz_when_ArraySlice_l450_4_2 = (realValue1_0_14 / aReg);
  assign _zz_selectReadFifo_4_14 = (selectReadFifo_4 - _zz_selectReadFifo_4_15);
  assign _zz_selectReadFifo_4_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_120 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_120_1);
  assign _zz_when_ArraySlice_l158_120_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_120_1 = {4'd0, _zz_when_ArraySlice_l158_120_2};
  assign _zz_when_ArraySlice_l158_120_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_120 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_120_1 = (_zz_when_ArraySlice_l159_120_2 - _zz_when_ArraySlice_l159_120_3);
  assign _zz_when_ArraySlice_l159_120_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_120_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_120_4);
  assign _zz_when_ArraySlice_l159_120_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_120_4 = {4'd0, _zz_when_ArraySlice_l159_120_5};
  assign _zz__zz_realValue_0_120 = {1'd0, wReg};
  assign _zz__zz_realValue_0_120_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_120_1 = (_zz_realValue_0_120_2 + _zz_realValue_0_120_3);
  assign _zz_realValue_0_120_2 = {1'd0, wReg};
  assign _zz_realValue_0_120_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_120 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_120_1 = (_zz_when_ArraySlice_l166_120_2 + _zz_when_ArraySlice_l166_120_6);
  assign _zz_when_ArraySlice_l166_120_2 = (realValue_0_120 - _zz_when_ArraySlice_l166_120_3);
  assign _zz_when_ArraySlice_l166_120_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_120_4);
  assign _zz_when_ArraySlice_l166_120_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_120_4 = {4'd0, _zz_when_ArraySlice_l166_120_5};
  assign _zz_when_ArraySlice_l166_120_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_121 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_121_1);
  assign _zz_when_ArraySlice_l158_121_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_121_1 = {3'd0, _zz_when_ArraySlice_l158_121_2};
  assign _zz_when_ArraySlice_l158_121_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_121_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_121 = {1'd0, _zz_when_ArraySlice_l159_121_1};
  assign _zz_when_ArraySlice_l159_121_2 = (_zz_when_ArraySlice_l159_121_3 - _zz_when_ArraySlice_l159_121_4);
  assign _zz_when_ArraySlice_l159_121_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_121_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_121_5);
  assign _zz_when_ArraySlice_l159_121_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_121_5 = {3'd0, _zz_when_ArraySlice_l159_121_6};
  assign _zz__zz_realValue_0_121 = {1'd0, wReg};
  assign _zz__zz_realValue_0_121_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_121_1 = (_zz_realValue_0_121_2 + _zz_realValue_0_121_3);
  assign _zz_realValue_0_121_2 = {1'd0, wReg};
  assign _zz_realValue_0_121_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_121_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_121 = {1'd0, _zz_when_ArraySlice_l166_121_1};
  assign _zz_when_ArraySlice_l166_121_2 = (_zz_when_ArraySlice_l166_121_3 + _zz_when_ArraySlice_l166_121_7);
  assign _zz_when_ArraySlice_l166_121_3 = (realValue_0_121 - _zz_when_ArraySlice_l166_121_4);
  assign _zz_when_ArraySlice_l166_121_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_121_5);
  assign _zz_when_ArraySlice_l166_121_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_121_5 = {3'd0, _zz_when_ArraySlice_l166_121_6};
  assign _zz_when_ArraySlice_l166_121_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_122 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_122_1);
  assign _zz_when_ArraySlice_l158_122_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_122_1 = {2'd0, _zz_when_ArraySlice_l158_122_2};
  assign _zz_when_ArraySlice_l158_122_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_122_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_122 = {1'd0, _zz_when_ArraySlice_l159_122_1};
  assign _zz_when_ArraySlice_l159_122_2 = (_zz_when_ArraySlice_l159_122_3 - _zz_when_ArraySlice_l159_122_4);
  assign _zz_when_ArraySlice_l159_122_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_122_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_122_5);
  assign _zz_when_ArraySlice_l159_122_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_122_5 = {2'd0, _zz_when_ArraySlice_l159_122_6};
  assign _zz__zz_realValue_0_122 = {1'd0, wReg};
  assign _zz__zz_realValue_0_122_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_122_1 = (_zz_realValue_0_122_2 + _zz_realValue_0_122_3);
  assign _zz_realValue_0_122_2 = {1'd0, wReg};
  assign _zz_realValue_0_122_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_122_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_122 = {1'd0, _zz_when_ArraySlice_l166_122_1};
  assign _zz_when_ArraySlice_l166_122_2 = (_zz_when_ArraySlice_l166_122_3 + _zz_when_ArraySlice_l166_122_7);
  assign _zz_when_ArraySlice_l166_122_3 = (realValue_0_122 - _zz_when_ArraySlice_l166_122_4);
  assign _zz_when_ArraySlice_l166_122_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_122_5);
  assign _zz_when_ArraySlice_l166_122_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_122_5 = {2'd0, _zz_when_ArraySlice_l166_122_6};
  assign _zz_when_ArraySlice_l166_122_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_123 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_123_1);
  assign _zz_when_ArraySlice_l158_123_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_123_1 = {2'd0, _zz_when_ArraySlice_l158_123_2};
  assign _zz_when_ArraySlice_l158_123_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_123_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_123 = {1'd0, _zz_when_ArraySlice_l159_123_1};
  assign _zz_when_ArraySlice_l159_123_2 = (_zz_when_ArraySlice_l159_123_3 - _zz_when_ArraySlice_l159_123_4);
  assign _zz_when_ArraySlice_l159_123_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_123_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_123_5);
  assign _zz_when_ArraySlice_l159_123_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_123_5 = {2'd0, _zz_when_ArraySlice_l159_123_6};
  assign _zz__zz_realValue_0_123 = {1'd0, wReg};
  assign _zz__zz_realValue_0_123_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_123_1 = (_zz_realValue_0_123_2 + _zz_realValue_0_123_3);
  assign _zz_realValue_0_123_2 = {1'd0, wReg};
  assign _zz_realValue_0_123_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_123_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_123 = {1'd0, _zz_when_ArraySlice_l166_123_1};
  assign _zz_when_ArraySlice_l166_123_2 = (_zz_when_ArraySlice_l166_123_3 + _zz_when_ArraySlice_l166_123_7);
  assign _zz_when_ArraySlice_l166_123_3 = (realValue_0_123 - _zz_when_ArraySlice_l166_123_4);
  assign _zz_when_ArraySlice_l166_123_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_123_5);
  assign _zz_when_ArraySlice_l166_123_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_123_5 = {2'd0, _zz_when_ArraySlice_l166_123_6};
  assign _zz_when_ArraySlice_l166_123_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_124 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_124_1);
  assign _zz_when_ArraySlice_l158_124_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_124_1 = {1'd0, _zz_when_ArraySlice_l158_124_2};
  assign _zz_when_ArraySlice_l158_124_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_124_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_124 = {1'd0, _zz_when_ArraySlice_l159_124_1};
  assign _zz_when_ArraySlice_l159_124_2 = (_zz_when_ArraySlice_l159_124_3 - _zz_when_ArraySlice_l159_124_4);
  assign _zz_when_ArraySlice_l159_124_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_124_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_124_5);
  assign _zz_when_ArraySlice_l159_124_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_124_5 = {1'd0, _zz_when_ArraySlice_l159_124_6};
  assign _zz__zz_realValue_0_124 = {1'd0, wReg};
  assign _zz__zz_realValue_0_124_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_124_1 = (_zz_realValue_0_124_2 + _zz_realValue_0_124_3);
  assign _zz_realValue_0_124_2 = {1'd0, wReg};
  assign _zz_realValue_0_124_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_124_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_124 = {1'd0, _zz_when_ArraySlice_l166_124_1};
  assign _zz_when_ArraySlice_l166_124_2 = (_zz_when_ArraySlice_l166_124_3 + _zz_when_ArraySlice_l166_124_7);
  assign _zz_when_ArraySlice_l166_124_3 = (realValue_0_124 - _zz_when_ArraySlice_l166_124_4);
  assign _zz_when_ArraySlice_l166_124_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_124_5);
  assign _zz_when_ArraySlice_l166_124_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_124_5 = {1'd0, _zz_when_ArraySlice_l166_124_6};
  assign _zz_when_ArraySlice_l166_124_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_125 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_125_1);
  assign _zz_when_ArraySlice_l158_125_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_125_1 = {1'd0, _zz_when_ArraySlice_l158_125_2};
  assign _zz_when_ArraySlice_l158_125_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_125_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_125 = {2'd0, _zz_when_ArraySlice_l159_125_1};
  assign _zz_when_ArraySlice_l159_125_2 = (_zz_when_ArraySlice_l159_125_3 - _zz_when_ArraySlice_l159_125_4);
  assign _zz_when_ArraySlice_l159_125_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_125_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_125_5);
  assign _zz_when_ArraySlice_l159_125_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_125_5 = {1'd0, _zz_when_ArraySlice_l159_125_6};
  assign _zz__zz_realValue_0_125 = {1'd0, wReg};
  assign _zz__zz_realValue_0_125_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_125_1 = (_zz_realValue_0_125_2 + _zz_realValue_0_125_3);
  assign _zz_realValue_0_125_2 = {1'd0, wReg};
  assign _zz_realValue_0_125_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_125_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_125 = {2'd0, _zz_when_ArraySlice_l166_125_1};
  assign _zz_when_ArraySlice_l166_125_2 = (_zz_when_ArraySlice_l166_125_3 + _zz_when_ArraySlice_l166_125_7);
  assign _zz_when_ArraySlice_l166_125_3 = (realValue_0_125 - _zz_when_ArraySlice_l166_125_4);
  assign _zz_when_ArraySlice_l166_125_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_125_5);
  assign _zz_when_ArraySlice_l166_125_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_125_5 = {1'd0, _zz_when_ArraySlice_l166_125_6};
  assign _zz_when_ArraySlice_l166_125_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_126 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_126_1);
  assign _zz_when_ArraySlice_l158_126_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_126_1 = {1'd0, _zz_when_ArraySlice_l158_126_2};
  assign _zz_when_ArraySlice_l158_126_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_126_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_126 = {2'd0, _zz_when_ArraySlice_l159_126_1};
  assign _zz_when_ArraySlice_l159_126_2 = (_zz_when_ArraySlice_l159_126_3 - _zz_when_ArraySlice_l159_126_4);
  assign _zz_when_ArraySlice_l159_126_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_126_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_126_5);
  assign _zz_when_ArraySlice_l159_126_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_126_5 = {1'd0, _zz_when_ArraySlice_l159_126_6};
  assign _zz__zz_realValue_0_126 = {1'd0, wReg};
  assign _zz__zz_realValue_0_126_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_126_1 = (_zz_realValue_0_126_2 + _zz_realValue_0_126_3);
  assign _zz_realValue_0_126_2 = {1'd0, wReg};
  assign _zz_realValue_0_126_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_126_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_126 = {2'd0, _zz_when_ArraySlice_l166_126_1};
  assign _zz_when_ArraySlice_l166_126_2 = (_zz_when_ArraySlice_l166_126_3 + _zz_when_ArraySlice_l166_126_7);
  assign _zz_when_ArraySlice_l166_126_3 = (realValue_0_126 - _zz_when_ArraySlice_l166_126_4);
  assign _zz_when_ArraySlice_l166_126_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_126_5);
  assign _zz_when_ArraySlice_l166_126_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_126_5 = {1'd0, _zz_when_ArraySlice_l166_126_6};
  assign _zz_when_ArraySlice_l166_126_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_127 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_127_1);
  assign _zz_when_ArraySlice_l158_127_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_127_1 = {1'd0, _zz_when_ArraySlice_l158_127_2};
  assign _zz_when_ArraySlice_l158_127_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_127_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_127 = {3'd0, _zz_when_ArraySlice_l159_127_1};
  assign _zz_when_ArraySlice_l159_127_2 = (_zz_when_ArraySlice_l159_127_3 - _zz_when_ArraySlice_l159_127_4);
  assign _zz_when_ArraySlice_l159_127_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_127_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_127_5);
  assign _zz_when_ArraySlice_l159_127_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_127_5 = {1'd0, _zz_when_ArraySlice_l159_127_6};
  assign _zz__zz_realValue_0_127 = {1'd0, wReg};
  assign _zz__zz_realValue_0_127_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_127_1 = (_zz_realValue_0_127_2 + _zz_realValue_0_127_3);
  assign _zz_realValue_0_127_2 = {1'd0, wReg};
  assign _zz_realValue_0_127_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_127_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_127 = {3'd0, _zz_when_ArraySlice_l166_127_1};
  assign _zz_when_ArraySlice_l166_127_2 = (_zz_when_ArraySlice_l166_127_3 + _zz_when_ArraySlice_l166_127_7);
  assign _zz_when_ArraySlice_l166_127_3 = (realValue_0_127 - _zz_when_ArraySlice_l166_127_4);
  assign _zz_when_ArraySlice_l166_127_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_127_5);
  assign _zz_when_ArraySlice_l166_127_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_127_5 = {1'd0, _zz_when_ArraySlice_l166_127_6};
  assign _zz_when_ArraySlice_l166_127_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_4 = (_zz_when_ArraySlice_l461_4_1 % aReg);
  assign _zz_when_ArraySlice_l461_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l447_4_2);
  assign _zz_when_ArraySlice_l447_4_3 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l447_4_2 = {1'd0, _zz_when_ArraySlice_l447_4_3};
  assign _zz_when_ArraySlice_l468_4_1 = (_zz_when_ArraySlice_l468_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l468_4 = {5'd0, _zz_when_ArraySlice_l468_4_1};
  assign _zz_when_ArraySlice_l468_4_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l376_5_1);
  assign _zz_when_ArraySlice_l376_5_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l376_5_1 = {1'd0, _zz_when_ArraySlice_l376_5_2};
  assign _zz_when_ArraySlice_l376_5_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l377_5_3);
  assign _zz_when_ArraySlice_l377_5_1 = _zz_when_ArraySlice_l377_5_2[6:0];
  assign _zz_when_ArraySlice_l377_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l377_5_3 = {1'd0, _zz_when_ArraySlice_l377_5_4};
  assign _zz__zz_outputStreamArrayData_5_valid_1 = (bReg * 3'b101);
  assign _zz__zz_outputStreamArrayData_5_valid = {1'd0, _zz__zz_outputStreamArrayData_5_valid_1};
  assign _zz__zz_8 = _zz_outputStreamArrayData_5_valid[6:0];
  assign _zz_outputStreamArrayData_5_valid_3 = _zz_outputStreamArrayData_5_valid[6:0];
  assign _zz_outputStreamArrayData_5_payload_1 = _zz_outputStreamArrayData_5_valid[6:0];
  assign _zz_when_ArraySlice_l383_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l383_5_3);
  assign _zz_when_ArraySlice_l383_5_1 = _zz_when_ArraySlice_l383_5_2[6:0];
  assign _zz_when_ArraySlice_l383_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l383_5_3 = {1'd0, _zz_when_ArraySlice_l383_5_4};
  assign _zz_when_ArraySlice_l384_5_1 = (_zz_when_ArraySlice_l384_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l384_5 = {5'd0, _zz_when_ArraySlice_l384_5_1};
  assign _zz_when_ArraySlice_l384_5_2 = (bReg * aReg);
  assign _zz_selectReadFifo_5 = (selectReadFifo_5 - _zz_selectReadFifo_5_1);
  assign _zz_selectReadFifo_5_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_5 = (_zz_when_ArraySlice_l387_5_1 % aReg);
  assign _zz_when_ArraySlice_l387_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l392_5_3);
  assign _zz_when_ArraySlice_l392_5_1 = _zz_when_ArraySlice_l392_5_2[6:0];
  assign _zz_when_ArraySlice_l392_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l392_5_3 = {1'd0, _zz_when_ArraySlice_l392_5_4};
  assign _zz_when_ArraySlice_l393_5_1 = (_zz_when_ArraySlice_l393_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l393_5 = {5'd0, _zz_when_ArraySlice_l393_5_1};
  assign _zz_when_ArraySlice_l393_5_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_15 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_15_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_15_1 = (_zz_realValue1_0_15_2 + _zz_realValue1_0_15_3);
  assign _zz_realValue1_0_15_2 = {1'd0, hReg};
  assign _zz_realValue1_0_15_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l395_5 = {1'd0, _zz_when_ArraySlice_l395_5_1};
  assign _zz_when_ArraySlice_l395_5_2 = (realValue1_0_15 / aReg);
  assign _zz_selectReadFifo_5_2 = (selectReadFifo_5 - _zz_selectReadFifo_5_3);
  assign _zz_selectReadFifo_5_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_5_5 = 1'b1;
  assign _zz_selectReadFifo_5_4 = {7'd0, _zz_selectReadFifo_5_5};
  assign _zz_when_ArraySlice_l158_128 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_128_1);
  assign _zz_when_ArraySlice_l158_128_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_128_1 = {4'd0, _zz_when_ArraySlice_l158_128_2};
  assign _zz_when_ArraySlice_l158_128_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_128 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_128_1 = (_zz_when_ArraySlice_l159_128_2 - _zz_when_ArraySlice_l159_128_3);
  assign _zz_when_ArraySlice_l159_128_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_128_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_128_4);
  assign _zz_when_ArraySlice_l159_128_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_128_4 = {4'd0, _zz_when_ArraySlice_l159_128_5};
  assign _zz__zz_realValue_0_128 = {1'd0, wReg};
  assign _zz__zz_realValue_0_128_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_128_1 = (_zz_realValue_0_128_2 + _zz_realValue_0_128_3);
  assign _zz_realValue_0_128_2 = {1'd0, wReg};
  assign _zz_realValue_0_128_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_128 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_128_1 = (_zz_when_ArraySlice_l166_128_2 + _zz_when_ArraySlice_l166_128_6);
  assign _zz_when_ArraySlice_l166_128_2 = (realValue_0_128 - _zz_when_ArraySlice_l166_128_3);
  assign _zz_when_ArraySlice_l166_128_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_128_4);
  assign _zz_when_ArraySlice_l166_128_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_128_4 = {4'd0, _zz_when_ArraySlice_l166_128_5};
  assign _zz_when_ArraySlice_l166_128_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_129 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_129_1);
  assign _zz_when_ArraySlice_l158_129_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_129_1 = {3'd0, _zz_when_ArraySlice_l158_129_2};
  assign _zz_when_ArraySlice_l158_129_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_129_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_129 = {1'd0, _zz_when_ArraySlice_l159_129_1};
  assign _zz_when_ArraySlice_l159_129_2 = (_zz_when_ArraySlice_l159_129_3 - _zz_when_ArraySlice_l159_129_4);
  assign _zz_when_ArraySlice_l159_129_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_129_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_129_5);
  assign _zz_when_ArraySlice_l159_129_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_129_5 = {3'd0, _zz_when_ArraySlice_l159_129_6};
  assign _zz__zz_realValue_0_129 = {1'd0, wReg};
  assign _zz__zz_realValue_0_129_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_129_1 = (_zz_realValue_0_129_2 + _zz_realValue_0_129_3);
  assign _zz_realValue_0_129_2 = {1'd0, wReg};
  assign _zz_realValue_0_129_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_129_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_129 = {1'd0, _zz_when_ArraySlice_l166_129_1};
  assign _zz_when_ArraySlice_l166_129_2 = (_zz_when_ArraySlice_l166_129_3 + _zz_when_ArraySlice_l166_129_7);
  assign _zz_when_ArraySlice_l166_129_3 = (realValue_0_129 - _zz_when_ArraySlice_l166_129_4);
  assign _zz_when_ArraySlice_l166_129_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_129_5);
  assign _zz_when_ArraySlice_l166_129_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_129_5 = {3'd0, _zz_when_ArraySlice_l166_129_6};
  assign _zz_when_ArraySlice_l166_129_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_130 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_130_1);
  assign _zz_when_ArraySlice_l158_130_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_130_1 = {2'd0, _zz_when_ArraySlice_l158_130_2};
  assign _zz_when_ArraySlice_l158_130_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_130_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_130 = {1'd0, _zz_when_ArraySlice_l159_130_1};
  assign _zz_when_ArraySlice_l159_130_2 = (_zz_when_ArraySlice_l159_130_3 - _zz_when_ArraySlice_l159_130_4);
  assign _zz_when_ArraySlice_l159_130_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_130_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_130_5);
  assign _zz_when_ArraySlice_l159_130_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_130_5 = {2'd0, _zz_when_ArraySlice_l159_130_6};
  assign _zz__zz_realValue_0_130 = {1'd0, wReg};
  assign _zz__zz_realValue_0_130_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_130_1 = (_zz_realValue_0_130_2 + _zz_realValue_0_130_3);
  assign _zz_realValue_0_130_2 = {1'd0, wReg};
  assign _zz_realValue_0_130_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_130_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_130 = {1'd0, _zz_when_ArraySlice_l166_130_1};
  assign _zz_when_ArraySlice_l166_130_2 = (_zz_when_ArraySlice_l166_130_3 + _zz_when_ArraySlice_l166_130_7);
  assign _zz_when_ArraySlice_l166_130_3 = (realValue_0_130 - _zz_when_ArraySlice_l166_130_4);
  assign _zz_when_ArraySlice_l166_130_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_130_5);
  assign _zz_when_ArraySlice_l166_130_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_130_5 = {2'd0, _zz_when_ArraySlice_l166_130_6};
  assign _zz_when_ArraySlice_l166_130_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_131 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_131_1);
  assign _zz_when_ArraySlice_l158_131_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_131_1 = {2'd0, _zz_when_ArraySlice_l158_131_2};
  assign _zz_when_ArraySlice_l158_131_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_131_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_131 = {1'd0, _zz_when_ArraySlice_l159_131_1};
  assign _zz_when_ArraySlice_l159_131_2 = (_zz_when_ArraySlice_l159_131_3 - _zz_when_ArraySlice_l159_131_4);
  assign _zz_when_ArraySlice_l159_131_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_131_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_131_5);
  assign _zz_when_ArraySlice_l159_131_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_131_5 = {2'd0, _zz_when_ArraySlice_l159_131_6};
  assign _zz__zz_realValue_0_131 = {1'd0, wReg};
  assign _zz__zz_realValue_0_131_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_131_1 = (_zz_realValue_0_131_2 + _zz_realValue_0_131_3);
  assign _zz_realValue_0_131_2 = {1'd0, wReg};
  assign _zz_realValue_0_131_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_131_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_131 = {1'd0, _zz_when_ArraySlice_l166_131_1};
  assign _zz_when_ArraySlice_l166_131_2 = (_zz_when_ArraySlice_l166_131_3 + _zz_when_ArraySlice_l166_131_7);
  assign _zz_when_ArraySlice_l166_131_3 = (realValue_0_131 - _zz_when_ArraySlice_l166_131_4);
  assign _zz_when_ArraySlice_l166_131_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_131_5);
  assign _zz_when_ArraySlice_l166_131_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_131_5 = {2'd0, _zz_when_ArraySlice_l166_131_6};
  assign _zz_when_ArraySlice_l166_131_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_132 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_132_1);
  assign _zz_when_ArraySlice_l158_132_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_132_1 = {1'd0, _zz_when_ArraySlice_l158_132_2};
  assign _zz_when_ArraySlice_l158_132_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_132_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_132 = {1'd0, _zz_when_ArraySlice_l159_132_1};
  assign _zz_when_ArraySlice_l159_132_2 = (_zz_when_ArraySlice_l159_132_3 - _zz_when_ArraySlice_l159_132_4);
  assign _zz_when_ArraySlice_l159_132_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_132_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_132_5);
  assign _zz_when_ArraySlice_l159_132_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_132_5 = {1'd0, _zz_when_ArraySlice_l159_132_6};
  assign _zz__zz_realValue_0_132 = {1'd0, wReg};
  assign _zz__zz_realValue_0_132_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_132_1 = (_zz_realValue_0_132_2 + _zz_realValue_0_132_3);
  assign _zz_realValue_0_132_2 = {1'd0, wReg};
  assign _zz_realValue_0_132_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_132_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_132 = {1'd0, _zz_when_ArraySlice_l166_132_1};
  assign _zz_when_ArraySlice_l166_132_2 = (_zz_when_ArraySlice_l166_132_3 + _zz_when_ArraySlice_l166_132_7);
  assign _zz_when_ArraySlice_l166_132_3 = (realValue_0_132 - _zz_when_ArraySlice_l166_132_4);
  assign _zz_when_ArraySlice_l166_132_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_132_5);
  assign _zz_when_ArraySlice_l166_132_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_132_5 = {1'd0, _zz_when_ArraySlice_l166_132_6};
  assign _zz_when_ArraySlice_l166_132_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_133 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_133_1);
  assign _zz_when_ArraySlice_l158_133_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_133_1 = {1'd0, _zz_when_ArraySlice_l158_133_2};
  assign _zz_when_ArraySlice_l158_133_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_133_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_133 = {2'd0, _zz_when_ArraySlice_l159_133_1};
  assign _zz_when_ArraySlice_l159_133_2 = (_zz_when_ArraySlice_l159_133_3 - _zz_when_ArraySlice_l159_133_4);
  assign _zz_when_ArraySlice_l159_133_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_133_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_133_5);
  assign _zz_when_ArraySlice_l159_133_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_133_5 = {1'd0, _zz_when_ArraySlice_l159_133_6};
  assign _zz__zz_realValue_0_133 = {1'd0, wReg};
  assign _zz__zz_realValue_0_133_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_133_1 = (_zz_realValue_0_133_2 + _zz_realValue_0_133_3);
  assign _zz_realValue_0_133_2 = {1'd0, wReg};
  assign _zz_realValue_0_133_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_133_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_133 = {2'd0, _zz_when_ArraySlice_l166_133_1};
  assign _zz_when_ArraySlice_l166_133_2 = (_zz_when_ArraySlice_l166_133_3 + _zz_when_ArraySlice_l166_133_7);
  assign _zz_when_ArraySlice_l166_133_3 = (realValue_0_133 - _zz_when_ArraySlice_l166_133_4);
  assign _zz_when_ArraySlice_l166_133_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_133_5);
  assign _zz_when_ArraySlice_l166_133_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_133_5 = {1'd0, _zz_when_ArraySlice_l166_133_6};
  assign _zz_when_ArraySlice_l166_133_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_134 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_134_1);
  assign _zz_when_ArraySlice_l158_134_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_134_1 = {1'd0, _zz_when_ArraySlice_l158_134_2};
  assign _zz_when_ArraySlice_l158_134_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_134_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_134 = {2'd0, _zz_when_ArraySlice_l159_134_1};
  assign _zz_when_ArraySlice_l159_134_2 = (_zz_when_ArraySlice_l159_134_3 - _zz_when_ArraySlice_l159_134_4);
  assign _zz_when_ArraySlice_l159_134_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_134_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_134_5);
  assign _zz_when_ArraySlice_l159_134_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_134_5 = {1'd0, _zz_when_ArraySlice_l159_134_6};
  assign _zz__zz_realValue_0_134 = {1'd0, wReg};
  assign _zz__zz_realValue_0_134_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_134_1 = (_zz_realValue_0_134_2 + _zz_realValue_0_134_3);
  assign _zz_realValue_0_134_2 = {1'd0, wReg};
  assign _zz_realValue_0_134_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_134_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_134 = {2'd0, _zz_when_ArraySlice_l166_134_1};
  assign _zz_when_ArraySlice_l166_134_2 = (_zz_when_ArraySlice_l166_134_3 + _zz_when_ArraySlice_l166_134_7);
  assign _zz_when_ArraySlice_l166_134_3 = (realValue_0_134 - _zz_when_ArraySlice_l166_134_4);
  assign _zz_when_ArraySlice_l166_134_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_134_5);
  assign _zz_when_ArraySlice_l166_134_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_134_5 = {1'd0, _zz_when_ArraySlice_l166_134_6};
  assign _zz_when_ArraySlice_l166_134_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_135 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_135_1);
  assign _zz_when_ArraySlice_l158_135_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_135_1 = {1'd0, _zz_when_ArraySlice_l158_135_2};
  assign _zz_when_ArraySlice_l158_135_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_135_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_135 = {3'd0, _zz_when_ArraySlice_l159_135_1};
  assign _zz_when_ArraySlice_l159_135_2 = (_zz_when_ArraySlice_l159_135_3 - _zz_when_ArraySlice_l159_135_4);
  assign _zz_when_ArraySlice_l159_135_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_135_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_135_5);
  assign _zz_when_ArraySlice_l159_135_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_135_5 = {1'd0, _zz_when_ArraySlice_l159_135_6};
  assign _zz__zz_realValue_0_135 = {1'd0, wReg};
  assign _zz__zz_realValue_0_135_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_135_1 = (_zz_realValue_0_135_2 + _zz_realValue_0_135_3);
  assign _zz_realValue_0_135_2 = {1'd0, wReg};
  assign _zz_realValue_0_135_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_135_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_135 = {3'd0, _zz_when_ArraySlice_l166_135_1};
  assign _zz_when_ArraySlice_l166_135_2 = (_zz_when_ArraySlice_l166_135_3 + _zz_when_ArraySlice_l166_135_7);
  assign _zz_when_ArraySlice_l166_135_3 = (realValue_0_135 - _zz_when_ArraySlice_l166_135_4);
  assign _zz_when_ArraySlice_l166_135_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_135_5);
  assign _zz_when_ArraySlice_l166_135_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_135_5 = {1'd0, _zz_when_ArraySlice_l166_135_6};
  assign _zz_when_ArraySlice_l166_135_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_5_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_5_2 = (_zz_when_ArraySlice_l403_5_3 + _zz_when_ArraySlice_l403_5_7);
  assign _zz_when_ArraySlice_l403_5_3 = (_zz_when_ArraySlice_l403_5_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l403_5_5);
  assign _zz_when_ArraySlice_l403_5_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_5_5 = {1'd0, _zz_when_ArraySlice_l403_5_6};
  assign _zz_when_ArraySlice_l403_5_8 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l403_5_7 = {1'd0, _zz_when_ArraySlice_l403_5_8};
  assign _zz_when_ArraySlice_l406_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_5_1 = (_zz_when_ArraySlice_l406_5_2 + 8'h01);
  assign _zz_when_ArraySlice_l406_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l406_5_3);
  assign _zz_when_ArraySlice_l406_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_5_3 = {1'd0, _zz_when_ArraySlice_l406_5_4};
  assign _zz_selectReadFifo_5_6 = (selectReadFifo_5 + _zz_selectReadFifo_5_7);
  assign _zz_selectReadFifo_5_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_7 = {1'd0, _zz_selectReadFifo_5_8};
  assign _zz_when_ArraySlice_l413_5 = (_zz_when_ArraySlice_l413_5_1 % aReg);
  assign _zz_when_ArraySlice_l413_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l417_5_3);
  assign _zz_when_ArraySlice_l417_5_1 = _zz_when_ArraySlice_l417_5_2[6:0];
  assign _zz_when_ArraySlice_l417_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l417_5_3 = {1'd0, _zz_when_ArraySlice_l417_5_4};
  assign _zz_when_ArraySlice_l418_5_1 = (_zz_when_ArraySlice_l418_5_2 - _zz_when_ArraySlice_l418_5_3);
  assign _zz_when_ArraySlice_l418_5 = {5'd0, _zz_when_ArraySlice_l418_5_1};
  assign _zz_when_ArraySlice_l418_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l418_5_3 = {7'd0, _zz_when_ArraySlice_l418_5_4};
  assign _zz__zz_realValue1_0_16 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_16_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_16_1 = (_zz_realValue1_0_16_2 + _zz_realValue1_0_16_3);
  assign _zz_realValue1_0_16_2 = {1'd0, hReg};
  assign _zz_realValue1_0_16_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l420_5 = {1'd0, _zz_when_ArraySlice_l420_5_1};
  assign _zz_when_ArraySlice_l420_5_2 = (realValue1_0_16 / aReg);
  assign _zz_selectReadFifo_5_9 = (selectReadFifo_5 - _zz_selectReadFifo_5_10);
  assign _zz_selectReadFifo_5_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_136 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_136_1);
  assign _zz_when_ArraySlice_l158_136_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_136_1 = {4'd0, _zz_when_ArraySlice_l158_136_2};
  assign _zz_when_ArraySlice_l158_136_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_136 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_136_1 = (_zz_when_ArraySlice_l159_136_2 - _zz_when_ArraySlice_l159_136_3);
  assign _zz_when_ArraySlice_l159_136_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_136_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_136_4);
  assign _zz_when_ArraySlice_l159_136_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_136_4 = {4'd0, _zz_when_ArraySlice_l159_136_5};
  assign _zz__zz_realValue_0_136 = {1'd0, wReg};
  assign _zz__zz_realValue_0_136_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_136_1 = (_zz_realValue_0_136_2 + _zz_realValue_0_136_3);
  assign _zz_realValue_0_136_2 = {1'd0, wReg};
  assign _zz_realValue_0_136_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_136 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_136_1 = (_zz_when_ArraySlice_l166_136_2 + _zz_when_ArraySlice_l166_136_6);
  assign _zz_when_ArraySlice_l166_136_2 = (realValue_0_136 - _zz_when_ArraySlice_l166_136_3);
  assign _zz_when_ArraySlice_l166_136_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_136_4);
  assign _zz_when_ArraySlice_l166_136_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_136_4 = {4'd0, _zz_when_ArraySlice_l166_136_5};
  assign _zz_when_ArraySlice_l166_136_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_137 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_137_1);
  assign _zz_when_ArraySlice_l158_137_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_137_1 = {3'd0, _zz_when_ArraySlice_l158_137_2};
  assign _zz_when_ArraySlice_l158_137_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_137_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_137 = {1'd0, _zz_when_ArraySlice_l159_137_1};
  assign _zz_when_ArraySlice_l159_137_2 = (_zz_when_ArraySlice_l159_137_3 - _zz_when_ArraySlice_l159_137_4);
  assign _zz_when_ArraySlice_l159_137_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_137_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_137_5);
  assign _zz_when_ArraySlice_l159_137_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_137_5 = {3'd0, _zz_when_ArraySlice_l159_137_6};
  assign _zz__zz_realValue_0_137 = {1'd0, wReg};
  assign _zz__zz_realValue_0_137_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_137_1 = (_zz_realValue_0_137_2 + _zz_realValue_0_137_3);
  assign _zz_realValue_0_137_2 = {1'd0, wReg};
  assign _zz_realValue_0_137_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_137_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_137 = {1'd0, _zz_when_ArraySlice_l166_137_1};
  assign _zz_when_ArraySlice_l166_137_2 = (_zz_when_ArraySlice_l166_137_3 + _zz_when_ArraySlice_l166_137_7);
  assign _zz_when_ArraySlice_l166_137_3 = (realValue_0_137 - _zz_when_ArraySlice_l166_137_4);
  assign _zz_when_ArraySlice_l166_137_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_137_5);
  assign _zz_when_ArraySlice_l166_137_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_137_5 = {3'd0, _zz_when_ArraySlice_l166_137_6};
  assign _zz_when_ArraySlice_l166_137_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_138 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_138_1);
  assign _zz_when_ArraySlice_l158_138_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_138_1 = {2'd0, _zz_when_ArraySlice_l158_138_2};
  assign _zz_when_ArraySlice_l158_138_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_138_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_138 = {1'd0, _zz_when_ArraySlice_l159_138_1};
  assign _zz_when_ArraySlice_l159_138_2 = (_zz_when_ArraySlice_l159_138_3 - _zz_when_ArraySlice_l159_138_4);
  assign _zz_when_ArraySlice_l159_138_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_138_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_138_5);
  assign _zz_when_ArraySlice_l159_138_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_138_5 = {2'd0, _zz_when_ArraySlice_l159_138_6};
  assign _zz__zz_realValue_0_138 = {1'd0, wReg};
  assign _zz__zz_realValue_0_138_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_138_1 = (_zz_realValue_0_138_2 + _zz_realValue_0_138_3);
  assign _zz_realValue_0_138_2 = {1'd0, wReg};
  assign _zz_realValue_0_138_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_138_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_138 = {1'd0, _zz_when_ArraySlice_l166_138_1};
  assign _zz_when_ArraySlice_l166_138_2 = (_zz_when_ArraySlice_l166_138_3 + _zz_when_ArraySlice_l166_138_7);
  assign _zz_when_ArraySlice_l166_138_3 = (realValue_0_138 - _zz_when_ArraySlice_l166_138_4);
  assign _zz_when_ArraySlice_l166_138_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_138_5);
  assign _zz_when_ArraySlice_l166_138_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_138_5 = {2'd0, _zz_when_ArraySlice_l166_138_6};
  assign _zz_when_ArraySlice_l166_138_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_139 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_139_1);
  assign _zz_when_ArraySlice_l158_139_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_139_1 = {2'd0, _zz_when_ArraySlice_l158_139_2};
  assign _zz_when_ArraySlice_l158_139_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_139_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_139 = {1'd0, _zz_when_ArraySlice_l159_139_1};
  assign _zz_when_ArraySlice_l159_139_2 = (_zz_when_ArraySlice_l159_139_3 - _zz_when_ArraySlice_l159_139_4);
  assign _zz_when_ArraySlice_l159_139_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_139_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_139_5);
  assign _zz_when_ArraySlice_l159_139_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_139_5 = {2'd0, _zz_when_ArraySlice_l159_139_6};
  assign _zz__zz_realValue_0_139 = {1'd0, wReg};
  assign _zz__zz_realValue_0_139_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_139_1 = (_zz_realValue_0_139_2 + _zz_realValue_0_139_3);
  assign _zz_realValue_0_139_2 = {1'd0, wReg};
  assign _zz_realValue_0_139_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_139_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_139 = {1'd0, _zz_when_ArraySlice_l166_139_1};
  assign _zz_when_ArraySlice_l166_139_2 = (_zz_when_ArraySlice_l166_139_3 + _zz_when_ArraySlice_l166_139_7);
  assign _zz_when_ArraySlice_l166_139_3 = (realValue_0_139 - _zz_when_ArraySlice_l166_139_4);
  assign _zz_when_ArraySlice_l166_139_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_139_5);
  assign _zz_when_ArraySlice_l166_139_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_139_5 = {2'd0, _zz_when_ArraySlice_l166_139_6};
  assign _zz_when_ArraySlice_l166_139_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_140 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_140_1);
  assign _zz_when_ArraySlice_l158_140_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_140_1 = {1'd0, _zz_when_ArraySlice_l158_140_2};
  assign _zz_when_ArraySlice_l158_140_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_140_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_140 = {1'd0, _zz_when_ArraySlice_l159_140_1};
  assign _zz_when_ArraySlice_l159_140_2 = (_zz_when_ArraySlice_l159_140_3 - _zz_when_ArraySlice_l159_140_4);
  assign _zz_when_ArraySlice_l159_140_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_140_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_140_5);
  assign _zz_when_ArraySlice_l159_140_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_140_5 = {1'd0, _zz_when_ArraySlice_l159_140_6};
  assign _zz__zz_realValue_0_140 = {1'd0, wReg};
  assign _zz__zz_realValue_0_140_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_140_1 = (_zz_realValue_0_140_2 + _zz_realValue_0_140_3);
  assign _zz_realValue_0_140_2 = {1'd0, wReg};
  assign _zz_realValue_0_140_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_140_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_140 = {1'd0, _zz_when_ArraySlice_l166_140_1};
  assign _zz_when_ArraySlice_l166_140_2 = (_zz_when_ArraySlice_l166_140_3 + _zz_when_ArraySlice_l166_140_7);
  assign _zz_when_ArraySlice_l166_140_3 = (realValue_0_140 - _zz_when_ArraySlice_l166_140_4);
  assign _zz_when_ArraySlice_l166_140_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_140_5);
  assign _zz_when_ArraySlice_l166_140_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_140_5 = {1'd0, _zz_when_ArraySlice_l166_140_6};
  assign _zz_when_ArraySlice_l166_140_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_141 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_141_1);
  assign _zz_when_ArraySlice_l158_141_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_141_1 = {1'd0, _zz_when_ArraySlice_l158_141_2};
  assign _zz_when_ArraySlice_l158_141_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_141_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_141 = {2'd0, _zz_when_ArraySlice_l159_141_1};
  assign _zz_when_ArraySlice_l159_141_2 = (_zz_when_ArraySlice_l159_141_3 - _zz_when_ArraySlice_l159_141_4);
  assign _zz_when_ArraySlice_l159_141_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_141_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_141_5);
  assign _zz_when_ArraySlice_l159_141_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_141_5 = {1'd0, _zz_when_ArraySlice_l159_141_6};
  assign _zz__zz_realValue_0_141 = {1'd0, wReg};
  assign _zz__zz_realValue_0_141_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_141_1 = (_zz_realValue_0_141_2 + _zz_realValue_0_141_3);
  assign _zz_realValue_0_141_2 = {1'd0, wReg};
  assign _zz_realValue_0_141_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_141_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_141 = {2'd0, _zz_when_ArraySlice_l166_141_1};
  assign _zz_when_ArraySlice_l166_141_2 = (_zz_when_ArraySlice_l166_141_3 + _zz_when_ArraySlice_l166_141_7);
  assign _zz_when_ArraySlice_l166_141_3 = (realValue_0_141 - _zz_when_ArraySlice_l166_141_4);
  assign _zz_when_ArraySlice_l166_141_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_141_5);
  assign _zz_when_ArraySlice_l166_141_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_141_5 = {1'd0, _zz_when_ArraySlice_l166_141_6};
  assign _zz_when_ArraySlice_l166_141_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_142 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_142_1);
  assign _zz_when_ArraySlice_l158_142_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_142_1 = {1'd0, _zz_when_ArraySlice_l158_142_2};
  assign _zz_when_ArraySlice_l158_142_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_142_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_142 = {2'd0, _zz_when_ArraySlice_l159_142_1};
  assign _zz_when_ArraySlice_l159_142_2 = (_zz_when_ArraySlice_l159_142_3 - _zz_when_ArraySlice_l159_142_4);
  assign _zz_when_ArraySlice_l159_142_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_142_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_142_5);
  assign _zz_when_ArraySlice_l159_142_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_142_5 = {1'd0, _zz_when_ArraySlice_l159_142_6};
  assign _zz__zz_realValue_0_142 = {1'd0, wReg};
  assign _zz__zz_realValue_0_142_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_142_1 = (_zz_realValue_0_142_2 + _zz_realValue_0_142_3);
  assign _zz_realValue_0_142_2 = {1'd0, wReg};
  assign _zz_realValue_0_142_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_142_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_142 = {2'd0, _zz_when_ArraySlice_l166_142_1};
  assign _zz_when_ArraySlice_l166_142_2 = (_zz_when_ArraySlice_l166_142_3 + _zz_when_ArraySlice_l166_142_7);
  assign _zz_when_ArraySlice_l166_142_3 = (realValue_0_142 - _zz_when_ArraySlice_l166_142_4);
  assign _zz_when_ArraySlice_l166_142_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_142_5);
  assign _zz_when_ArraySlice_l166_142_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_142_5 = {1'd0, _zz_when_ArraySlice_l166_142_6};
  assign _zz_when_ArraySlice_l166_142_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_143 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_143_1);
  assign _zz_when_ArraySlice_l158_143_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_143_1 = {1'd0, _zz_when_ArraySlice_l158_143_2};
  assign _zz_when_ArraySlice_l158_143_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_143_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_143 = {3'd0, _zz_when_ArraySlice_l159_143_1};
  assign _zz_when_ArraySlice_l159_143_2 = (_zz_when_ArraySlice_l159_143_3 - _zz_when_ArraySlice_l159_143_4);
  assign _zz_when_ArraySlice_l159_143_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_143_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_143_5);
  assign _zz_when_ArraySlice_l159_143_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_143_5 = {1'd0, _zz_when_ArraySlice_l159_143_6};
  assign _zz__zz_realValue_0_143 = {1'd0, wReg};
  assign _zz__zz_realValue_0_143_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_143_1 = (_zz_realValue_0_143_2 + _zz_realValue_0_143_3);
  assign _zz_realValue_0_143_2 = {1'd0, wReg};
  assign _zz_realValue_0_143_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_143_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_143 = {3'd0, _zz_when_ArraySlice_l166_143_1};
  assign _zz_when_ArraySlice_l166_143_2 = (_zz_when_ArraySlice_l166_143_3 + _zz_when_ArraySlice_l166_143_7);
  assign _zz_when_ArraySlice_l166_143_3 = (realValue_0_143 - _zz_when_ArraySlice_l166_143_4);
  assign _zz_when_ArraySlice_l166_143_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_143_5);
  assign _zz_when_ArraySlice_l166_143_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_143_5 = {1'd0, _zz_when_ArraySlice_l166_143_6};
  assign _zz_when_ArraySlice_l166_143_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_5_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_5_2 = (_zz_when_ArraySlice_l428_5_3 + _zz_when_ArraySlice_l428_5_7);
  assign _zz_when_ArraySlice_l428_5_3 = (_zz_when_ArraySlice_l428_5_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l428_5_5);
  assign _zz_when_ArraySlice_l428_5_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_5_5 = {1'd0, _zz_when_ArraySlice_l428_5_6};
  assign _zz_when_ArraySlice_l428_5_8 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l428_5_7 = {1'd0, _zz_when_ArraySlice_l428_5_8};
  assign _zz_when_ArraySlice_l431_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_5_1 = (_zz_when_ArraySlice_l431_5_2 + 8'h01);
  assign _zz_when_ArraySlice_l431_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l431_5_3);
  assign _zz_when_ArraySlice_l431_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_5_3 = {1'd0, _zz_when_ArraySlice_l431_5_4};
  assign _zz_selectReadFifo_5_11 = (selectReadFifo_5 + _zz_selectReadFifo_5_12);
  assign _zz_selectReadFifo_5_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_12 = {1'd0, _zz_selectReadFifo_5_13};
  assign _zz_when_ArraySlice_l438_5 = (_zz_when_ArraySlice_l438_5_1 % aReg);
  assign _zz_when_ArraySlice_l438_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_5_1 = (_zz_when_ArraySlice_l449_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l449_5 = {5'd0, _zz_when_ArraySlice_l449_5_1};
  assign _zz_when_ArraySlice_l449_5_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_17 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_17_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_17_1 = (_zz_realValue1_0_17_2 + _zz_realValue1_0_17_3);
  assign _zz_realValue1_0_17_2 = {1'd0, hReg};
  assign _zz_realValue1_0_17_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l450_5 = {1'd0, _zz_when_ArraySlice_l450_5_1};
  assign _zz_when_ArraySlice_l450_5_2 = (realValue1_0_17 / aReg);
  assign _zz_selectReadFifo_5_14 = (selectReadFifo_5 - _zz_selectReadFifo_5_15);
  assign _zz_selectReadFifo_5_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_144 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_144_1);
  assign _zz_when_ArraySlice_l158_144_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_144_1 = {4'd0, _zz_when_ArraySlice_l158_144_2};
  assign _zz_when_ArraySlice_l158_144_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_144 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_144_1 = (_zz_when_ArraySlice_l159_144_2 - _zz_when_ArraySlice_l159_144_3);
  assign _zz_when_ArraySlice_l159_144_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_144_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_144_4);
  assign _zz_when_ArraySlice_l159_144_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_144_4 = {4'd0, _zz_when_ArraySlice_l159_144_5};
  assign _zz__zz_realValue_0_144 = {1'd0, wReg};
  assign _zz__zz_realValue_0_144_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_144_1 = (_zz_realValue_0_144_2 + _zz_realValue_0_144_3);
  assign _zz_realValue_0_144_2 = {1'd0, wReg};
  assign _zz_realValue_0_144_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_144 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_144_1 = (_zz_when_ArraySlice_l166_144_2 + _zz_when_ArraySlice_l166_144_6);
  assign _zz_when_ArraySlice_l166_144_2 = (realValue_0_144 - _zz_when_ArraySlice_l166_144_3);
  assign _zz_when_ArraySlice_l166_144_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_144_4);
  assign _zz_when_ArraySlice_l166_144_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_144_4 = {4'd0, _zz_when_ArraySlice_l166_144_5};
  assign _zz_when_ArraySlice_l166_144_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_145 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_145_1);
  assign _zz_when_ArraySlice_l158_145_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_145_1 = {3'd0, _zz_when_ArraySlice_l158_145_2};
  assign _zz_when_ArraySlice_l158_145_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_145_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_145 = {1'd0, _zz_when_ArraySlice_l159_145_1};
  assign _zz_when_ArraySlice_l159_145_2 = (_zz_when_ArraySlice_l159_145_3 - _zz_when_ArraySlice_l159_145_4);
  assign _zz_when_ArraySlice_l159_145_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_145_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_145_5);
  assign _zz_when_ArraySlice_l159_145_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_145_5 = {3'd0, _zz_when_ArraySlice_l159_145_6};
  assign _zz__zz_realValue_0_145 = {1'd0, wReg};
  assign _zz__zz_realValue_0_145_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_145_1 = (_zz_realValue_0_145_2 + _zz_realValue_0_145_3);
  assign _zz_realValue_0_145_2 = {1'd0, wReg};
  assign _zz_realValue_0_145_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_145_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_145 = {1'd0, _zz_when_ArraySlice_l166_145_1};
  assign _zz_when_ArraySlice_l166_145_2 = (_zz_when_ArraySlice_l166_145_3 + _zz_when_ArraySlice_l166_145_7);
  assign _zz_when_ArraySlice_l166_145_3 = (realValue_0_145 - _zz_when_ArraySlice_l166_145_4);
  assign _zz_when_ArraySlice_l166_145_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_145_5);
  assign _zz_when_ArraySlice_l166_145_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_145_5 = {3'd0, _zz_when_ArraySlice_l166_145_6};
  assign _zz_when_ArraySlice_l166_145_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_146 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_146_1);
  assign _zz_when_ArraySlice_l158_146_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_146_1 = {2'd0, _zz_when_ArraySlice_l158_146_2};
  assign _zz_when_ArraySlice_l158_146_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_146_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_146 = {1'd0, _zz_when_ArraySlice_l159_146_1};
  assign _zz_when_ArraySlice_l159_146_2 = (_zz_when_ArraySlice_l159_146_3 - _zz_when_ArraySlice_l159_146_4);
  assign _zz_when_ArraySlice_l159_146_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_146_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_146_5);
  assign _zz_when_ArraySlice_l159_146_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_146_5 = {2'd0, _zz_when_ArraySlice_l159_146_6};
  assign _zz__zz_realValue_0_146 = {1'd0, wReg};
  assign _zz__zz_realValue_0_146_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_146_1 = (_zz_realValue_0_146_2 + _zz_realValue_0_146_3);
  assign _zz_realValue_0_146_2 = {1'd0, wReg};
  assign _zz_realValue_0_146_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_146_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_146 = {1'd0, _zz_when_ArraySlice_l166_146_1};
  assign _zz_when_ArraySlice_l166_146_2 = (_zz_when_ArraySlice_l166_146_3 + _zz_when_ArraySlice_l166_146_7);
  assign _zz_when_ArraySlice_l166_146_3 = (realValue_0_146 - _zz_when_ArraySlice_l166_146_4);
  assign _zz_when_ArraySlice_l166_146_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_146_5);
  assign _zz_when_ArraySlice_l166_146_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_146_5 = {2'd0, _zz_when_ArraySlice_l166_146_6};
  assign _zz_when_ArraySlice_l166_146_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_147 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_147_1);
  assign _zz_when_ArraySlice_l158_147_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_147_1 = {2'd0, _zz_when_ArraySlice_l158_147_2};
  assign _zz_when_ArraySlice_l158_147_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_147_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_147 = {1'd0, _zz_when_ArraySlice_l159_147_1};
  assign _zz_when_ArraySlice_l159_147_2 = (_zz_when_ArraySlice_l159_147_3 - _zz_when_ArraySlice_l159_147_4);
  assign _zz_when_ArraySlice_l159_147_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_147_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_147_5);
  assign _zz_when_ArraySlice_l159_147_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_147_5 = {2'd0, _zz_when_ArraySlice_l159_147_6};
  assign _zz__zz_realValue_0_147 = {1'd0, wReg};
  assign _zz__zz_realValue_0_147_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_147_1 = (_zz_realValue_0_147_2 + _zz_realValue_0_147_3);
  assign _zz_realValue_0_147_2 = {1'd0, wReg};
  assign _zz_realValue_0_147_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_147_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_147 = {1'd0, _zz_when_ArraySlice_l166_147_1};
  assign _zz_when_ArraySlice_l166_147_2 = (_zz_when_ArraySlice_l166_147_3 + _zz_when_ArraySlice_l166_147_7);
  assign _zz_when_ArraySlice_l166_147_3 = (realValue_0_147 - _zz_when_ArraySlice_l166_147_4);
  assign _zz_when_ArraySlice_l166_147_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_147_5);
  assign _zz_when_ArraySlice_l166_147_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_147_5 = {2'd0, _zz_when_ArraySlice_l166_147_6};
  assign _zz_when_ArraySlice_l166_147_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_148 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_148_1);
  assign _zz_when_ArraySlice_l158_148_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_148_1 = {1'd0, _zz_when_ArraySlice_l158_148_2};
  assign _zz_when_ArraySlice_l158_148_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_148_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_148 = {1'd0, _zz_when_ArraySlice_l159_148_1};
  assign _zz_when_ArraySlice_l159_148_2 = (_zz_when_ArraySlice_l159_148_3 - _zz_when_ArraySlice_l159_148_4);
  assign _zz_when_ArraySlice_l159_148_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_148_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_148_5);
  assign _zz_when_ArraySlice_l159_148_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_148_5 = {1'd0, _zz_when_ArraySlice_l159_148_6};
  assign _zz__zz_realValue_0_148 = {1'd0, wReg};
  assign _zz__zz_realValue_0_148_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_148_1 = (_zz_realValue_0_148_2 + _zz_realValue_0_148_3);
  assign _zz_realValue_0_148_2 = {1'd0, wReg};
  assign _zz_realValue_0_148_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_148_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_148 = {1'd0, _zz_when_ArraySlice_l166_148_1};
  assign _zz_when_ArraySlice_l166_148_2 = (_zz_when_ArraySlice_l166_148_3 + _zz_when_ArraySlice_l166_148_7);
  assign _zz_when_ArraySlice_l166_148_3 = (realValue_0_148 - _zz_when_ArraySlice_l166_148_4);
  assign _zz_when_ArraySlice_l166_148_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_148_5);
  assign _zz_when_ArraySlice_l166_148_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_148_5 = {1'd0, _zz_when_ArraySlice_l166_148_6};
  assign _zz_when_ArraySlice_l166_148_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_149 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_149_1);
  assign _zz_when_ArraySlice_l158_149_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_149_1 = {1'd0, _zz_when_ArraySlice_l158_149_2};
  assign _zz_when_ArraySlice_l158_149_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_149_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_149 = {2'd0, _zz_when_ArraySlice_l159_149_1};
  assign _zz_when_ArraySlice_l159_149_2 = (_zz_when_ArraySlice_l159_149_3 - _zz_when_ArraySlice_l159_149_4);
  assign _zz_when_ArraySlice_l159_149_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_149_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_149_5);
  assign _zz_when_ArraySlice_l159_149_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_149_5 = {1'd0, _zz_when_ArraySlice_l159_149_6};
  assign _zz__zz_realValue_0_149 = {1'd0, wReg};
  assign _zz__zz_realValue_0_149_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_149_1 = (_zz_realValue_0_149_2 + _zz_realValue_0_149_3);
  assign _zz_realValue_0_149_2 = {1'd0, wReg};
  assign _zz_realValue_0_149_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_149_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_149 = {2'd0, _zz_when_ArraySlice_l166_149_1};
  assign _zz_when_ArraySlice_l166_149_2 = (_zz_when_ArraySlice_l166_149_3 + _zz_when_ArraySlice_l166_149_7);
  assign _zz_when_ArraySlice_l166_149_3 = (realValue_0_149 - _zz_when_ArraySlice_l166_149_4);
  assign _zz_when_ArraySlice_l166_149_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_149_5);
  assign _zz_when_ArraySlice_l166_149_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_149_5 = {1'd0, _zz_when_ArraySlice_l166_149_6};
  assign _zz_when_ArraySlice_l166_149_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_150 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_150_1);
  assign _zz_when_ArraySlice_l158_150_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_150_1 = {1'd0, _zz_when_ArraySlice_l158_150_2};
  assign _zz_when_ArraySlice_l158_150_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_150_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_150 = {2'd0, _zz_when_ArraySlice_l159_150_1};
  assign _zz_when_ArraySlice_l159_150_2 = (_zz_when_ArraySlice_l159_150_3 - _zz_when_ArraySlice_l159_150_4);
  assign _zz_when_ArraySlice_l159_150_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_150_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_150_5);
  assign _zz_when_ArraySlice_l159_150_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_150_5 = {1'd0, _zz_when_ArraySlice_l159_150_6};
  assign _zz__zz_realValue_0_150 = {1'd0, wReg};
  assign _zz__zz_realValue_0_150_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_150_1 = (_zz_realValue_0_150_2 + _zz_realValue_0_150_3);
  assign _zz_realValue_0_150_2 = {1'd0, wReg};
  assign _zz_realValue_0_150_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_150_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_150 = {2'd0, _zz_when_ArraySlice_l166_150_1};
  assign _zz_when_ArraySlice_l166_150_2 = (_zz_when_ArraySlice_l166_150_3 + _zz_when_ArraySlice_l166_150_7);
  assign _zz_when_ArraySlice_l166_150_3 = (realValue_0_150 - _zz_when_ArraySlice_l166_150_4);
  assign _zz_when_ArraySlice_l166_150_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_150_5);
  assign _zz_when_ArraySlice_l166_150_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_150_5 = {1'd0, _zz_when_ArraySlice_l166_150_6};
  assign _zz_when_ArraySlice_l166_150_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_151 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_151_1);
  assign _zz_when_ArraySlice_l158_151_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_151_1 = {1'd0, _zz_when_ArraySlice_l158_151_2};
  assign _zz_when_ArraySlice_l158_151_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_151_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_151 = {3'd0, _zz_when_ArraySlice_l159_151_1};
  assign _zz_when_ArraySlice_l159_151_2 = (_zz_when_ArraySlice_l159_151_3 - _zz_when_ArraySlice_l159_151_4);
  assign _zz_when_ArraySlice_l159_151_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_151_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_151_5);
  assign _zz_when_ArraySlice_l159_151_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_151_5 = {1'd0, _zz_when_ArraySlice_l159_151_6};
  assign _zz__zz_realValue_0_151 = {1'd0, wReg};
  assign _zz__zz_realValue_0_151_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_151_1 = (_zz_realValue_0_151_2 + _zz_realValue_0_151_3);
  assign _zz_realValue_0_151_2 = {1'd0, wReg};
  assign _zz_realValue_0_151_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_151_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_151 = {3'd0, _zz_when_ArraySlice_l166_151_1};
  assign _zz_when_ArraySlice_l166_151_2 = (_zz_when_ArraySlice_l166_151_3 + _zz_when_ArraySlice_l166_151_7);
  assign _zz_when_ArraySlice_l166_151_3 = (realValue_0_151 - _zz_when_ArraySlice_l166_151_4);
  assign _zz_when_ArraySlice_l166_151_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_151_5);
  assign _zz_when_ArraySlice_l166_151_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_151_5 = {1'd0, _zz_when_ArraySlice_l166_151_6};
  assign _zz_when_ArraySlice_l166_151_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_5 = (_zz_when_ArraySlice_l461_5_1 % aReg);
  assign _zz_when_ArraySlice_l461_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l447_5_2);
  assign _zz_when_ArraySlice_l447_5_3 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l447_5_2 = {1'd0, _zz_when_ArraySlice_l447_5_3};
  assign _zz_when_ArraySlice_l468_5_1 = (_zz_when_ArraySlice_l468_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l468_5 = {5'd0, _zz_when_ArraySlice_l468_5_1};
  assign _zz_when_ArraySlice_l468_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l376_6_1);
  assign _zz_when_ArraySlice_l376_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l376_6_1 = {1'd0, _zz_when_ArraySlice_l376_6_2};
  assign _zz_when_ArraySlice_l376_6_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l377_6_3);
  assign _zz_when_ArraySlice_l377_6_1 = _zz_when_ArraySlice_l377_6_2[6:0];
  assign _zz_when_ArraySlice_l377_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l377_6_3 = {1'd0, _zz_when_ArraySlice_l377_6_4};
  assign _zz__zz_outputStreamArrayData_6_valid_1 = (bReg * 3'b110);
  assign _zz__zz_outputStreamArrayData_6_valid = {1'd0, _zz__zz_outputStreamArrayData_6_valid_1};
  assign _zz__zz_9 = _zz_outputStreamArrayData_6_valid[6:0];
  assign _zz_outputStreamArrayData_6_valid_3 = _zz_outputStreamArrayData_6_valid[6:0];
  assign _zz_outputStreamArrayData_6_payload_1 = _zz_outputStreamArrayData_6_valid[6:0];
  assign _zz_when_ArraySlice_l383_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l383_6_3);
  assign _zz_when_ArraySlice_l383_6_1 = _zz_when_ArraySlice_l383_6_2[6:0];
  assign _zz_when_ArraySlice_l383_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l383_6_3 = {1'd0, _zz_when_ArraySlice_l383_6_4};
  assign _zz_when_ArraySlice_l384_6_1 = (_zz_when_ArraySlice_l384_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l384_6 = {5'd0, _zz_when_ArraySlice_l384_6_1};
  assign _zz_when_ArraySlice_l384_6_2 = (bReg * aReg);
  assign _zz_selectReadFifo_6 = (selectReadFifo_6 - _zz_selectReadFifo_6_1);
  assign _zz_selectReadFifo_6_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_6 = (_zz_when_ArraySlice_l387_6_1 % aReg);
  assign _zz_when_ArraySlice_l387_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l392_6_3);
  assign _zz_when_ArraySlice_l392_6_1 = _zz_when_ArraySlice_l392_6_2[6:0];
  assign _zz_when_ArraySlice_l392_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l392_6_3 = {1'd0, _zz_when_ArraySlice_l392_6_4};
  assign _zz_when_ArraySlice_l393_6_1 = (_zz_when_ArraySlice_l393_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l393_6 = {5'd0, _zz_when_ArraySlice_l393_6_1};
  assign _zz_when_ArraySlice_l393_6_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_18 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_18_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_18_1 = (_zz_realValue1_0_18_2 + _zz_realValue1_0_18_3);
  assign _zz_realValue1_0_18_2 = {1'd0, hReg};
  assign _zz_realValue1_0_18_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l395_6 = {1'd0, _zz_when_ArraySlice_l395_6_1};
  assign _zz_when_ArraySlice_l395_6_2 = (realValue1_0_18 / aReg);
  assign _zz_selectReadFifo_6_2 = (selectReadFifo_6 - _zz_selectReadFifo_6_3);
  assign _zz_selectReadFifo_6_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_6_5 = 1'b1;
  assign _zz_selectReadFifo_6_4 = {7'd0, _zz_selectReadFifo_6_5};
  assign _zz_when_ArraySlice_l158_152 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_152_1);
  assign _zz_when_ArraySlice_l158_152_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_152_1 = {4'd0, _zz_when_ArraySlice_l158_152_2};
  assign _zz_when_ArraySlice_l158_152_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_152 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_152_1 = (_zz_when_ArraySlice_l159_152_2 - _zz_when_ArraySlice_l159_152_3);
  assign _zz_when_ArraySlice_l159_152_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_152_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_152_4);
  assign _zz_when_ArraySlice_l159_152_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_152_4 = {4'd0, _zz_when_ArraySlice_l159_152_5};
  assign _zz__zz_realValue_0_152 = {1'd0, wReg};
  assign _zz__zz_realValue_0_152_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_152_1 = (_zz_realValue_0_152_2 + _zz_realValue_0_152_3);
  assign _zz_realValue_0_152_2 = {1'd0, wReg};
  assign _zz_realValue_0_152_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_152 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_152_1 = (_zz_when_ArraySlice_l166_152_2 + _zz_when_ArraySlice_l166_152_6);
  assign _zz_when_ArraySlice_l166_152_2 = (realValue_0_152 - _zz_when_ArraySlice_l166_152_3);
  assign _zz_when_ArraySlice_l166_152_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_152_4);
  assign _zz_when_ArraySlice_l166_152_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_152_4 = {4'd0, _zz_when_ArraySlice_l166_152_5};
  assign _zz_when_ArraySlice_l166_152_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_153 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_153_1);
  assign _zz_when_ArraySlice_l158_153_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_153_1 = {3'd0, _zz_when_ArraySlice_l158_153_2};
  assign _zz_when_ArraySlice_l158_153_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_153_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_153 = {1'd0, _zz_when_ArraySlice_l159_153_1};
  assign _zz_when_ArraySlice_l159_153_2 = (_zz_when_ArraySlice_l159_153_3 - _zz_when_ArraySlice_l159_153_4);
  assign _zz_when_ArraySlice_l159_153_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_153_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_153_5);
  assign _zz_when_ArraySlice_l159_153_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_153_5 = {3'd0, _zz_when_ArraySlice_l159_153_6};
  assign _zz__zz_realValue_0_153 = {1'd0, wReg};
  assign _zz__zz_realValue_0_153_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_153_1 = (_zz_realValue_0_153_2 + _zz_realValue_0_153_3);
  assign _zz_realValue_0_153_2 = {1'd0, wReg};
  assign _zz_realValue_0_153_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_153_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_153 = {1'd0, _zz_when_ArraySlice_l166_153_1};
  assign _zz_when_ArraySlice_l166_153_2 = (_zz_when_ArraySlice_l166_153_3 + _zz_when_ArraySlice_l166_153_7);
  assign _zz_when_ArraySlice_l166_153_3 = (realValue_0_153 - _zz_when_ArraySlice_l166_153_4);
  assign _zz_when_ArraySlice_l166_153_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_153_5);
  assign _zz_when_ArraySlice_l166_153_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_153_5 = {3'd0, _zz_when_ArraySlice_l166_153_6};
  assign _zz_when_ArraySlice_l166_153_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_154 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_154_1);
  assign _zz_when_ArraySlice_l158_154_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_154_1 = {2'd0, _zz_when_ArraySlice_l158_154_2};
  assign _zz_when_ArraySlice_l158_154_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_154_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_154 = {1'd0, _zz_when_ArraySlice_l159_154_1};
  assign _zz_when_ArraySlice_l159_154_2 = (_zz_when_ArraySlice_l159_154_3 - _zz_when_ArraySlice_l159_154_4);
  assign _zz_when_ArraySlice_l159_154_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_154_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_154_5);
  assign _zz_when_ArraySlice_l159_154_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_154_5 = {2'd0, _zz_when_ArraySlice_l159_154_6};
  assign _zz__zz_realValue_0_154 = {1'd0, wReg};
  assign _zz__zz_realValue_0_154_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_154_1 = (_zz_realValue_0_154_2 + _zz_realValue_0_154_3);
  assign _zz_realValue_0_154_2 = {1'd0, wReg};
  assign _zz_realValue_0_154_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_154_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_154 = {1'd0, _zz_when_ArraySlice_l166_154_1};
  assign _zz_when_ArraySlice_l166_154_2 = (_zz_when_ArraySlice_l166_154_3 + _zz_when_ArraySlice_l166_154_7);
  assign _zz_when_ArraySlice_l166_154_3 = (realValue_0_154 - _zz_when_ArraySlice_l166_154_4);
  assign _zz_when_ArraySlice_l166_154_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_154_5);
  assign _zz_when_ArraySlice_l166_154_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_154_5 = {2'd0, _zz_when_ArraySlice_l166_154_6};
  assign _zz_when_ArraySlice_l166_154_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_155 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_155_1);
  assign _zz_when_ArraySlice_l158_155_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_155_1 = {2'd0, _zz_when_ArraySlice_l158_155_2};
  assign _zz_when_ArraySlice_l158_155_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_155_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_155 = {1'd0, _zz_when_ArraySlice_l159_155_1};
  assign _zz_when_ArraySlice_l159_155_2 = (_zz_when_ArraySlice_l159_155_3 - _zz_when_ArraySlice_l159_155_4);
  assign _zz_when_ArraySlice_l159_155_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_155_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_155_5);
  assign _zz_when_ArraySlice_l159_155_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_155_5 = {2'd0, _zz_when_ArraySlice_l159_155_6};
  assign _zz__zz_realValue_0_155 = {1'd0, wReg};
  assign _zz__zz_realValue_0_155_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_155_1 = (_zz_realValue_0_155_2 + _zz_realValue_0_155_3);
  assign _zz_realValue_0_155_2 = {1'd0, wReg};
  assign _zz_realValue_0_155_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_155_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_155 = {1'd0, _zz_when_ArraySlice_l166_155_1};
  assign _zz_when_ArraySlice_l166_155_2 = (_zz_when_ArraySlice_l166_155_3 + _zz_when_ArraySlice_l166_155_7);
  assign _zz_when_ArraySlice_l166_155_3 = (realValue_0_155 - _zz_when_ArraySlice_l166_155_4);
  assign _zz_when_ArraySlice_l166_155_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_155_5);
  assign _zz_when_ArraySlice_l166_155_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_155_5 = {2'd0, _zz_when_ArraySlice_l166_155_6};
  assign _zz_when_ArraySlice_l166_155_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_156 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_156_1);
  assign _zz_when_ArraySlice_l158_156_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_156_1 = {1'd0, _zz_when_ArraySlice_l158_156_2};
  assign _zz_when_ArraySlice_l158_156_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_156_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_156 = {1'd0, _zz_when_ArraySlice_l159_156_1};
  assign _zz_when_ArraySlice_l159_156_2 = (_zz_when_ArraySlice_l159_156_3 - _zz_when_ArraySlice_l159_156_4);
  assign _zz_when_ArraySlice_l159_156_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_156_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_156_5);
  assign _zz_when_ArraySlice_l159_156_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_156_5 = {1'd0, _zz_when_ArraySlice_l159_156_6};
  assign _zz__zz_realValue_0_156 = {1'd0, wReg};
  assign _zz__zz_realValue_0_156_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_156_1 = (_zz_realValue_0_156_2 + _zz_realValue_0_156_3);
  assign _zz_realValue_0_156_2 = {1'd0, wReg};
  assign _zz_realValue_0_156_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_156_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_156 = {1'd0, _zz_when_ArraySlice_l166_156_1};
  assign _zz_when_ArraySlice_l166_156_2 = (_zz_when_ArraySlice_l166_156_3 + _zz_when_ArraySlice_l166_156_7);
  assign _zz_when_ArraySlice_l166_156_3 = (realValue_0_156 - _zz_when_ArraySlice_l166_156_4);
  assign _zz_when_ArraySlice_l166_156_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_156_5);
  assign _zz_when_ArraySlice_l166_156_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_156_5 = {1'd0, _zz_when_ArraySlice_l166_156_6};
  assign _zz_when_ArraySlice_l166_156_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_157 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_157_1);
  assign _zz_when_ArraySlice_l158_157_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_157_1 = {1'd0, _zz_when_ArraySlice_l158_157_2};
  assign _zz_when_ArraySlice_l158_157_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_157_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_157 = {2'd0, _zz_when_ArraySlice_l159_157_1};
  assign _zz_when_ArraySlice_l159_157_2 = (_zz_when_ArraySlice_l159_157_3 - _zz_when_ArraySlice_l159_157_4);
  assign _zz_when_ArraySlice_l159_157_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_157_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_157_5);
  assign _zz_when_ArraySlice_l159_157_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_157_5 = {1'd0, _zz_when_ArraySlice_l159_157_6};
  assign _zz__zz_realValue_0_157 = {1'd0, wReg};
  assign _zz__zz_realValue_0_157_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_157_1 = (_zz_realValue_0_157_2 + _zz_realValue_0_157_3);
  assign _zz_realValue_0_157_2 = {1'd0, wReg};
  assign _zz_realValue_0_157_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_157_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_157 = {2'd0, _zz_when_ArraySlice_l166_157_1};
  assign _zz_when_ArraySlice_l166_157_2 = (_zz_when_ArraySlice_l166_157_3 + _zz_when_ArraySlice_l166_157_7);
  assign _zz_when_ArraySlice_l166_157_3 = (realValue_0_157 - _zz_when_ArraySlice_l166_157_4);
  assign _zz_when_ArraySlice_l166_157_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_157_5);
  assign _zz_when_ArraySlice_l166_157_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_157_5 = {1'd0, _zz_when_ArraySlice_l166_157_6};
  assign _zz_when_ArraySlice_l166_157_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_158 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_158_1);
  assign _zz_when_ArraySlice_l158_158_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_158_1 = {1'd0, _zz_when_ArraySlice_l158_158_2};
  assign _zz_when_ArraySlice_l158_158_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_158_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_158 = {2'd0, _zz_when_ArraySlice_l159_158_1};
  assign _zz_when_ArraySlice_l159_158_2 = (_zz_when_ArraySlice_l159_158_3 - _zz_when_ArraySlice_l159_158_4);
  assign _zz_when_ArraySlice_l159_158_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_158_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_158_5);
  assign _zz_when_ArraySlice_l159_158_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_158_5 = {1'd0, _zz_when_ArraySlice_l159_158_6};
  assign _zz__zz_realValue_0_158 = {1'd0, wReg};
  assign _zz__zz_realValue_0_158_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_158_1 = (_zz_realValue_0_158_2 + _zz_realValue_0_158_3);
  assign _zz_realValue_0_158_2 = {1'd0, wReg};
  assign _zz_realValue_0_158_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_158_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_158 = {2'd0, _zz_when_ArraySlice_l166_158_1};
  assign _zz_when_ArraySlice_l166_158_2 = (_zz_when_ArraySlice_l166_158_3 + _zz_when_ArraySlice_l166_158_7);
  assign _zz_when_ArraySlice_l166_158_3 = (realValue_0_158 - _zz_when_ArraySlice_l166_158_4);
  assign _zz_when_ArraySlice_l166_158_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_158_5);
  assign _zz_when_ArraySlice_l166_158_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_158_5 = {1'd0, _zz_when_ArraySlice_l166_158_6};
  assign _zz_when_ArraySlice_l166_158_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_159 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_159_1);
  assign _zz_when_ArraySlice_l158_159_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_159_1 = {1'd0, _zz_when_ArraySlice_l158_159_2};
  assign _zz_when_ArraySlice_l158_159_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_159_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_159 = {3'd0, _zz_when_ArraySlice_l159_159_1};
  assign _zz_when_ArraySlice_l159_159_2 = (_zz_when_ArraySlice_l159_159_3 - _zz_when_ArraySlice_l159_159_4);
  assign _zz_when_ArraySlice_l159_159_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_159_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_159_5);
  assign _zz_when_ArraySlice_l159_159_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_159_5 = {1'd0, _zz_when_ArraySlice_l159_159_6};
  assign _zz__zz_realValue_0_159 = {1'd0, wReg};
  assign _zz__zz_realValue_0_159_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_159_1 = (_zz_realValue_0_159_2 + _zz_realValue_0_159_3);
  assign _zz_realValue_0_159_2 = {1'd0, wReg};
  assign _zz_realValue_0_159_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_159_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_159 = {3'd0, _zz_when_ArraySlice_l166_159_1};
  assign _zz_when_ArraySlice_l166_159_2 = (_zz_when_ArraySlice_l166_159_3 + _zz_when_ArraySlice_l166_159_7);
  assign _zz_when_ArraySlice_l166_159_3 = (realValue_0_159 - _zz_when_ArraySlice_l166_159_4);
  assign _zz_when_ArraySlice_l166_159_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_159_5);
  assign _zz_when_ArraySlice_l166_159_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_159_5 = {1'd0, _zz_when_ArraySlice_l166_159_6};
  assign _zz_when_ArraySlice_l166_159_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_6_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_6_2 = (_zz_when_ArraySlice_l403_6_3 + _zz_when_ArraySlice_l403_6_7);
  assign _zz_when_ArraySlice_l403_6_3 = (_zz_when_ArraySlice_l403_6_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_6_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l403_6_5);
  assign _zz_when_ArraySlice_l403_6_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_6_5 = {1'd0, _zz_when_ArraySlice_l403_6_6};
  assign _zz_when_ArraySlice_l403_6_8 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l403_6_7 = {1'd0, _zz_when_ArraySlice_l403_6_8};
  assign _zz_when_ArraySlice_l406_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_6_1 = (_zz_when_ArraySlice_l406_6_2 + 8'h01);
  assign _zz_when_ArraySlice_l406_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l406_6_3);
  assign _zz_when_ArraySlice_l406_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_6_3 = {1'd0, _zz_when_ArraySlice_l406_6_4};
  assign _zz_selectReadFifo_6_6 = (selectReadFifo_6 + _zz_selectReadFifo_6_7);
  assign _zz_selectReadFifo_6_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_7 = {1'd0, _zz_selectReadFifo_6_8};
  assign _zz_when_ArraySlice_l413_6 = (_zz_when_ArraySlice_l413_6_1 % aReg);
  assign _zz_when_ArraySlice_l413_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l417_6_3);
  assign _zz_when_ArraySlice_l417_6_1 = _zz_when_ArraySlice_l417_6_2[6:0];
  assign _zz_when_ArraySlice_l417_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l417_6_3 = {1'd0, _zz_when_ArraySlice_l417_6_4};
  assign _zz_when_ArraySlice_l418_6_1 = (_zz_when_ArraySlice_l418_6_2 - _zz_when_ArraySlice_l418_6_3);
  assign _zz_when_ArraySlice_l418_6 = {5'd0, _zz_when_ArraySlice_l418_6_1};
  assign _zz_when_ArraySlice_l418_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l418_6_3 = {7'd0, _zz_when_ArraySlice_l418_6_4};
  assign _zz__zz_realValue1_0_19 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_19_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_19_1 = (_zz_realValue1_0_19_2 + _zz_realValue1_0_19_3);
  assign _zz_realValue1_0_19_2 = {1'd0, hReg};
  assign _zz_realValue1_0_19_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l420_6 = {1'd0, _zz_when_ArraySlice_l420_6_1};
  assign _zz_when_ArraySlice_l420_6_2 = (realValue1_0_19 / aReg);
  assign _zz_selectReadFifo_6_9 = (selectReadFifo_6 - _zz_selectReadFifo_6_10);
  assign _zz_selectReadFifo_6_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_160 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_160_1);
  assign _zz_when_ArraySlice_l158_160_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_160_1 = {4'd0, _zz_when_ArraySlice_l158_160_2};
  assign _zz_when_ArraySlice_l158_160_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_160 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_160_1 = (_zz_when_ArraySlice_l159_160_2 - _zz_when_ArraySlice_l159_160_3);
  assign _zz_when_ArraySlice_l159_160_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_160_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_160_4);
  assign _zz_when_ArraySlice_l159_160_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_160_4 = {4'd0, _zz_when_ArraySlice_l159_160_5};
  assign _zz__zz_realValue_0_160 = {1'd0, wReg};
  assign _zz__zz_realValue_0_160_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_160_1 = (_zz_realValue_0_160_2 + _zz_realValue_0_160_3);
  assign _zz_realValue_0_160_2 = {1'd0, wReg};
  assign _zz_realValue_0_160_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_160 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_160_1 = (_zz_when_ArraySlice_l166_160_2 + _zz_when_ArraySlice_l166_160_6);
  assign _zz_when_ArraySlice_l166_160_2 = (realValue_0_160 - _zz_when_ArraySlice_l166_160_3);
  assign _zz_when_ArraySlice_l166_160_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_160_4);
  assign _zz_when_ArraySlice_l166_160_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_160_4 = {4'd0, _zz_when_ArraySlice_l166_160_5};
  assign _zz_when_ArraySlice_l166_160_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_161 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_161_1);
  assign _zz_when_ArraySlice_l158_161_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_161_1 = {3'd0, _zz_when_ArraySlice_l158_161_2};
  assign _zz_when_ArraySlice_l158_161_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_161_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_161 = {1'd0, _zz_when_ArraySlice_l159_161_1};
  assign _zz_when_ArraySlice_l159_161_2 = (_zz_when_ArraySlice_l159_161_3 - _zz_when_ArraySlice_l159_161_4);
  assign _zz_when_ArraySlice_l159_161_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_161_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_161_5);
  assign _zz_when_ArraySlice_l159_161_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_161_5 = {3'd0, _zz_when_ArraySlice_l159_161_6};
  assign _zz__zz_realValue_0_161 = {1'd0, wReg};
  assign _zz__zz_realValue_0_161_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_161_1 = (_zz_realValue_0_161_2 + _zz_realValue_0_161_3);
  assign _zz_realValue_0_161_2 = {1'd0, wReg};
  assign _zz_realValue_0_161_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_161_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_161 = {1'd0, _zz_when_ArraySlice_l166_161_1};
  assign _zz_when_ArraySlice_l166_161_2 = (_zz_when_ArraySlice_l166_161_3 + _zz_when_ArraySlice_l166_161_7);
  assign _zz_when_ArraySlice_l166_161_3 = (realValue_0_161 - _zz_when_ArraySlice_l166_161_4);
  assign _zz_when_ArraySlice_l166_161_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_161_5);
  assign _zz_when_ArraySlice_l166_161_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_161_5 = {3'd0, _zz_when_ArraySlice_l166_161_6};
  assign _zz_when_ArraySlice_l166_161_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_162 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_162_1);
  assign _zz_when_ArraySlice_l158_162_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_162_1 = {2'd0, _zz_when_ArraySlice_l158_162_2};
  assign _zz_when_ArraySlice_l158_162_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_162_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_162 = {1'd0, _zz_when_ArraySlice_l159_162_1};
  assign _zz_when_ArraySlice_l159_162_2 = (_zz_when_ArraySlice_l159_162_3 - _zz_when_ArraySlice_l159_162_4);
  assign _zz_when_ArraySlice_l159_162_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_162_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_162_5);
  assign _zz_when_ArraySlice_l159_162_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_162_5 = {2'd0, _zz_when_ArraySlice_l159_162_6};
  assign _zz__zz_realValue_0_162 = {1'd0, wReg};
  assign _zz__zz_realValue_0_162_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_162_1 = (_zz_realValue_0_162_2 + _zz_realValue_0_162_3);
  assign _zz_realValue_0_162_2 = {1'd0, wReg};
  assign _zz_realValue_0_162_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_162_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_162 = {1'd0, _zz_when_ArraySlice_l166_162_1};
  assign _zz_when_ArraySlice_l166_162_2 = (_zz_when_ArraySlice_l166_162_3 + _zz_when_ArraySlice_l166_162_7);
  assign _zz_when_ArraySlice_l166_162_3 = (realValue_0_162 - _zz_when_ArraySlice_l166_162_4);
  assign _zz_when_ArraySlice_l166_162_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_162_5);
  assign _zz_when_ArraySlice_l166_162_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_162_5 = {2'd0, _zz_when_ArraySlice_l166_162_6};
  assign _zz_when_ArraySlice_l166_162_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_163 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_163_1);
  assign _zz_when_ArraySlice_l158_163_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_163_1 = {2'd0, _zz_when_ArraySlice_l158_163_2};
  assign _zz_when_ArraySlice_l158_163_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_163_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_163 = {1'd0, _zz_when_ArraySlice_l159_163_1};
  assign _zz_when_ArraySlice_l159_163_2 = (_zz_when_ArraySlice_l159_163_3 - _zz_when_ArraySlice_l159_163_4);
  assign _zz_when_ArraySlice_l159_163_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_163_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_163_5);
  assign _zz_when_ArraySlice_l159_163_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_163_5 = {2'd0, _zz_when_ArraySlice_l159_163_6};
  assign _zz__zz_realValue_0_163 = {1'd0, wReg};
  assign _zz__zz_realValue_0_163_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_163_1 = (_zz_realValue_0_163_2 + _zz_realValue_0_163_3);
  assign _zz_realValue_0_163_2 = {1'd0, wReg};
  assign _zz_realValue_0_163_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_163_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_163 = {1'd0, _zz_when_ArraySlice_l166_163_1};
  assign _zz_when_ArraySlice_l166_163_2 = (_zz_when_ArraySlice_l166_163_3 + _zz_when_ArraySlice_l166_163_7);
  assign _zz_when_ArraySlice_l166_163_3 = (realValue_0_163 - _zz_when_ArraySlice_l166_163_4);
  assign _zz_when_ArraySlice_l166_163_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_163_5);
  assign _zz_when_ArraySlice_l166_163_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_163_5 = {2'd0, _zz_when_ArraySlice_l166_163_6};
  assign _zz_when_ArraySlice_l166_163_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_164 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_164_1);
  assign _zz_when_ArraySlice_l158_164_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_164_1 = {1'd0, _zz_when_ArraySlice_l158_164_2};
  assign _zz_when_ArraySlice_l158_164_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_164_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_164 = {1'd0, _zz_when_ArraySlice_l159_164_1};
  assign _zz_when_ArraySlice_l159_164_2 = (_zz_when_ArraySlice_l159_164_3 - _zz_when_ArraySlice_l159_164_4);
  assign _zz_when_ArraySlice_l159_164_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_164_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_164_5);
  assign _zz_when_ArraySlice_l159_164_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_164_5 = {1'd0, _zz_when_ArraySlice_l159_164_6};
  assign _zz__zz_realValue_0_164 = {1'd0, wReg};
  assign _zz__zz_realValue_0_164_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_164_1 = (_zz_realValue_0_164_2 + _zz_realValue_0_164_3);
  assign _zz_realValue_0_164_2 = {1'd0, wReg};
  assign _zz_realValue_0_164_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_164_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_164 = {1'd0, _zz_when_ArraySlice_l166_164_1};
  assign _zz_when_ArraySlice_l166_164_2 = (_zz_when_ArraySlice_l166_164_3 + _zz_when_ArraySlice_l166_164_7);
  assign _zz_when_ArraySlice_l166_164_3 = (realValue_0_164 - _zz_when_ArraySlice_l166_164_4);
  assign _zz_when_ArraySlice_l166_164_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_164_5);
  assign _zz_when_ArraySlice_l166_164_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_164_5 = {1'd0, _zz_when_ArraySlice_l166_164_6};
  assign _zz_when_ArraySlice_l166_164_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_165 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_165_1);
  assign _zz_when_ArraySlice_l158_165_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_165_1 = {1'd0, _zz_when_ArraySlice_l158_165_2};
  assign _zz_when_ArraySlice_l158_165_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_165_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_165 = {2'd0, _zz_when_ArraySlice_l159_165_1};
  assign _zz_when_ArraySlice_l159_165_2 = (_zz_when_ArraySlice_l159_165_3 - _zz_when_ArraySlice_l159_165_4);
  assign _zz_when_ArraySlice_l159_165_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_165_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_165_5);
  assign _zz_when_ArraySlice_l159_165_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_165_5 = {1'd0, _zz_when_ArraySlice_l159_165_6};
  assign _zz__zz_realValue_0_165 = {1'd0, wReg};
  assign _zz__zz_realValue_0_165_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_165_1 = (_zz_realValue_0_165_2 + _zz_realValue_0_165_3);
  assign _zz_realValue_0_165_2 = {1'd0, wReg};
  assign _zz_realValue_0_165_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_165_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_165 = {2'd0, _zz_when_ArraySlice_l166_165_1};
  assign _zz_when_ArraySlice_l166_165_2 = (_zz_when_ArraySlice_l166_165_3 + _zz_when_ArraySlice_l166_165_7);
  assign _zz_when_ArraySlice_l166_165_3 = (realValue_0_165 - _zz_when_ArraySlice_l166_165_4);
  assign _zz_when_ArraySlice_l166_165_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_165_5);
  assign _zz_when_ArraySlice_l166_165_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_165_5 = {1'd0, _zz_when_ArraySlice_l166_165_6};
  assign _zz_when_ArraySlice_l166_165_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_166 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_166_1);
  assign _zz_when_ArraySlice_l158_166_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_166_1 = {1'd0, _zz_when_ArraySlice_l158_166_2};
  assign _zz_when_ArraySlice_l158_166_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_166_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_166 = {2'd0, _zz_when_ArraySlice_l159_166_1};
  assign _zz_when_ArraySlice_l159_166_2 = (_zz_when_ArraySlice_l159_166_3 - _zz_when_ArraySlice_l159_166_4);
  assign _zz_when_ArraySlice_l159_166_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_166_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_166_5);
  assign _zz_when_ArraySlice_l159_166_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_166_5 = {1'd0, _zz_when_ArraySlice_l159_166_6};
  assign _zz__zz_realValue_0_166 = {1'd0, wReg};
  assign _zz__zz_realValue_0_166_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_166_1 = (_zz_realValue_0_166_2 + _zz_realValue_0_166_3);
  assign _zz_realValue_0_166_2 = {1'd0, wReg};
  assign _zz_realValue_0_166_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_166_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_166 = {2'd0, _zz_when_ArraySlice_l166_166_1};
  assign _zz_when_ArraySlice_l166_166_2 = (_zz_when_ArraySlice_l166_166_3 + _zz_when_ArraySlice_l166_166_7);
  assign _zz_when_ArraySlice_l166_166_3 = (realValue_0_166 - _zz_when_ArraySlice_l166_166_4);
  assign _zz_when_ArraySlice_l166_166_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_166_5);
  assign _zz_when_ArraySlice_l166_166_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_166_5 = {1'd0, _zz_when_ArraySlice_l166_166_6};
  assign _zz_when_ArraySlice_l166_166_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_167 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_167_1);
  assign _zz_when_ArraySlice_l158_167_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_167_1 = {1'd0, _zz_when_ArraySlice_l158_167_2};
  assign _zz_when_ArraySlice_l158_167_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_167_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_167 = {3'd0, _zz_when_ArraySlice_l159_167_1};
  assign _zz_when_ArraySlice_l159_167_2 = (_zz_when_ArraySlice_l159_167_3 - _zz_when_ArraySlice_l159_167_4);
  assign _zz_when_ArraySlice_l159_167_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_167_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_167_5);
  assign _zz_when_ArraySlice_l159_167_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_167_5 = {1'd0, _zz_when_ArraySlice_l159_167_6};
  assign _zz__zz_realValue_0_167 = {1'd0, wReg};
  assign _zz__zz_realValue_0_167_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_167_1 = (_zz_realValue_0_167_2 + _zz_realValue_0_167_3);
  assign _zz_realValue_0_167_2 = {1'd0, wReg};
  assign _zz_realValue_0_167_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_167_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_167 = {3'd0, _zz_when_ArraySlice_l166_167_1};
  assign _zz_when_ArraySlice_l166_167_2 = (_zz_when_ArraySlice_l166_167_3 + _zz_when_ArraySlice_l166_167_7);
  assign _zz_when_ArraySlice_l166_167_3 = (realValue_0_167 - _zz_when_ArraySlice_l166_167_4);
  assign _zz_when_ArraySlice_l166_167_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_167_5);
  assign _zz_when_ArraySlice_l166_167_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_167_5 = {1'd0, _zz_when_ArraySlice_l166_167_6};
  assign _zz_when_ArraySlice_l166_167_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_6_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_6_2 = (_zz_when_ArraySlice_l428_6_3 + _zz_when_ArraySlice_l428_6_7);
  assign _zz_when_ArraySlice_l428_6_3 = (_zz_when_ArraySlice_l428_6_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_6_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l428_6_5);
  assign _zz_when_ArraySlice_l428_6_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_6_5 = {1'd0, _zz_when_ArraySlice_l428_6_6};
  assign _zz_when_ArraySlice_l428_6_8 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l428_6_7 = {1'd0, _zz_when_ArraySlice_l428_6_8};
  assign _zz_when_ArraySlice_l431_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_6_1 = (_zz_when_ArraySlice_l431_6_2 + 8'h01);
  assign _zz_when_ArraySlice_l431_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l431_6_3);
  assign _zz_when_ArraySlice_l431_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_6_3 = {1'd0, _zz_when_ArraySlice_l431_6_4};
  assign _zz_selectReadFifo_6_11 = (selectReadFifo_6 + _zz_selectReadFifo_6_12);
  assign _zz_selectReadFifo_6_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_12 = {1'd0, _zz_selectReadFifo_6_13};
  assign _zz_when_ArraySlice_l438_6 = (_zz_when_ArraySlice_l438_6_1 % aReg);
  assign _zz_when_ArraySlice_l438_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_6_1 = (_zz_when_ArraySlice_l449_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l449_6 = {5'd0, _zz_when_ArraySlice_l449_6_1};
  assign _zz_when_ArraySlice_l449_6_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_20 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_20_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_20_1 = (_zz_realValue1_0_20_2 + _zz_realValue1_0_20_3);
  assign _zz_realValue1_0_20_2 = {1'd0, hReg};
  assign _zz_realValue1_0_20_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l450_6 = {1'd0, _zz_when_ArraySlice_l450_6_1};
  assign _zz_when_ArraySlice_l450_6_2 = (realValue1_0_20 / aReg);
  assign _zz_selectReadFifo_6_14 = (selectReadFifo_6 - _zz_selectReadFifo_6_15);
  assign _zz_selectReadFifo_6_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_168 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_168_1);
  assign _zz_when_ArraySlice_l158_168_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_168_1 = {4'd0, _zz_when_ArraySlice_l158_168_2};
  assign _zz_when_ArraySlice_l158_168_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_168 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_168_1 = (_zz_when_ArraySlice_l159_168_2 - _zz_when_ArraySlice_l159_168_3);
  assign _zz_when_ArraySlice_l159_168_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_168_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_168_4);
  assign _zz_when_ArraySlice_l159_168_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_168_4 = {4'd0, _zz_when_ArraySlice_l159_168_5};
  assign _zz__zz_realValue_0_168 = {1'd0, wReg};
  assign _zz__zz_realValue_0_168_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_168_1 = (_zz_realValue_0_168_2 + _zz_realValue_0_168_3);
  assign _zz_realValue_0_168_2 = {1'd0, wReg};
  assign _zz_realValue_0_168_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_168 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_168_1 = (_zz_when_ArraySlice_l166_168_2 + _zz_when_ArraySlice_l166_168_6);
  assign _zz_when_ArraySlice_l166_168_2 = (realValue_0_168 - _zz_when_ArraySlice_l166_168_3);
  assign _zz_when_ArraySlice_l166_168_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_168_4);
  assign _zz_when_ArraySlice_l166_168_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_168_4 = {4'd0, _zz_when_ArraySlice_l166_168_5};
  assign _zz_when_ArraySlice_l166_168_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_169 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_169_1);
  assign _zz_when_ArraySlice_l158_169_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_169_1 = {3'd0, _zz_when_ArraySlice_l158_169_2};
  assign _zz_when_ArraySlice_l158_169_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_169_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_169 = {1'd0, _zz_when_ArraySlice_l159_169_1};
  assign _zz_when_ArraySlice_l159_169_2 = (_zz_when_ArraySlice_l159_169_3 - _zz_when_ArraySlice_l159_169_4);
  assign _zz_when_ArraySlice_l159_169_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_169_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_169_5);
  assign _zz_when_ArraySlice_l159_169_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_169_5 = {3'd0, _zz_when_ArraySlice_l159_169_6};
  assign _zz__zz_realValue_0_169 = {1'd0, wReg};
  assign _zz__zz_realValue_0_169_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_169_1 = (_zz_realValue_0_169_2 + _zz_realValue_0_169_3);
  assign _zz_realValue_0_169_2 = {1'd0, wReg};
  assign _zz_realValue_0_169_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_169_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_169 = {1'd0, _zz_when_ArraySlice_l166_169_1};
  assign _zz_when_ArraySlice_l166_169_2 = (_zz_when_ArraySlice_l166_169_3 + _zz_when_ArraySlice_l166_169_7);
  assign _zz_when_ArraySlice_l166_169_3 = (realValue_0_169 - _zz_when_ArraySlice_l166_169_4);
  assign _zz_when_ArraySlice_l166_169_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_169_5);
  assign _zz_when_ArraySlice_l166_169_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_169_5 = {3'd0, _zz_when_ArraySlice_l166_169_6};
  assign _zz_when_ArraySlice_l166_169_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_170 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_170_1);
  assign _zz_when_ArraySlice_l158_170_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_170_1 = {2'd0, _zz_when_ArraySlice_l158_170_2};
  assign _zz_when_ArraySlice_l158_170_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_170_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_170 = {1'd0, _zz_when_ArraySlice_l159_170_1};
  assign _zz_when_ArraySlice_l159_170_2 = (_zz_when_ArraySlice_l159_170_3 - _zz_when_ArraySlice_l159_170_4);
  assign _zz_when_ArraySlice_l159_170_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_170_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_170_5);
  assign _zz_when_ArraySlice_l159_170_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_170_5 = {2'd0, _zz_when_ArraySlice_l159_170_6};
  assign _zz__zz_realValue_0_170 = {1'd0, wReg};
  assign _zz__zz_realValue_0_170_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_170_1 = (_zz_realValue_0_170_2 + _zz_realValue_0_170_3);
  assign _zz_realValue_0_170_2 = {1'd0, wReg};
  assign _zz_realValue_0_170_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_170_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_170 = {1'd0, _zz_when_ArraySlice_l166_170_1};
  assign _zz_when_ArraySlice_l166_170_2 = (_zz_when_ArraySlice_l166_170_3 + _zz_when_ArraySlice_l166_170_7);
  assign _zz_when_ArraySlice_l166_170_3 = (realValue_0_170 - _zz_when_ArraySlice_l166_170_4);
  assign _zz_when_ArraySlice_l166_170_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_170_5);
  assign _zz_when_ArraySlice_l166_170_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_170_5 = {2'd0, _zz_when_ArraySlice_l166_170_6};
  assign _zz_when_ArraySlice_l166_170_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_171 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_171_1);
  assign _zz_when_ArraySlice_l158_171_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_171_1 = {2'd0, _zz_when_ArraySlice_l158_171_2};
  assign _zz_when_ArraySlice_l158_171_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_171_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_171 = {1'd0, _zz_when_ArraySlice_l159_171_1};
  assign _zz_when_ArraySlice_l159_171_2 = (_zz_when_ArraySlice_l159_171_3 - _zz_when_ArraySlice_l159_171_4);
  assign _zz_when_ArraySlice_l159_171_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_171_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_171_5);
  assign _zz_when_ArraySlice_l159_171_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_171_5 = {2'd0, _zz_when_ArraySlice_l159_171_6};
  assign _zz__zz_realValue_0_171 = {1'd0, wReg};
  assign _zz__zz_realValue_0_171_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_171_1 = (_zz_realValue_0_171_2 + _zz_realValue_0_171_3);
  assign _zz_realValue_0_171_2 = {1'd0, wReg};
  assign _zz_realValue_0_171_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_171_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_171 = {1'd0, _zz_when_ArraySlice_l166_171_1};
  assign _zz_when_ArraySlice_l166_171_2 = (_zz_when_ArraySlice_l166_171_3 + _zz_when_ArraySlice_l166_171_7);
  assign _zz_when_ArraySlice_l166_171_3 = (realValue_0_171 - _zz_when_ArraySlice_l166_171_4);
  assign _zz_when_ArraySlice_l166_171_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_171_5);
  assign _zz_when_ArraySlice_l166_171_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_171_5 = {2'd0, _zz_when_ArraySlice_l166_171_6};
  assign _zz_when_ArraySlice_l166_171_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_172 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_172_1);
  assign _zz_when_ArraySlice_l158_172_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_172_1 = {1'd0, _zz_when_ArraySlice_l158_172_2};
  assign _zz_when_ArraySlice_l158_172_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_172_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_172 = {1'd0, _zz_when_ArraySlice_l159_172_1};
  assign _zz_when_ArraySlice_l159_172_2 = (_zz_when_ArraySlice_l159_172_3 - _zz_when_ArraySlice_l159_172_4);
  assign _zz_when_ArraySlice_l159_172_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_172_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_172_5);
  assign _zz_when_ArraySlice_l159_172_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_172_5 = {1'd0, _zz_when_ArraySlice_l159_172_6};
  assign _zz__zz_realValue_0_172 = {1'd0, wReg};
  assign _zz__zz_realValue_0_172_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_172_1 = (_zz_realValue_0_172_2 + _zz_realValue_0_172_3);
  assign _zz_realValue_0_172_2 = {1'd0, wReg};
  assign _zz_realValue_0_172_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_172_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_172 = {1'd0, _zz_when_ArraySlice_l166_172_1};
  assign _zz_when_ArraySlice_l166_172_2 = (_zz_when_ArraySlice_l166_172_3 + _zz_when_ArraySlice_l166_172_7);
  assign _zz_when_ArraySlice_l166_172_3 = (realValue_0_172 - _zz_when_ArraySlice_l166_172_4);
  assign _zz_when_ArraySlice_l166_172_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_172_5);
  assign _zz_when_ArraySlice_l166_172_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_172_5 = {1'd0, _zz_when_ArraySlice_l166_172_6};
  assign _zz_when_ArraySlice_l166_172_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_173 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_173_1);
  assign _zz_when_ArraySlice_l158_173_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_173_1 = {1'd0, _zz_when_ArraySlice_l158_173_2};
  assign _zz_when_ArraySlice_l158_173_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_173_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_173 = {2'd0, _zz_when_ArraySlice_l159_173_1};
  assign _zz_when_ArraySlice_l159_173_2 = (_zz_when_ArraySlice_l159_173_3 - _zz_when_ArraySlice_l159_173_4);
  assign _zz_when_ArraySlice_l159_173_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_173_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_173_5);
  assign _zz_when_ArraySlice_l159_173_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_173_5 = {1'd0, _zz_when_ArraySlice_l159_173_6};
  assign _zz__zz_realValue_0_173 = {1'd0, wReg};
  assign _zz__zz_realValue_0_173_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_173_1 = (_zz_realValue_0_173_2 + _zz_realValue_0_173_3);
  assign _zz_realValue_0_173_2 = {1'd0, wReg};
  assign _zz_realValue_0_173_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_173_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_173 = {2'd0, _zz_when_ArraySlice_l166_173_1};
  assign _zz_when_ArraySlice_l166_173_2 = (_zz_when_ArraySlice_l166_173_3 + _zz_when_ArraySlice_l166_173_7);
  assign _zz_when_ArraySlice_l166_173_3 = (realValue_0_173 - _zz_when_ArraySlice_l166_173_4);
  assign _zz_when_ArraySlice_l166_173_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_173_5);
  assign _zz_when_ArraySlice_l166_173_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_173_5 = {1'd0, _zz_when_ArraySlice_l166_173_6};
  assign _zz_when_ArraySlice_l166_173_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_174 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_174_1);
  assign _zz_when_ArraySlice_l158_174_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_174_1 = {1'd0, _zz_when_ArraySlice_l158_174_2};
  assign _zz_when_ArraySlice_l158_174_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_174_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_174 = {2'd0, _zz_when_ArraySlice_l159_174_1};
  assign _zz_when_ArraySlice_l159_174_2 = (_zz_when_ArraySlice_l159_174_3 - _zz_when_ArraySlice_l159_174_4);
  assign _zz_when_ArraySlice_l159_174_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_174_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_174_5);
  assign _zz_when_ArraySlice_l159_174_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_174_5 = {1'd0, _zz_when_ArraySlice_l159_174_6};
  assign _zz__zz_realValue_0_174 = {1'd0, wReg};
  assign _zz__zz_realValue_0_174_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_174_1 = (_zz_realValue_0_174_2 + _zz_realValue_0_174_3);
  assign _zz_realValue_0_174_2 = {1'd0, wReg};
  assign _zz_realValue_0_174_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_174_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_174 = {2'd0, _zz_when_ArraySlice_l166_174_1};
  assign _zz_when_ArraySlice_l166_174_2 = (_zz_when_ArraySlice_l166_174_3 + _zz_when_ArraySlice_l166_174_7);
  assign _zz_when_ArraySlice_l166_174_3 = (realValue_0_174 - _zz_when_ArraySlice_l166_174_4);
  assign _zz_when_ArraySlice_l166_174_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_174_5);
  assign _zz_when_ArraySlice_l166_174_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_174_5 = {1'd0, _zz_when_ArraySlice_l166_174_6};
  assign _zz_when_ArraySlice_l166_174_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_175 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_175_1);
  assign _zz_when_ArraySlice_l158_175_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_175_1 = {1'd0, _zz_when_ArraySlice_l158_175_2};
  assign _zz_when_ArraySlice_l158_175_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_175_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_175 = {3'd0, _zz_when_ArraySlice_l159_175_1};
  assign _zz_when_ArraySlice_l159_175_2 = (_zz_when_ArraySlice_l159_175_3 - _zz_when_ArraySlice_l159_175_4);
  assign _zz_when_ArraySlice_l159_175_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_175_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_175_5);
  assign _zz_when_ArraySlice_l159_175_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_175_5 = {1'd0, _zz_when_ArraySlice_l159_175_6};
  assign _zz__zz_realValue_0_175 = {1'd0, wReg};
  assign _zz__zz_realValue_0_175_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_175_1 = (_zz_realValue_0_175_2 + _zz_realValue_0_175_3);
  assign _zz_realValue_0_175_2 = {1'd0, wReg};
  assign _zz_realValue_0_175_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_175_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_175 = {3'd0, _zz_when_ArraySlice_l166_175_1};
  assign _zz_when_ArraySlice_l166_175_2 = (_zz_when_ArraySlice_l166_175_3 + _zz_when_ArraySlice_l166_175_7);
  assign _zz_when_ArraySlice_l166_175_3 = (realValue_0_175 - _zz_when_ArraySlice_l166_175_4);
  assign _zz_when_ArraySlice_l166_175_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_175_5);
  assign _zz_when_ArraySlice_l166_175_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_175_5 = {1'd0, _zz_when_ArraySlice_l166_175_6};
  assign _zz_when_ArraySlice_l166_175_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_6 = (_zz_when_ArraySlice_l461_6_1 % aReg);
  assign _zz_when_ArraySlice_l461_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l447_6_2);
  assign _zz_when_ArraySlice_l447_6_3 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l447_6_2 = {1'd0, _zz_when_ArraySlice_l447_6_3};
  assign _zz_when_ArraySlice_l468_6_1 = (_zz_when_ArraySlice_l468_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l468_6 = {5'd0, _zz_when_ArraySlice_l468_6_1};
  assign _zz_when_ArraySlice_l468_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l376_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l376_7_1);
  assign _zz_when_ArraySlice_l376_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l376_7_1 = {1'd0, _zz_when_ArraySlice_l376_7_2};
  assign _zz_when_ArraySlice_l376_7_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l377_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l377_7_3);
  assign _zz_when_ArraySlice_l377_7_1 = _zz_when_ArraySlice_l377_7_2[6:0];
  assign _zz_when_ArraySlice_l377_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l377_7_3 = {1'd0, _zz_when_ArraySlice_l377_7_4};
  assign _zz__zz_outputStreamArrayData_7_valid_1 = (bReg * 3'b111);
  assign _zz__zz_outputStreamArrayData_7_valid = {1'd0, _zz__zz_outputStreamArrayData_7_valid_1};
  assign _zz__zz_10 = _zz_outputStreamArrayData_7_valid[6:0];
  assign _zz_outputStreamArrayData_7_valid_3 = _zz_outputStreamArrayData_7_valid[6:0];
  assign _zz_outputStreamArrayData_7_payload_1 = _zz_outputStreamArrayData_7_valid[6:0];
  assign _zz_when_ArraySlice_l383_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l383_7_3);
  assign _zz_when_ArraySlice_l383_7_1 = _zz_when_ArraySlice_l383_7_2[6:0];
  assign _zz_when_ArraySlice_l383_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l383_7_3 = {1'd0, _zz_when_ArraySlice_l383_7_4};
  assign _zz_when_ArraySlice_l384_7_1 = (_zz_when_ArraySlice_l384_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l384_7 = {5'd0, _zz_when_ArraySlice_l384_7_1};
  assign _zz_when_ArraySlice_l384_7_2 = (bReg * aReg);
  assign _zz_selectReadFifo_7 = (selectReadFifo_7 - _zz_selectReadFifo_7_1);
  assign _zz_selectReadFifo_7_1 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l387_7 = (_zz_when_ArraySlice_l387_7_1 % aReg);
  assign _zz_when_ArraySlice_l387_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l392_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l392_7_3);
  assign _zz_when_ArraySlice_l392_7_1 = _zz_when_ArraySlice_l392_7_2[6:0];
  assign _zz_when_ArraySlice_l392_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l392_7_3 = {1'd0, _zz_when_ArraySlice_l392_7_4};
  assign _zz_when_ArraySlice_l393_7_1 = (_zz_when_ArraySlice_l393_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l393_7 = {5'd0, _zz_when_ArraySlice_l393_7_1};
  assign _zz_when_ArraySlice_l393_7_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_21 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_21_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_21_1 = (_zz_realValue1_0_21_2 + _zz_realValue1_0_21_3);
  assign _zz_realValue1_0_21_2 = {1'd0, hReg};
  assign _zz_realValue1_0_21_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l395_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l395_7 = {1'd0, _zz_when_ArraySlice_l395_7_1};
  assign _zz_when_ArraySlice_l395_7_2 = (realValue1_0_21 / aReg);
  assign _zz_selectReadFifo_7_2 = (selectReadFifo_7 - _zz_selectReadFifo_7_3);
  assign _zz_selectReadFifo_7_3 = {4'd0, bReg};
  assign _zz_selectReadFifo_7_5 = 1'b1;
  assign _zz_selectReadFifo_7_4 = {7'd0, _zz_selectReadFifo_7_5};
  assign _zz_when_ArraySlice_l158_176 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_176_1);
  assign _zz_when_ArraySlice_l158_176_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_176_1 = {4'd0, _zz_when_ArraySlice_l158_176_2};
  assign _zz_when_ArraySlice_l158_176_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_176 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_176_1 = (_zz_when_ArraySlice_l159_176_2 - _zz_when_ArraySlice_l159_176_3);
  assign _zz_when_ArraySlice_l159_176_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_176_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_176_4);
  assign _zz_when_ArraySlice_l159_176_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_176_4 = {4'd0, _zz_when_ArraySlice_l159_176_5};
  assign _zz__zz_realValue_0_176 = {1'd0, wReg};
  assign _zz__zz_realValue_0_176_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_176_1 = (_zz_realValue_0_176_2 + _zz_realValue_0_176_3);
  assign _zz_realValue_0_176_2 = {1'd0, wReg};
  assign _zz_realValue_0_176_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_176 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_176_1 = (_zz_when_ArraySlice_l166_176_2 + _zz_when_ArraySlice_l166_176_6);
  assign _zz_when_ArraySlice_l166_176_2 = (realValue_0_176 - _zz_when_ArraySlice_l166_176_3);
  assign _zz_when_ArraySlice_l166_176_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_176_4);
  assign _zz_when_ArraySlice_l166_176_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_176_4 = {4'd0, _zz_when_ArraySlice_l166_176_5};
  assign _zz_when_ArraySlice_l166_176_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_177 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_177_1);
  assign _zz_when_ArraySlice_l158_177_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_177_1 = {3'd0, _zz_when_ArraySlice_l158_177_2};
  assign _zz_when_ArraySlice_l158_177_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_177_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_177 = {1'd0, _zz_when_ArraySlice_l159_177_1};
  assign _zz_when_ArraySlice_l159_177_2 = (_zz_when_ArraySlice_l159_177_3 - _zz_when_ArraySlice_l159_177_4);
  assign _zz_when_ArraySlice_l159_177_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_177_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_177_5);
  assign _zz_when_ArraySlice_l159_177_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_177_5 = {3'd0, _zz_when_ArraySlice_l159_177_6};
  assign _zz__zz_realValue_0_177 = {1'd0, wReg};
  assign _zz__zz_realValue_0_177_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_177_1 = (_zz_realValue_0_177_2 + _zz_realValue_0_177_3);
  assign _zz_realValue_0_177_2 = {1'd0, wReg};
  assign _zz_realValue_0_177_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_177_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_177 = {1'd0, _zz_when_ArraySlice_l166_177_1};
  assign _zz_when_ArraySlice_l166_177_2 = (_zz_when_ArraySlice_l166_177_3 + _zz_when_ArraySlice_l166_177_7);
  assign _zz_when_ArraySlice_l166_177_3 = (realValue_0_177 - _zz_when_ArraySlice_l166_177_4);
  assign _zz_when_ArraySlice_l166_177_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_177_5);
  assign _zz_when_ArraySlice_l166_177_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_177_5 = {3'd0, _zz_when_ArraySlice_l166_177_6};
  assign _zz_when_ArraySlice_l166_177_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_178 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_178_1);
  assign _zz_when_ArraySlice_l158_178_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_178_1 = {2'd0, _zz_when_ArraySlice_l158_178_2};
  assign _zz_when_ArraySlice_l158_178_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_178_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_178 = {1'd0, _zz_when_ArraySlice_l159_178_1};
  assign _zz_when_ArraySlice_l159_178_2 = (_zz_when_ArraySlice_l159_178_3 - _zz_when_ArraySlice_l159_178_4);
  assign _zz_when_ArraySlice_l159_178_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_178_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_178_5);
  assign _zz_when_ArraySlice_l159_178_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_178_5 = {2'd0, _zz_when_ArraySlice_l159_178_6};
  assign _zz__zz_realValue_0_178 = {1'd0, wReg};
  assign _zz__zz_realValue_0_178_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_178_1 = (_zz_realValue_0_178_2 + _zz_realValue_0_178_3);
  assign _zz_realValue_0_178_2 = {1'd0, wReg};
  assign _zz_realValue_0_178_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_178_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_178 = {1'd0, _zz_when_ArraySlice_l166_178_1};
  assign _zz_when_ArraySlice_l166_178_2 = (_zz_when_ArraySlice_l166_178_3 + _zz_when_ArraySlice_l166_178_7);
  assign _zz_when_ArraySlice_l166_178_3 = (realValue_0_178 - _zz_when_ArraySlice_l166_178_4);
  assign _zz_when_ArraySlice_l166_178_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_178_5);
  assign _zz_when_ArraySlice_l166_178_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_178_5 = {2'd0, _zz_when_ArraySlice_l166_178_6};
  assign _zz_when_ArraySlice_l166_178_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_179 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_179_1);
  assign _zz_when_ArraySlice_l158_179_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_179_1 = {2'd0, _zz_when_ArraySlice_l158_179_2};
  assign _zz_when_ArraySlice_l158_179_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_179_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_179 = {1'd0, _zz_when_ArraySlice_l159_179_1};
  assign _zz_when_ArraySlice_l159_179_2 = (_zz_when_ArraySlice_l159_179_3 - _zz_when_ArraySlice_l159_179_4);
  assign _zz_when_ArraySlice_l159_179_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_179_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_179_5);
  assign _zz_when_ArraySlice_l159_179_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_179_5 = {2'd0, _zz_when_ArraySlice_l159_179_6};
  assign _zz__zz_realValue_0_179 = {1'd0, wReg};
  assign _zz__zz_realValue_0_179_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_179_1 = (_zz_realValue_0_179_2 + _zz_realValue_0_179_3);
  assign _zz_realValue_0_179_2 = {1'd0, wReg};
  assign _zz_realValue_0_179_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_179_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_179 = {1'd0, _zz_when_ArraySlice_l166_179_1};
  assign _zz_when_ArraySlice_l166_179_2 = (_zz_when_ArraySlice_l166_179_3 + _zz_when_ArraySlice_l166_179_7);
  assign _zz_when_ArraySlice_l166_179_3 = (realValue_0_179 - _zz_when_ArraySlice_l166_179_4);
  assign _zz_when_ArraySlice_l166_179_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_179_5);
  assign _zz_when_ArraySlice_l166_179_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_179_5 = {2'd0, _zz_when_ArraySlice_l166_179_6};
  assign _zz_when_ArraySlice_l166_179_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_180 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_180_1);
  assign _zz_when_ArraySlice_l158_180_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_180_1 = {1'd0, _zz_when_ArraySlice_l158_180_2};
  assign _zz_when_ArraySlice_l158_180_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_180_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_180 = {1'd0, _zz_when_ArraySlice_l159_180_1};
  assign _zz_when_ArraySlice_l159_180_2 = (_zz_when_ArraySlice_l159_180_3 - _zz_when_ArraySlice_l159_180_4);
  assign _zz_when_ArraySlice_l159_180_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_180_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_180_5);
  assign _zz_when_ArraySlice_l159_180_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_180_5 = {1'd0, _zz_when_ArraySlice_l159_180_6};
  assign _zz__zz_realValue_0_180 = {1'd0, wReg};
  assign _zz__zz_realValue_0_180_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_180_1 = (_zz_realValue_0_180_2 + _zz_realValue_0_180_3);
  assign _zz_realValue_0_180_2 = {1'd0, wReg};
  assign _zz_realValue_0_180_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_180_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_180 = {1'd0, _zz_when_ArraySlice_l166_180_1};
  assign _zz_when_ArraySlice_l166_180_2 = (_zz_when_ArraySlice_l166_180_3 + _zz_when_ArraySlice_l166_180_7);
  assign _zz_when_ArraySlice_l166_180_3 = (realValue_0_180 - _zz_when_ArraySlice_l166_180_4);
  assign _zz_when_ArraySlice_l166_180_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_180_5);
  assign _zz_when_ArraySlice_l166_180_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_180_5 = {1'd0, _zz_when_ArraySlice_l166_180_6};
  assign _zz_when_ArraySlice_l166_180_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_181 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_181_1);
  assign _zz_when_ArraySlice_l158_181_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_181_1 = {1'd0, _zz_when_ArraySlice_l158_181_2};
  assign _zz_when_ArraySlice_l158_181_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_181_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_181 = {2'd0, _zz_when_ArraySlice_l159_181_1};
  assign _zz_when_ArraySlice_l159_181_2 = (_zz_when_ArraySlice_l159_181_3 - _zz_when_ArraySlice_l159_181_4);
  assign _zz_when_ArraySlice_l159_181_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_181_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_181_5);
  assign _zz_when_ArraySlice_l159_181_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_181_5 = {1'd0, _zz_when_ArraySlice_l159_181_6};
  assign _zz__zz_realValue_0_181 = {1'd0, wReg};
  assign _zz__zz_realValue_0_181_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_181_1 = (_zz_realValue_0_181_2 + _zz_realValue_0_181_3);
  assign _zz_realValue_0_181_2 = {1'd0, wReg};
  assign _zz_realValue_0_181_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_181_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_181 = {2'd0, _zz_when_ArraySlice_l166_181_1};
  assign _zz_when_ArraySlice_l166_181_2 = (_zz_when_ArraySlice_l166_181_3 + _zz_when_ArraySlice_l166_181_7);
  assign _zz_when_ArraySlice_l166_181_3 = (realValue_0_181 - _zz_when_ArraySlice_l166_181_4);
  assign _zz_when_ArraySlice_l166_181_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_181_5);
  assign _zz_when_ArraySlice_l166_181_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_181_5 = {1'd0, _zz_when_ArraySlice_l166_181_6};
  assign _zz_when_ArraySlice_l166_181_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_182 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_182_1);
  assign _zz_when_ArraySlice_l158_182_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_182_1 = {1'd0, _zz_when_ArraySlice_l158_182_2};
  assign _zz_when_ArraySlice_l158_182_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_182_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_182 = {2'd0, _zz_when_ArraySlice_l159_182_1};
  assign _zz_when_ArraySlice_l159_182_2 = (_zz_when_ArraySlice_l159_182_3 - _zz_when_ArraySlice_l159_182_4);
  assign _zz_when_ArraySlice_l159_182_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_182_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_182_5);
  assign _zz_when_ArraySlice_l159_182_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_182_5 = {1'd0, _zz_when_ArraySlice_l159_182_6};
  assign _zz__zz_realValue_0_182 = {1'd0, wReg};
  assign _zz__zz_realValue_0_182_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_182_1 = (_zz_realValue_0_182_2 + _zz_realValue_0_182_3);
  assign _zz_realValue_0_182_2 = {1'd0, wReg};
  assign _zz_realValue_0_182_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_182_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_182 = {2'd0, _zz_when_ArraySlice_l166_182_1};
  assign _zz_when_ArraySlice_l166_182_2 = (_zz_when_ArraySlice_l166_182_3 + _zz_when_ArraySlice_l166_182_7);
  assign _zz_when_ArraySlice_l166_182_3 = (realValue_0_182 - _zz_when_ArraySlice_l166_182_4);
  assign _zz_when_ArraySlice_l166_182_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_182_5);
  assign _zz_when_ArraySlice_l166_182_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_182_5 = {1'd0, _zz_when_ArraySlice_l166_182_6};
  assign _zz_when_ArraySlice_l166_182_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_183 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_183_1);
  assign _zz_when_ArraySlice_l158_183_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_183_1 = {1'd0, _zz_when_ArraySlice_l158_183_2};
  assign _zz_when_ArraySlice_l158_183_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_183_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_183 = {3'd0, _zz_when_ArraySlice_l159_183_1};
  assign _zz_when_ArraySlice_l159_183_2 = (_zz_when_ArraySlice_l159_183_3 - _zz_when_ArraySlice_l159_183_4);
  assign _zz_when_ArraySlice_l159_183_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_183_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_183_5);
  assign _zz_when_ArraySlice_l159_183_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_183_5 = {1'd0, _zz_when_ArraySlice_l159_183_6};
  assign _zz__zz_realValue_0_183 = {1'd0, wReg};
  assign _zz__zz_realValue_0_183_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_183_1 = (_zz_realValue_0_183_2 + _zz_realValue_0_183_3);
  assign _zz_realValue_0_183_2 = {1'd0, wReg};
  assign _zz_realValue_0_183_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_183_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_183 = {3'd0, _zz_when_ArraySlice_l166_183_1};
  assign _zz_when_ArraySlice_l166_183_2 = (_zz_when_ArraySlice_l166_183_3 + _zz_when_ArraySlice_l166_183_7);
  assign _zz_when_ArraySlice_l166_183_3 = (realValue_0_183 - _zz_when_ArraySlice_l166_183_4);
  assign _zz_when_ArraySlice_l166_183_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_183_5);
  assign _zz_when_ArraySlice_l166_183_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_183_5 = {1'd0, _zz_when_ArraySlice_l166_183_6};
  assign _zz_when_ArraySlice_l166_183_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l403_7_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l403_7_2 = (_zz_when_ArraySlice_l403_7_3 + _zz_when_ArraySlice_l403_7_7);
  assign _zz_when_ArraySlice_l403_7_3 = (_zz_when_ArraySlice_l403_7_4 + 8'h01);
  assign _zz_when_ArraySlice_l403_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l403_7_5);
  assign _zz_when_ArraySlice_l403_7_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l403_7_5 = {1'd0, _zz_when_ArraySlice_l403_7_6};
  assign _zz_when_ArraySlice_l403_7_8 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l403_7_7 = {1'd0, _zz_when_ArraySlice_l403_7_8};
  assign _zz_when_ArraySlice_l406_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l406_7_1 = (_zz_when_ArraySlice_l406_7_2 + 8'h01);
  assign _zz_when_ArraySlice_l406_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l406_7_3);
  assign _zz_when_ArraySlice_l406_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l406_7_3 = {1'd0, _zz_when_ArraySlice_l406_7_4};
  assign _zz_selectReadFifo_7_6 = (selectReadFifo_7 + _zz_selectReadFifo_7_7);
  assign _zz_selectReadFifo_7_8 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_7 = {1'd0, _zz_selectReadFifo_7_8};
  assign _zz_when_ArraySlice_l413_7 = (_zz_when_ArraySlice_l413_7_1 % aReg);
  assign _zz_when_ArraySlice_l413_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l417_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l417_7_3);
  assign _zz_when_ArraySlice_l417_7_1 = _zz_when_ArraySlice_l417_7_2[6:0];
  assign _zz_when_ArraySlice_l417_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l417_7_3 = {1'd0, _zz_when_ArraySlice_l417_7_4};
  assign _zz_when_ArraySlice_l418_7_1 = (_zz_when_ArraySlice_l418_7_2 - _zz_when_ArraySlice_l418_7_3);
  assign _zz_when_ArraySlice_l418_7 = {5'd0, _zz_when_ArraySlice_l418_7_1};
  assign _zz_when_ArraySlice_l418_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l418_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l418_7_3 = {7'd0, _zz_when_ArraySlice_l418_7_4};
  assign _zz__zz_realValue1_0_22 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_22_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_22_1 = (_zz_realValue1_0_22_2 + _zz_realValue1_0_22_3);
  assign _zz_realValue1_0_22_2 = {1'd0, hReg};
  assign _zz_realValue1_0_22_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l420_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l420_7 = {1'd0, _zz_when_ArraySlice_l420_7_1};
  assign _zz_when_ArraySlice_l420_7_2 = (realValue1_0_22 / aReg);
  assign _zz_selectReadFifo_7_9 = (selectReadFifo_7 - _zz_selectReadFifo_7_10);
  assign _zz_selectReadFifo_7_10 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_184 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_184_1);
  assign _zz_when_ArraySlice_l158_184_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_184_1 = {4'd0, _zz_when_ArraySlice_l158_184_2};
  assign _zz_when_ArraySlice_l158_184_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_184 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_184_1 = (_zz_when_ArraySlice_l159_184_2 - _zz_when_ArraySlice_l159_184_3);
  assign _zz_when_ArraySlice_l159_184_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_184_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_184_4);
  assign _zz_when_ArraySlice_l159_184_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_184_4 = {4'd0, _zz_when_ArraySlice_l159_184_5};
  assign _zz__zz_realValue_0_184 = {1'd0, wReg};
  assign _zz__zz_realValue_0_184_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_184_1 = (_zz_realValue_0_184_2 + _zz_realValue_0_184_3);
  assign _zz_realValue_0_184_2 = {1'd0, wReg};
  assign _zz_realValue_0_184_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_184 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_184_1 = (_zz_when_ArraySlice_l166_184_2 + _zz_when_ArraySlice_l166_184_6);
  assign _zz_when_ArraySlice_l166_184_2 = (realValue_0_184 - _zz_when_ArraySlice_l166_184_3);
  assign _zz_when_ArraySlice_l166_184_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_184_4);
  assign _zz_when_ArraySlice_l166_184_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_184_4 = {4'd0, _zz_when_ArraySlice_l166_184_5};
  assign _zz_when_ArraySlice_l166_184_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_185 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_185_1);
  assign _zz_when_ArraySlice_l158_185_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_185_1 = {3'd0, _zz_when_ArraySlice_l158_185_2};
  assign _zz_when_ArraySlice_l158_185_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_185_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_185 = {1'd0, _zz_when_ArraySlice_l159_185_1};
  assign _zz_when_ArraySlice_l159_185_2 = (_zz_when_ArraySlice_l159_185_3 - _zz_when_ArraySlice_l159_185_4);
  assign _zz_when_ArraySlice_l159_185_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_185_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_185_5);
  assign _zz_when_ArraySlice_l159_185_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_185_5 = {3'd0, _zz_when_ArraySlice_l159_185_6};
  assign _zz__zz_realValue_0_185 = {1'd0, wReg};
  assign _zz__zz_realValue_0_185_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_185_1 = (_zz_realValue_0_185_2 + _zz_realValue_0_185_3);
  assign _zz_realValue_0_185_2 = {1'd0, wReg};
  assign _zz_realValue_0_185_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_185_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_185 = {1'd0, _zz_when_ArraySlice_l166_185_1};
  assign _zz_when_ArraySlice_l166_185_2 = (_zz_when_ArraySlice_l166_185_3 + _zz_when_ArraySlice_l166_185_7);
  assign _zz_when_ArraySlice_l166_185_3 = (realValue_0_185 - _zz_when_ArraySlice_l166_185_4);
  assign _zz_when_ArraySlice_l166_185_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_185_5);
  assign _zz_when_ArraySlice_l166_185_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_185_5 = {3'd0, _zz_when_ArraySlice_l166_185_6};
  assign _zz_when_ArraySlice_l166_185_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_186 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_186_1);
  assign _zz_when_ArraySlice_l158_186_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_186_1 = {2'd0, _zz_when_ArraySlice_l158_186_2};
  assign _zz_when_ArraySlice_l158_186_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_186_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_186 = {1'd0, _zz_when_ArraySlice_l159_186_1};
  assign _zz_when_ArraySlice_l159_186_2 = (_zz_when_ArraySlice_l159_186_3 - _zz_when_ArraySlice_l159_186_4);
  assign _zz_when_ArraySlice_l159_186_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_186_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_186_5);
  assign _zz_when_ArraySlice_l159_186_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_186_5 = {2'd0, _zz_when_ArraySlice_l159_186_6};
  assign _zz__zz_realValue_0_186 = {1'd0, wReg};
  assign _zz__zz_realValue_0_186_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_186_1 = (_zz_realValue_0_186_2 + _zz_realValue_0_186_3);
  assign _zz_realValue_0_186_2 = {1'd0, wReg};
  assign _zz_realValue_0_186_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_186_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_186 = {1'd0, _zz_when_ArraySlice_l166_186_1};
  assign _zz_when_ArraySlice_l166_186_2 = (_zz_when_ArraySlice_l166_186_3 + _zz_when_ArraySlice_l166_186_7);
  assign _zz_when_ArraySlice_l166_186_3 = (realValue_0_186 - _zz_when_ArraySlice_l166_186_4);
  assign _zz_when_ArraySlice_l166_186_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_186_5);
  assign _zz_when_ArraySlice_l166_186_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_186_5 = {2'd0, _zz_when_ArraySlice_l166_186_6};
  assign _zz_when_ArraySlice_l166_186_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_187 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_187_1);
  assign _zz_when_ArraySlice_l158_187_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_187_1 = {2'd0, _zz_when_ArraySlice_l158_187_2};
  assign _zz_when_ArraySlice_l158_187_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_187_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_187 = {1'd0, _zz_when_ArraySlice_l159_187_1};
  assign _zz_when_ArraySlice_l159_187_2 = (_zz_when_ArraySlice_l159_187_3 - _zz_when_ArraySlice_l159_187_4);
  assign _zz_when_ArraySlice_l159_187_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_187_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_187_5);
  assign _zz_when_ArraySlice_l159_187_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_187_5 = {2'd0, _zz_when_ArraySlice_l159_187_6};
  assign _zz__zz_realValue_0_187 = {1'd0, wReg};
  assign _zz__zz_realValue_0_187_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_187_1 = (_zz_realValue_0_187_2 + _zz_realValue_0_187_3);
  assign _zz_realValue_0_187_2 = {1'd0, wReg};
  assign _zz_realValue_0_187_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_187_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_187 = {1'd0, _zz_when_ArraySlice_l166_187_1};
  assign _zz_when_ArraySlice_l166_187_2 = (_zz_when_ArraySlice_l166_187_3 + _zz_when_ArraySlice_l166_187_7);
  assign _zz_when_ArraySlice_l166_187_3 = (realValue_0_187 - _zz_when_ArraySlice_l166_187_4);
  assign _zz_when_ArraySlice_l166_187_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_187_5);
  assign _zz_when_ArraySlice_l166_187_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_187_5 = {2'd0, _zz_when_ArraySlice_l166_187_6};
  assign _zz_when_ArraySlice_l166_187_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_188 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_188_1);
  assign _zz_when_ArraySlice_l158_188_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_188_1 = {1'd0, _zz_when_ArraySlice_l158_188_2};
  assign _zz_when_ArraySlice_l158_188_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_188_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_188 = {1'd0, _zz_when_ArraySlice_l159_188_1};
  assign _zz_when_ArraySlice_l159_188_2 = (_zz_when_ArraySlice_l159_188_3 - _zz_when_ArraySlice_l159_188_4);
  assign _zz_when_ArraySlice_l159_188_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_188_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_188_5);
  assign _zz_when_ArraySlice_l159_188_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_188_5 = {1'd0, _zz_when_ArraySlice_l159_188_6};
  assign _zz__zz_realValue_0_188 = {1'd0, wReg};
  assign _zz__zz_realValue_0_188_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_188_1 = (_zz_realValue_0_188_2 + _zz_realValue_0_188_3);
  assign _zz_realValue_0_188_2 = {1'd0, wReg};
  assign _zz_realValue_0_188_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_188_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_188 = {1'd0, _zz_when_ArraySlice_l166_188_1};
  assign _zz_when_ArraySlice_l166_188_2 = (_zz_when_ArraySlice_l166_188_3 + _zz_when_ArraySlice_l166_188_7);
  assign _zz_when_ArraySlice_l166_188_3 = (realValue_0_188 - _zz_when_ArraySlice_l166_188_4);
  assign _zz_when_ArraySlice_l166_188_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_188_5);
  assign _zz_when_ArraySlice_l166_188_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_188_5 = {1'd0, _zz_when_ArraySlice_l166_188_6};
  assign _zz_when_ArraySlice_l166_188_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_189 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_189_1);
  assign _zz_when_ArraySlice_l158_189_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_189_1 = {1'd0, _zz_when_ArraySlice_l158_189_2};
  assign _zz_when_ArraySlice_l158_189_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_189_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_189 = {2'd0, _zz_when_ArraySlice_l159_189_1};
  assign _zz_when_ArraySlice_l159_189_2 = (_zz_when_ArraySlice_l159_189_3 - _zz_when_ArraySlice_l159_189_4);
  assign _zz_when_ArraySlice_l159_189_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_189_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_189_5);
  assign _zz_when_ArraySlice_l159_189_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_189_5 = {1'd0, _zz_when_ArraySlice_l159_189_6};
  assign _zz__zz_realValue_0_189 = {1'd0, wReg};
  assign _zz__zz_realValue_0_189_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_189_1 = (_zz_realValue_0_189_2 + _zz_realValue_0_189_3);
  assign _zz_realValue_0_189_2 = {1'd0, wReg};
  assign _zz_realValue_0_189_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_189_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_189 = {2'd0, _zz_when_ArraySlice_l166_189_1};
  assign _zz_when_ArraySlice_l166_189_2 = (_zz_when_ArraySlice_l166_189_3 + _zz_when_ArraySlice_l166_189_7);
  assign _zz_when_ArraySlice_l166_189_3 = (realValue_0_189 - _zz_when_ArraySlice_l166_189_4);
  assign _zz_when_ArraySlice_l166_189_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_189_5);
  assign _zz_when_ArraySlice_l166_189_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_189_5 = {1'd0, _zz_when_ArraySlice_l166_189_6};
  assign _zz_when_ArraySlice_l166_189_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_190 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_190_1);
  assign _zz_when_ArraySlice_l158_190_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_190_1 = {1'd0, _zz_when_ArraySlice_l158_190_2};
  assign _zz_when_ArraySlice_l158_190_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_190_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_190 = {2'd0, _zz_when_ArraySlice_l159_190_1};
  assign _zz_when_ArraySlice_l159_190_2 = (_zz_when_ArraySlice_l159_190_3 - _zz_when_ArraySlice_l159_190_4);
  assign _zz_when_ArraySlice_l159_190_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_190_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_190_5);
  assign _zz_when_ArraySlice_l159_190_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_190_5 = {1'd0, _zz_when_ArraySlice_l159_190_6};
  assign _zz__zz_realValue_0_190 = {1'd0, wReg};
  assign _zz__zz_realValue_0_190_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_190_1 = (_zz_realValue_0_190_2 + _zz_realValue_0_190_3);
  assign _zz_realValue_0_190_2 = {1'd0, wReg};
  assign _zz_realValue_0_190_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_190_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_190 = {2'd0, _zz_when_ArraySlice_l166_190_1};
  assign _zz_when_ArraySlice_l166_190_2 = (_zz_when_ArraySlice_l166_190_3 + _zz_when_ArraySlice_l166_190_7);
  assign _zz_when_ArraySlice_l166_190_3 = (realValue_0_190 - _zz_when_ArraySlice_l166_190_4);
  assign _zz_when_ArraySlice_l166_190_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_190_5);
  assign _zz_when_ArraySlice_l166_190_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_190_5 = {1'd0, _zz_when_ArraySlice_l166_190_6};
  assign _zz_when_ArraySlice_l166_190_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_191 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_191_1);
  assign _zz_when_ArraySlice_l158_191_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_191_1 = {1'd0, _zz_when_ArraySlice_l158_191_2};
  assign _zz_when_ArraySlice_l158_191_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_191_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_191 = {3'd0, _zz_when_ArraySlice_l159_191_1};
  assign _zz_when_ArraySlice_l159_191_2 = (_zz_when_ArraySlice_l159_191_3 - _zz_when_ArraySlice_l159_191_4);
  assign _zz_when_ArraySlice_l159_191_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_191_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_191_5);
  assign _zz_when_ArraySlice_l159_191_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_191_5 = {1'd0, _zz_when_ArraySlice_l159_191_6};
  assign _zz__zz_realValue_0_191 = {1'd0, wReg};
  assign _zz__zz_realValue_0_191_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_191_1 = (_zz_realValue_0_191_2 + _zz_realValue_0_191_3);
  assign _zz_realValue_0_191_2 = {1'd0, wReg};
  assign _zz_realValue_0_191_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_191_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_191 = {3'd0, _zz_when_ArraySlice_l166_191_1};
  assign _zz_when_ArraySlice_l166_191_2 = (_zz_when_ArraySlice_l166_191_3 + _zz_when_ArraySlice_l166_191_7);
  assign _zz_when_ArraySlice_l166_191_3 = (realValue_0_191 - _zz_when_ArraySlice_l166_191_4);
  assign _zz_when_ArraySlice_l166_191_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_191_5);
  assign _zz_when_ArraySlice_l166_191_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_191_5 = {1'd0, _zz_when_ArraySlice_l166_191_6};
  assign _zz_when_ArraySlice_l166_191_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l428_7_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l428_7_2 = (_zz_when_ArraySlice_l428_7_3 + _zz_when_ArraySlice_l428_7_7);
  assign _zz_when_ArraySlice_l428_7_3 = (_zz_when_ArraySlice_l428_7_4 + 8'h01);
  assign _zz_when_ArraySlice_l428_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l428_7_5);
  assign _zz_when_ArraySlice_l428_7_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l428_7_5 = {1'd0, _zz_when_ArraySlice_l428_7_6};
  assign _zz_when_ArraySlice_l428_7_8 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l428_7_7 = {1'd0, _zz_when_ArraySlice_l428_7_8};
  assign _zz_when_ArraySlice_l431_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l431_7_1 = (_zz_when_ArraySlice_l431_7_2 + 8'h01);
  assign _zz_when_ArraySlice_l431_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l431_7_3);
  assign _zz_when_ArraySlice_l431_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l431_7_3 = {1'd0, _zz_when_ArraySlice_l431_7_4};
  assign _zz_selectReadFifo_7_11 = (selectReadFifo_7 + _zz_selectReadFifo_7_12);
  assign _zz_selectReadFifo_7_13 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_12 = {1'd0, _zz_selectReadFifo_7_13};
  assign _zz_when_ArraySlice_l438_7 = (_zz_when_ArraySlice_l438_7_1 % aReg);
  assign _zz_when_ArraySlice_l438_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l449_7_1 = (_zz_when_ArraySlice_l449_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l449_7 = {5'd0, _zz_when_ArraySlice_l449_7_1};
  assign _zz_when_ArraySlice_l449_7_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_23 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_23_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_23_1 = (_zz_realValue1_0_23_2 + _zz_realValue1_0_23_3);
  assign _zz_realValue1_0_23_2 = {1'd0, hReg};
  assign _zz_realValue1_0_23_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l450_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l450_7 = {1'd0, _zz_when_ArraySlice_l450_7_1};
  assign _zz_when_ArraySlice_l450_7_2 = (realValue1_0_23 / aReg);
  assign _zz_selectReadFifo_7_14 = (selectReadFifo_7 - _zz_selectReadFifo_7_15);
  assign _zz_selectReadFifo_7_15 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_192 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_192_1);
  assign _zz_when_ArraySlice_l158_192_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_192_1 = {4'd0, _zz_when_ArraySlice_l158_192_2};
  assign _zz_when_ArraySlice_l158_192_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_192 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_192_1 = (_zz_when_ArraySlice_l159_192_2 - _zz_when_ArraySlice_l159_192_3);
  assign _zz_when_ArraySlice_l159_192_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_192_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_192_4);
  assign _zz_when_ArraySlice_l159_192_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_192_4 = {4'd0, _zz_when_ArraySlice_l159_192_5};
  assign _zz__zz_realValue_0_192 = {1'd0, wReg};
  assign _zz__zz_realValue_0_192_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_192_1 = (_zz_realValue_0_192_2 + _zz_realValue_0_192_3);
  assign _zz_realValue_0_192_2 = {1'd0, wReg};
  assign _zz_realValue_0_192_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_192 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_192_1 = (_zz_when_ArraySlice_l166_192_2 + _zz_when_ArraySlice_l166_192_6);
  assign _zz_when_ArraySlice_l166_192_2 = (realValue_0_192 - _zz_when_ArraySlice_l166_192_3);
  assign _zz_when_ArraySlice_l166_192_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_192_4);
  assign _zz_when_ArraySlice_l166_192_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_192_4 = {4'd0, _zz_when_ArraySlice_l166_192_5};
  assign _zz_when_ArraySlice_l166_192_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_193 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_193_1);
  assign _zz_when_ArraySlice_l158_193_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_193_1 = {3'd0, _zz_when_ArraySlice_l158_193_2};
  assign _zz_when_ArraySlice_l158_193_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_193_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_193 = {1'd0, _zz_when_ArraySlice_l159_193_1};
  assign _zz_when_ArraySlice_l159_193_2 = (_zz_when_ArraySlice_l159_193_3 - _zz_when_ArraySlice_l159_193_4);
  assign _zz_when_ArraySlice_l159_193_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_193_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_193_5);
  assign _zz_when_ArraySlice_l159_193_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_193_5 = {3'd0, _zz_when_ArraySlice_l159_193_6};
  assign _zz__zz_realValue_0_193 = {1'd0, wReg};
  assign _zz__zz_realValue_0_193_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_193_1 = (_zz_realValue_0_193_2 + _zz_realValue_0_193_3);
  assign _zz_realValue_0_193_2 = {1'd0, wReg};
  assign _zz_realValue_0_193_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_193_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_193 = {1'd0, _zz_when_ArraySlice_l166_193_1};
  assign _zz_when_ArraySlice_l166_193_2 = (_zz_when_ArraySlice_l166_193_3 + _zz_when_ArraySlice_l166_193_7);
  assign _zz_when_ArraySlice_l166_193_3 = (realValue_0_193 - _zz_when_ArraySlice_l166_193_4);
  assign _zz_when_ArraySlice_l166_193_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_193_5);
  assign _zz_when_ArraySlice_l166_193_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_193_5 = {3'd0, _zz_when_ArraySlice_l166_193_6};
  assign _zz_when_ArraySlice_l166_193_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_194 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_194_1);
  assign _zz_when_ArraySlice_l158_194_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_194_1 = {2'd0, _zz_when_ArraySlice_l158_194_2};
  assign _zz_when_ArraySlice_l158_194_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_194_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_194 = {1'd0, _zz_when_ArraySlice_l159_194_1};
  assign _zz_when_ArraySlice_l159_194_2 = (_zz_when_ArraySlice_l159_194_3 - _zz_when_ArraySlice_l159_194_4);
  assign _zz_when_ArraySlice_l159_194_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_194_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_194_5);
  assign _zz_when_ArraySlice_l159_194_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_194_5 = {2'd0, _zz_when_ArraySlice_l159_194_6};
  assign _zz__zz_realValue_0_194 = {1'd0, wReg};
  assign _zz__zz_realValue_0_194_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_194_1 = (_zz_realValue_0_194_2 + _zz_realValue_0_194_3);
  assign _zz_realValue_0_194_2 = {1'd0, wReg};
  assign _zz_realValue_0_194_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_194_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_194 = {1'd0, _zz_when_ArraySlice_l166_194_1};
  assign _zz_when_ArraySlice_l166_194_2 = (_zz_when_ArraySlice_l166_194_3 + _zz_when_ArraySlice_l166_194_7);
  assign _zz_when_ArraySlice_l166_194_3 = (realValue_0_194 - _zz_when_ArraySlice_l166_194_4);
  assign _zz_when_ArraySlice_l166_194_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_194_5);
  assign _zz_when_ArraySlice_l166_194_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_194_5 = {2'd0, _zz_when_ArraySlice_l166_194_6};
  assign _zz_when_ArraySlice_l166_194_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_195 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_195_1);
  assign _zz_when_ArraySlice_l158_195_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_195_1 = {2'd0, _zz_when_ArraySlice_l158_195_2};
  assign _zz_when_ArraySlice_l158_195_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_195_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_195 = {1'd0, _zz_when_ArraySlice_l159_195_1};
  assign _zz_when_ArraySlice_l159_195_2 = (_zz_when_ArraySlice_l159_195_3 - _zz_when_ArraySlice_l159_195_4);
  assign _zz_when_ArraySlice_l159_195_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_195_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_195_5);
  assign _zz_when_ArraySlice_l159_195_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_195_5 = {2'd0, _zz_when_ArraySlice_l159_195_6};
  assign _zz__zz_realValue_0_195 = {1'd0, wReg};
  assign _zz__zz_realValue_0_195_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_195_1 = (_zz_realValue_0_195_2 + _zz_realValue_0_195_3);
  assign _zz_realValue_0_195_2 = {1'd0, wReg};
  assign _zz_realValue_0_195_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_195_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_195 = {1'd0, _zz_when_ArraySlice_l166_195_1};
  assign _zz_when_ArraySlice_l166_195_2 = (_zz_when_ArraySlice_l166_195_3 + _zz_when_ArraySlice_l166_195_7);
  assign _zz_when_ArraySlice_l166_195_3 = (realValue_0_195 - _zz_when_ArraySlice_l166_195_4);
  assign _zz_when_ArraySlice_l166_195_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_195_5);
  assign _zz_when_ArraySlice_l166_195_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_195_5 = {2'd0, _zz_when_ArraySlice_l166_195_6};
  assign _zz_when_ArraySlice_l166_195_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_196 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_196_1);
  assign _zz_when_ArraySlice_l158_196_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_196_1 = {1'd0, _zz_when_ArraySlice_l158_196_2};
  assign _zz_when_ArraySlice_l158_196_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_196_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_196 = {1'd0, _zz_when_ArraySlice_l159_196_1};
  assign _zz_when_ArraySlice_l159_196_2 = (_zz_when_ArraySlice_l159_196_3 - _zz_when_ArraySlice_l159_196_4);
  assign _zz_when_ArraySlice_l159_196_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_196_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_196_5);
  assign _zz_when_ArraySlice_l159_196_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_196_5 = {1'd0, _zz_when_ArraySlice_l159_196_6};
  assign _zz__zz_realValue_0_196 = {1'd0, wReg};
  assign _zz__zz_realValue_0_196_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_196_1 = (_zz_realValue_0_196_2 + _zz_realValue_0_196_3);
  assign _zz_realValue_0_196_2 = {1'd0, wReg};
  assign _zz_realValue_0_196_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_196_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_196 = {1'd0, _zz_when_ArraySlice_l166_196_1};
  assign _zz_when_ArraySlice_l166_196_2 = (_zz_when_ArraySlice_l166_196_3 + _zz_when_ArraySlice_l166_196_7);
  assign _zz_when_ArraySlice_l166_196_3 = (realValue_0_196 - _zz_when_ArraySlice_l166_196_4);
  assign _zz_when_ArraySlice_l166_196_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_196_5);
  assign _zz_when_ArraySlice_l166_196_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_196_5 = {1'd0, _zz_when_ArraySlice_l166_196_6};
  assign _zz_when_ArraySlice_l166_196_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_197 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_197_1);
  assign _zz_when_ArraySlice_l158_197_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_197_1 = {1'd0, _zz_when_ArraySlice_l158_197_2};
  assign _zz_when_ArraySlice_l158_197_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_197_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_197 = {2'd0, _zz_when_ArraySlice_l159_197_1};
  assign _zz_when_ArraySlice_l159_197_2 = (_zz_when_ArraySlice_l159_197_3 - _zz_when_ArraySlice_l159_197_4);
  assign _zz_when_ArraySlice_l159_197_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_197_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_197_5);
  assign _zz_when_ArraySlice_l159_197_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_197_5 = {1'd0, _zz_when_ArraySlice_l159_197_6};
  assign _zz__zz_realValue_0_197 = {1'd0, wReg};
  assign _zz__zz_realValue_0_197_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_197_1 = (_zz_realValue_0_197_2 + _zz_realValue_0_197_3);
  assign _zz_realValue_0_197_2 = {1'd0, wReg};
  assign _zz_realValue_0_197_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_197_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_197 = {2'd0, _zz_when_ArraySlice_l166_197_1};
  assign _zz_when_ArraySlice_l166_197_2 = (_zz_when_ArraySlice_l166_197_3 + _zz_when_ArraySlice_l166_197_7);
  assign _zz_when_ArraySlice_l166_197_3 = (realValue_0_197 - _zz_when_ArraySlice_l166_197_4);
  assign _zz_when_ArraySlice_l166_197_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_197_5);
  assign _zz_when_ArraySlice_l166_197_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_197_5 = {1'd0, _zz_when_ArraySlice_l166_197_6};
  assign _zz_when_ArraySlice_l166_197_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_198 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_198_1);
  assign _zz_when_ArraySlice_l158_198_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_198_1 = {1'd0, _zz_when_ArraySlice_l158_198_2};
  assign _zz_when_ArraySlice_l158_198_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_198_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_198 = {2'd0, _zz_when_ArraySlice_l159_198_1};
  assign _zz_when_ArraySlice_l159_198_2 = (_zz_when_ArraySlice_l159_198_3 - _zz_when_ArraySlice_l159_198_4);
  assign _zz_when_ArraySlice_l159_198_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_198_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_198_5);
  assign _zz_when_ArraySlice_l159_198_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_198_5 = {1'd0, _zz_when_ArraySlice_l159_198_6};
  assign _zz__zz_realValue_0_198 = {1'd0, wReg};
  assign _zz__zz_realValue_0_198_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_198_1 = (_zz_realValue_0_198_2 + _zz_realValue_0_198_3);
  assign _zz_realValue_0_198_2 = {1'd0, wReg};
  assign _zz_realValue_0_198_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_198_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_198 = {2'd0, _zz_when_ArraySlice_l166_198_1};
  assign _zz_when_ArraySlice_l166_198_2 = (_zz_when_ArraySlice_l166_198_3 + _zz_when_ArraySlice_l166_198_7);
  assign _zz_when_ArraySlice_l166_198_3 = (realValue_0_198 - _zz_when_ArraySlice_l166_198_4);
  assign _zz_when_ArraySlice_l166_198_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_198_5);
  assign _zz_when_ArraySlice_l166_198_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_198_5 = {1'd0, _zz_when_ArraySlice_l166_198_6};
  assign _zz_when_ArraySlice_l166_198_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_199 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_199_1);
  assign _zz_when_ArraySlice_l158_199_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_199_1 = {1'd0, _zz_when_ArraySlice_l158_199_2};
  assign _zz_when_ArraySlice_l158_199_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_199_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_199 = {3'd0, _zz_when_ArraySlice_l159_199_1};
  assign _zz_when_ArraySlice_l159_199_2 = (_zz_when_ArraySlice_l159_199_3 - _zz_when_ArraySlice_l159_199_4);
  assign _zz_when_ArraySlice_l159_199_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_199_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_199_5);
  assign _zz_when_ArraySlice_l159_199_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_199_5 = {1'd0, _zz_when_ArraySlice_l159_199_6};
  assign _zz__zz_realValue_0_199 = {1'd0, wReg};
  assign _zz__zz_realValue_0_199_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_199_1 = (_zz_realValue_0_199_2 + _zz_realValue_0_199_3);
  assign _zz_realValue_0_199_2 = {1'd0, wReg};
  assign _zz_realValue_0_199_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_199_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_199 = {3'd0, _zz_when_ArraySlice_l166_199_1};
  assign _zz_when_ArraySlice_l166_199_2 = (_zz_when_ArraySlice_l166_199_3 + _zz_when_ArraySlice_l166_199_7);
  assign _zz_when_ArraySlice_l166_199_3 = (realValue_0_199 - _zz_when_ArraySlice_l166_199_4);
  assign _zz_when_ArraySlice_l166_199_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_199_5);
  assign _zz_when_ArraySlice_l166_199_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_199_5 = {1'd0, _zz_when_ArraySlice_l166_199_6};
  assign _zz_when_ArraySlice_l166_199_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l461_7 = (_zz_when_ArraySlice_l461_7_1 % aReg);
  assign _zz_when_ArraySlice_l461_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l447_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l447_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l447_7_2);
  assign _zz_when_ArraySlice_l447_7_3 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l447_7_2 = {1'd0, _zz_when_ArraySlice_l447_7_3};
  assign _zz_when_ArraySlice_l468_7_1 = (_zz_when_ArraySlice_l468_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l468_7 = {5'd0, _zz_when_ArraySlice_l468_7_1};
  assign _zz_when_ArraySlice_l468_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l158_200 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_200_1);
  assign _zz_when_ArraySlice_l158_200_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_200_1 = {4'd0, _zz_when_ArraySlice_l158_200_2};
  assign _zz_when_ArraySlice_l158_200_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_200 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_200_1 = (_zz_when_ArraySlice_l159_200_2 - _zz_when_ArraySlice_l159_200_3);
  assign _zz_when_ArraySlice_l159_200_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_200_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_200_4);
  assign _zz_when_ArraySlice_l159_200_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_200_4 = {4'd0, _zz_when_ArraySlice_l159_200_5};
  assign _zz__zz_realValue_0_200 = {1'd0, wReg};
  assign _zz__zz_realValue_0_200_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_200_1 = (_zz_realValue_0_200_2 + _zz_realValue_0_200_3);
  assign _zz_realValue_0_200_2 = {1'd0, wReg};
  assign _zz_realValue_0_200_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_200 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_200_1 = (_zz_when_ArraySlice_l166_200_2 + _zz_when_ArraySlice_l166_200_6);
  assign _zz_when_ArraySlice_l166_200_2 = (realValue_0_200 - _zz_when_ArraySlice_l166_200_3);
  assign _zz_when_ArraySlice_l166_200_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_200_4);
  assign _zz_when_ArraySlice_l166_200_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_200_4 = {4'd0, _zz_when_ArraySlice_l166_200_5};
  assign _zz_when_ArraySlice_l166_200_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_201 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_201_1);
  assign _zz_when_ArraySlice_l158_201_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_201_1 = {3'd0, _zz_when_ArraySlice_l158_201_2};
  assign _zz_when_ArraySlice_l158_201_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_201_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_201 = {1'd0, _zz_when_ArraySlice_l159_201_1};
  assign _zz_when_ArraySlice_l159_201_2 = (_zz_when_ArraySlice_l159_201_3 - _zz_when_ArraySlice_l159_201_4);
  assign _zz_when_ArraySlice_l159_201_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_201_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_201_5);
  assign _zz_when_ArraySlice_l159_201_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_201_5 = {3'd0, _zz_when_ArraySlice_l159_201_6};
  assign _zz__zz_realValue_0_201 = {1'd0, wReg};
  assign _zz__zz_realValue_0_201_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_201_1 = (_zz_realValue_0_201_2 + _zz_realValue_0_201_3);
  assign _zz_realValue_0_201_2 = {1'd0, wReg};
  assign _zz_realValue_0_201_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_201_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_201 = {1'd0, _zz_when_ArraySlice_l166_201_1};
  assign _zz_when_ArraySlice_l166_201_2 = (_zz_when_ArraySlice_l166_201_3 + _zz_when_ArraySlice_l166_201_7);
  assign _zz_when_ArraySlice_l166_201_3 = (realValue_0_201 - _zz_when_ArraySlice_l166_201_4);
  assign _zz_when_ArraySlice_l166_201_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_201_5);
  assign _zz_when_ArraySlice_l166_201_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_201_5 = {3'd0, _zz_when_ArraySlice_l166_201_6};
  assign _zz_when_ArraySlice_l166_201_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_202 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_202_1);
  assign _zz_when_ArraySlice_l158_202_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_202_1 = {2'd0, _zz_when_ArraySlice_l158_202_2};
  assign _zz_when_ArraySlice_l158_202_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_202_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_202 = {1'd0, _zz_when_ArraySlice_l159_202_1};
  assign _zz_when_ArraySlice_l159_202_2 = (_zz_when_ArraySlice_l159_202_3 - _zz_when_ArraySlice_l159_202_4);
  assign _zz_when_ArraySlice_l159_202_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_202_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_202_5);
  assign _zz_when_ArraySlice_l159_202_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_202_5 = {2'd0, _zz_when_ArraySlice_l159_202_6};
  assign _zz__zz_realValue_0_202 = {1'd0, wReg};
  assign _zz__zz_realValue_0_202_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_202_1 = (_zz_realValue_0_202_2 + _zz_realValue_0_202_3);
  assign _zz_realValue_0_202_2 = {1'd0, wReg};
  assign _zz_realValue_0_202_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_202_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_202 = {1'd0, _zz_when_ArraySlice_l166_202_1};
  assign _zz_when_ArraySlice_l166_202_2 = (_zz_when_ArraySlice_l166_202_3 + _zz_when_ArraySlice_l166_202_7);
  assign _zz_when_ArraySlice_l166_202_3 = (realValue_0_202 - _zz_when_ArraySlice_l166_202_4);
  assign _zz_when_ArraySlice_l166_202_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_202_5);
  assign _zz_when_ArraySlice_l166_202_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_202_5 = {2'd0, _zz_when_ArraySlice_l166_202_6};
  assign _zz_when_ArraySlice_l166_202_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_203 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_203_1);
  assign _zz_when_ArraySlice_l158_203_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_203_1 = {2'd0, _zz_when_ArraySlice_l158_203_2};
  assign _zz_when_ArraySlice_l158_203_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_203_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_203 = {1'd0, _zz_when_ArraySlice_l159_203_1};
  assign _zz_when_ArraySlice_l159_203_2 = (_zz_when_ArraySlice_l159_203_3 - _zz_when_ArraySlice_l159_203_4);
  assign _zz_when_ArraySlice_l159_203_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_203_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_203_5);
  assign _zz_when_ArraySlice_l159_203_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_203_5 = {2'd0, _zz_when_ArraySlice_l159_203_6};
  assign _zz__zz_realValue_0_203 = {1'd0, wReg};
  assign _zz__zz_realValue_0_203_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_203_1 = (_zz_realValue_0_203_2 + _zz_realValue_0_203_3);
  assign _zz_realValue_0_203_2 = {1'd0, wReg};
  assign _zz_realValue_0_203_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_203_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_203 = {1'd0, _zz_when_ArraySlice_l166_203_1};
  assign _zz_when_ArraySlice_l166_203_2 = (_zz_when_ArraySlice_l166_203_3 + _zz_when_ArraySlice_l166_203_7);
  assign _zz_when_ArraySlice_l166_203_3 = (realValue_0_203 - _zz_when_ArraySlice_l166_203_4);
  assign _zz_when_ArraySlice_l166_203_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_203_5);
  assign _zz_when_ArraySlice_l166_203_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_203_5 = {2'd0, _zz_when_ArraySlice_l166_203_6};
  assign _zz_when_ArraySlice_l166_203_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_204 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_204_1);
  assign _zz_when_ArraySlice_l158_204_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_204_1 = {1'd0, _zz_when_ArraySlice_l158_204_2};
  assign _zz_when_ArraySlice_l158_204_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_204_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_204 = {1'd0, _zz_when_ArraySlice_l159_204_1};
  assign _zz_when_ArraySlice_l159_204_2 = (_zz_when_ArraySlice_l159_204_3 - _zz_when_ArraySlice_l159_204_4);
  assign _zz_when_ArraySlice_l159_204_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_204_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_204_5);
  assign _zz_when_ArraySlice_l159_204_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_204_5 = {1'd0, _zz_when_ArraySlice_l159_204_6};
  assign _zz__zz_realValue_0_204 = {1'd0, wReg};
  assign _zz__zz_realValue_0_204_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_204_1 = (_zz_realValue_0_204_2 + _zz_realValue_0_204_3);
  assign _zz_realValue_0_204_2 = {1'd0, wReg};
  assign _zz_realValue_0_204_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_204_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_204 = {1'd0, _zz_when_ArraySlice_l166_204_1};
  assign _zz_when_ArraySlice_l166_204_2 = (_zz_when_ArraySlice_l166_204_3 + _zz_when_ArraySlice_l166_204_7);
  assign _zz_when_ArraySlice_l166_204_3 = (realValue_0_204 - _zz_when_ArraySlice_l166_204_4);
  assign _zz_when_ArraySlice_l166_204_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_204_5);
  assign _zz_when_ArraySlice_l166_204_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_204_5 = {1'd0, _zz_when_ArraySlice_l166_204_6};
  assign _zz_when_ArraySlice_l166_204_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_205 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_205_1);
  assign _zz_when_ArraySlice_l158_205_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_205_1 = {1'd0, _zz_when_ArraySlice_l158_205_2};
  assign _zz_when_ArraySlice_l158_205_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_205_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_205 = {2'd0, _zz_when_ArraySlice_l159_205_1};
  assign _zz_when_ArraySlice_l159_205_2 = (_zz_when_ArraySlice_l159_205_3 - _zz_when_ArraySlice_l159_205_4);
  assign _zz_when_ArraySlice_l159_205_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_205_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_205_5);
  assign _zz_when_ArraySlice_l159_205_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_205_5 = {1'd0, _zz_when_ArraySlice_l159_205_6};
  assign _zz__zz_realValue_0_205 = {1'd0, wReg};
  assign _zz__zz_realValue_0_205_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_205_1 = (_zz_realValue_0_205_2 + _zz_realValue_0_205_3);
  assign _zz_realValue_0_205_2 = {1'd0, wReg};
  assign _zz_realValue_0_205_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_205_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_205 = {2'd0, _zz_when_ArraySlice_l166_205_1};
  assign _zz_when_ArraySlice_l166_205_2 = (_zz_when_ArraySlice_l166_205_3 + _zz_when_ArraySlice_l166_205_7);
  assign _zz_when_ArraySlice_l166_205_3 = (realValue_0_205 - _zz_when_ArraySlice_l166_205_4);
  assign _zz_when_ArraySlice_l166_205_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_205_5);
  assign _zz_when_ArraySlice_l166_205_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_205_5 = {1'd0, _zz_when_ArraySlice_l166_205_6};
  assign _zz_when_ArraySlice_l166_205_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_206 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_206_1);
  assign _zz_when_ArraySlice_l158_206_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_206_1 = {1'd0, _zz_when_ArraySlice_l158_206_2};
  assign _zz_when_ArraySlice_l158_206_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_206_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_206 = {2'd0, _zz_when_ArraySlice_l159_206_1};
  assign _zz_when_ArraySlice_l159_206_2 = (_zz_when_ArraySlice_l159_206_3 - _zz_when_ArraySlice_l159_206_4);
  assign _zz_when_ArraySlice_l159_206_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_206_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_206_5);
  assign _zz_when_ArraySlice_l159_206_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_206_5 = {1'd0, _zz_when_ArraySlice_l159_206_6};
  assign _zz__zz_realValue_0_206 = {1'd0, wReg};
  assign _zz__zz_realValue_0_206_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_206_1 = (_zz_realValue_0_206_2 + _zz_realValue_0_206_3);
  assign _zz_realValue_0_206_2 = {1'd0, wReg};
  assign _zz_realValue_0_206_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_206_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_206 = {2'd0, _zz_when_ArraySlice_l166_206_1};
  assign _zz_when_ArraySlice_l166_206_2 = (_zz_when_ArraySlice_l166_206_3 + _zz_when_ArraySlice_l166_206_7);
  assign _zz_when_ArraySlice_l166_206_3 = (realValue_0_206 - _zz_when_ArraySlice_l166_206_4);
  assign _zz_when_ArraySlice_l166_206_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_206_5);
  assign _zz_when_ArraySlice_l166_206_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_206_5 = {1'd0, _zz_when_ArraySlice_l166_206_6};
  assign _zz_when_ArraySlice_l166_206_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_207 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_207_1);
  assign _zz_when_ArraySlice_l158_207_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_207_1 = {1'd0, _zz_when_ArraySlice_l158_207_2};
  assign _zz_when_ArraySlice_l158_207_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_207_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_207 = {3'd0, _zz_when_ArraySlice_l159_207_1};
  assign _zz_when_ArraySlice_l159_207_2 = (_zz_when_ArraySlice_l159_207_3 - _zz_when_ArraySlice_l159_207_4);
  assign _zz_when_ArraySlice_l159_207_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_207_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_207_5);
  assign _zz_when_ArraySlice_l159_207_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_207_5 = {1'd0, _zz_when_ArraySlice_l159_207_6};
  assign _zz__zz_realValue_0_207 = {1'd0, wReg};
  assign _zz__zz_realValue_0_207_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_207_1 = (_zz_realValue_0_207_2 + _zz_realValue_0_207_3);
  assign _zz_realValue_0_207_2 = {1'd0, wReg};
  assign _zz_realValue_0_207_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_207_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_207 = {3'd0, _zz_when_ArraySlice_l166_207_1};
  assign _zz_when_ArraySlice_l166_207_2 = (_zz_when_ArraySlice_l166_207_3 + _zz_when_ArraySlice_l166_207_7);
  assign _zz_when_ArraySlice_l166_207_3 = (realValue_0_207 - _zz_when_ArraySlice_l166_207_4);
  assign _zz_when_ArraySlice_l166_207_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_207_5);
  assign _zz_when_ArraySlice_l166_207_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_207_5 = {1'd0, _zz_when_ArraySlice_l166_207_6};
  assign _zz_when_ArraySlice_l166_207_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l233 = (selectReadFifo_0 + _zz_when_ArraySlice_l233_1);
  assign _zz_when_ArraySlice_l233_2 = 4'b0000;
  assign _zz_when_ArraySlice_l233_1 = {4'd0, _zz_when_ArraySlice_l233_2};
  assign _zz_when_ArraySlice_l233_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l234_3);
  assign _zz_when_ArraySlice_l234_1 = _zz_when_ArraySlice_l234_2[6:0];
  assign _zz_when_ArraySlice_l234_4 = 4'b0000;
  assign _zz_when_ArraySlice_l234_3 = {4'd0, _zz_when_ArraySlice_l234_4};
  assign _zz__zz_outputStreamArrayData_0_valid_1_2 = 4'b0000;
  assign _zz__zz_outputStreamArrayData_0_valid_1_1 = {4'd0, _zz__zz_outputStreamArrayData_0_valid_1_2};
  assign _zz__zz_11 = _zz_outputStreamArrayData_0_valid_1[6:0];
  assign _zz_outputStreamArrayData_0_valid_5 = _zz_outputStreamArrayData_0_valid_1[6:0];
  assign _zz_outputStreamArrayData_0_payload_3 = _zz_outputStreamArrayData_0_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l240_3);
  assign _zz_when_ArraySlice_l240_1 = _zz_when_ArraySlice_l240_2[6:0];
  assign _zz_when_ArraySlice_l240_4 = 4'b0000;
  assign _zz_when_ArraySlice_l240_3 = {4'd0, _zz_when_ArraySlice_l240_4};
  assign _zz_when_ArraySlice_l241_1 = (_zz_when_ArraySlice_l241_2 - 8'h01);
  assign _zz_when_ArraySlice_l241 = {5'd0, _zz_when_ArraySlice_l241_1};
  assign _zz_when_ArraySlice_l241_2 = (bReg * aReg);
  assign _zz_selectReadFifo_0_16 = (selectReadFifo_0 - _zz_selectReadFifo_0_17);
  assign _zz_selectReadFifo_0_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244 = (_zz_when_ArraySlice_l244_1 % aReg);
  assign _zz_when_ArraySlice_l244_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l249_3);
  assign _zz_when_ArraySlice_l249_1 = _zz_when_ArraySlice_l249_2[6:0];
  assign _zz_when_ArraySlice_l249_4 = 4'b0000;
  assign _zz_when_ArraySlice_l249_3 = {4'd0, _zz_when_ArraySlice_l249_4};
  assign _zz_when_ArraySlice_l250_1 = (_zz_when_ArraySlice_l250_2 - 8'h01);
  assign _zz_when_ArraySlice_l250 = {5'd0, _zz_when_ArraySlice_l250_1};
  assign _zz_when_ArraySlice_l250_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_24 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_24_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_24_1 = (_zz_realValue1_0_24_2 + _zz_realValue1_0_24_3);
  assign _zz_realValue1_0_24_2 = {1'd0, hReg};
  assign _zz_realValue1_0_24_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l252 = {1'd0, _zz_when_ArraySlice_l252_1};
  assign _zz_when_ArraySlice_l252_2 = (realValue1_0_24 / aReg);
  assign _zz_selectReadFifo_0_18 = (selectReadFifo_0 - _zz_selectReadFifo_0_19);
  assign _zz_selectReadFifo_0_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_0_21 = 1'b1;
  assign _zz_selectReadFifo_0_20 = {7'd0, _zz_selectReadFifo_0_21};
  assign _zz_when_ArraySlice_l158_208 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_208_1);
  assign _zz_when_ArraySlice_l158_208_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_208_1 = {4'd0, _zz_when_ArraySlice_l158_208_2};
  assign _zz_when_ArraySlice_l158_208_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_208 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_208_1 = (_zz_when_ArraySlice_l159_208_2 - _zz_when_ArraySlice_l159_208_3);
  assign _zz_when_ArraySlice_l159_208_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_208_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_208_4);
  assign _zz_when_ArraySlice_l159_208_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_208_4 = {4'd0, _zz_when_ArraySlice_l159_208_5};
  assign _zz__zz_realValue_0_208 = {1'd0, wReg};
  assign _zz__zz_realValue_0_208_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_208_1 = (_zz_realValue_0_208_2 + _zz_realValue_0_208_3);
  assign _zz_realValue_0_208_2 = {1'd0, wReg};
  assign _zz_realValue_0_208_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_208 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_208_1 = (_zz_when_ArraySlice_l166_208_2 + _zz_when_ArraySlice_l166_208_6);
  assign _zz_when_ArraySlice_l166_208_2 = (realValue_0_208 - _zz_when_ArraySlice_l166_208_3);
  assign _zz_when_ArraySlice_l166_208_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_208_4);
  assign _zz_when_ArraySlice_l166_208_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_208_4 = {4'd0, _zz_when_ArraySlice_l166_208_5};
  assign _zz_when_ArraySlice_l166_208_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_209 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_209_1);
  assign _zz_when_ArraySlice_l158_209_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_209_1 = {3'd0, _zz_when_ArraySlice_l158_209_2};
  assign _zz_when_ArraySlice_l158_209_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_209_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_209 = {1'd0, _zz_when_ArraySlice_l159_209_1};
  assign _zz_when_ArraySlice_l159_209_2 = (_zz_when_ArraySlice_l159_209_3 - _zz_when_ArraySlice_l159_209_4);
  assign _zz_when_ArraySlice_l159_209_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_209_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_209_5);
  assign _zz_when_ArraySlice_l159_209_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_209_5 = {3'd0, _zz_when_ArraySlice_l159_209_6};
  assign _zz__zz_realValue_0_209 = {1'd0, wReg};
  assign _zz__zz_realValue_0_209_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_209_1 = (_zz_realValue_0_209_2 + _zz_realValue_0_209_3);
  assign _zz_realValue_0_209_2 = {1'd0, wReg};
  assign _zz_realValue_0_209_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_209_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_209 = {1'd0, _zz_when_ArraySlice_l166_209_1};
  assign _zz_when_ArraySlice_l166_209_2 = (_zz_when_ArraySlice_l166_209_3 + _zz_when_ArraySlice_l166_209_7);
  assign _zz_when_ArraySlice_l166_209_3 = (realValue_0_209 - _zz_when_ArraySlice_l166_209_4);
  assign _zz_when_ArraySlice_l166_209_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_209_5);
  assign _zz_when_ArraySlice_l166_209_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_209_5 = {3'd0, _zz_when_ArraySlice_l166_209_6};
  assign _zz_when_ArraySlice_l166_209_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_210 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_210_1);
  assign _zz_when_ArraySlice_l158_210_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_210_1 = {2'd0, _zz_when_ArraySlice_l158_210_2};
  assign _zz_when_ArraySlice_l158_210_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_210_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_210 = {1'd0, _zz_when_ArraySlice_l159_210_1};
  assign _zz_when_ArraySlice_l159_210_2 = (_zz_when_ArraySlice_l159_210_3 - _zz_when_ArraySlice_l159_210_4);
  assign _zz_when_ArraySlice_l159_210_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_210_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_210_5);
  assign _zz_when_ArraySlice_l159_210_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_210_5 = {2'd0, _zz_when_ArraySlice_l159_210_6};
  assign _zz__zz_realValue_0_210 = {1'd0, wReg};
  assign _zz__zz_realValue_0_210_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_210_1 = (_zz_realValue_0_210_2 + _zz_realValue_0_210_3);
  assign _zz_realValue_0_210_2 = {1'd0, wReg};
  assign _zz_realValue_0_210_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_210_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_210 = {1'd0, _zz_when_ArraySlice_l166_210_1};
  assign _zz_when_ArraySlice_l166_210_2 = (_zz_when_ArraySlice_l166_210_3 + _zz_when_ArraySlice_l166_210_7);
  assign _zz_when_ArraySlice_l166_210_3 = (realValue_0_210 - _zz_when_ArraySlice_l166_210_4);
  assign _zz_when_ArraySlice_l166_210_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_210_5);
  assign _zz_when_ArraySlice_l166_210_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_210_5 = {2'd0, _zz_when_ArraySlice_l166_210_6};
  assign _zz_when_ArraySlice_l166_210_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_211 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_211_1);
  assign _zz_when_ArraySlice_l158_211_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_211_1 = {2'd0, _zz_when_ArraySlice_l158_211_2};
  assign _zz_when_ArraySlice_l158_211_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_211_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_211 = {1'd0, _zz_when_ArraySlice_l159_211_1};
  assign _zz_when_ArraySlice_l159_211_2 = (_zz_when_ArraySlice_l159_211_3 - _zz_when_ArraySlice_l159_211_4);
  assign _zz_when_ArraySlice_l159_211_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_211_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_211_5);
  assign _zz_when_ArraySlice_l159_211_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_211_5 = {2'd0, _zz_when_ArraySlice_l159_211_6};
  assign _zz__zz_realValue_0_211 = {1'd0, wReg};
  assign _zz__zz_realValue_0_211_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_211_1 = (_zz_realValue_0_211_2 + _zz_realValue_0_211_3);
  assign _zz_realValue_0_211_2 = {1'd0, wReg};
  assign _zz_realValue_0_211_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_211_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_211 = {1'd0, _zz_when_ArraySlice_l166_211_1};
  assign _zz_when_ArraySlice_l166_211_2 = (_zz_when_ArraySlice_l166_211_3 + _zz_when_ArraySlice_l166_211_7);
  assign _zz_when_ArraySlice_l166_211_3 = (realValue_0_211 - _zz_when_ArraySlice_l166_211_4);
  assign _zz_when_ArraySlice_l166_211_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_211_5);
  assign _zz_when_ArraySlice_l166_211_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_211_5 = {2'd0, _zz_when_ArraySlice_l166_211_6};
  assign _zz_when_ArraySlice_l166_211_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_212 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_212_1);
  assign _zz_when_ArraySlice_l158_212_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_212_1 = {1'd0, _zz_when_ArraySlice_l158_212_2};
  assign _zz_when_ArraySlice_l158_212_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_212_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_212 = {1'd0, _zz_when_ArraySlice_l159_212_1};
  assign _zz_when_ArraySlice_l159_212_2 = (_zz_when_ArraySlice_l159_212_3 - _zz_when_ArraySlice_l159_212_4);
  assign _zz_when_ArraySlice_l159_212_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_212_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_212_5);
  assign _zz_when_ArraySlice_l159_212_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_212_5 = {1'd0, _zz_when_ArraySlice_l159_212_6};
  assign _zz__zz_realValue_0_212 = {1'd0, wReg};
  assign _zz__zz_realValue_0_212_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_212_1 = (_zz_realValue_0_212_2 + _zz_realValue_0_212_3);
  assign _zz_realValue_0_212_2 = {1'd0, wReg};
  assign _zz_realValue_0_212_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_212_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_212 = {1'd0, _zz_when_ArraySlice_l166_212_1};
  assign _zz_when_ArraySlice_l166_212_2 = (_zz_when_ArraySlice_l166_212_3 + _zz_when_ArraySlice_l166_212_7);
  assign _zz_when_ArraySlice_l166_212_3 = (realValue_0_212 - _zz_when_ArraySlice_l166_212_4);
  assign _zz_when_ArraySlice_l166_212_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_212_5);
  assign _zz_when_ArraySlice_l166_212_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_212_5 = {1'd0, _zz_when_ArraySlice_l166_212_6};
  assign _zz_when_ArraySlice_l166_212_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_213 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_213_1);
  assign _zz_when_ArraySlice_l158_213_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_213_1 = {1'd0, _zz_when_ArraySlice_l158_213_2};
  assign _zz_when_ArraySlice_l158_213_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_213_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_213 = {2'd0, _zz_when_ArraySlice_l159_213_1};
  assign _zz_when_ArraySlice_l159_213_2 = (_zz_when_ArraySlice_l159_213_3 - _zz_when_ArraySlice_l159_213_4);
  assign _zz_when_ArraySlice_l159_213_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_213_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_213_5);
  assign _zz_when_ArraySlice_l159_213_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_213_5 = {1'd0, _zz_when_ArraySlice_l159_213_6};
  assign _zz__zz_realValue_0_213 = {1'd0, wReg};
  assign _zz__zz_realValue_0_213_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_213_1 = (_zz_realValue_0_213_2 + _zz_realValue_0_213_3);
  assign _zz_realValue_0_213_2 = {1'd0, wReg};
  assign _zz_realValue_0_213_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_213_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_213 = {2'd0, _zz_when_ArraySlice_l166_213_1};
  assign _zz_when_ArraySlice_l166_213_2 = (_zz_when_ArraySlice_l166_213_3 + _zz_when_ArraySlice_l166_213_7);
  assign _zz_when_ArraySlice_l166_213_3 = (realValue_0_213 - _zz_when_ArraySlice_l166_213_4);
  assign _zz_when_ArraySlice_l166_213_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_213_5);
  assign _zz_when_ArraySlice_l166_213_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_213_5 = {1'd0, _zz_when_ArraySlice_l166_213_6};
  assign _zz_when_ArraySlice_l166_213_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_214 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_214_1);
  assign _zz_when_ArraySlice_l158_214_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_214_1 = {1'd0, _zz_when_ArraySlice_l158_214_2};
  assign _zz_when_ArraySlice_l158_214_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_214_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_214 = {2'd0, _zz_when_ArraySlice_l159_214_1};
  assign _zz_when_ArraySlice_l159_214_2 = (_zz_when_ArraySlice_l159_214_3 - _zz_when_ArraySlice_l159_214_4);
  assign _zz_when_ArraySlice_l159_214_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_214_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_214_5);
  assign _zz_when_ArraySlice_l159_214_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_214_5 = {1'd0, _zz_when_ArraySlice_l159_214_6};
  assign _zz__zz_realValue_0_214 = {1'd0, wReg};
  assign _zz__zz_realValue_0_214_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_214_1 = (_zz_realValue_0_214_2 + _zz_realValue_0_214_3);
  assign _zz_realValue_0_214_2 = {1'd0, wReg};
  assign _zz_realValue_0_214_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_214_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_214 = {2'd0, _zz_when_ArraySlice_l166_214_1};
  assign _zz_when_ArraySlice_l166_214_2 = (_zz_when_ArraySlice_l166_214_3 + _zz_when_ArraySlice_l166_214_7);
  assign _zz_when_ArraySlice_l166_214_3 = (realValue_0_214 - _zz_when_ArraySlice_l166_214_4);
  assign _zz_when_ArraySlice_l166_214_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_214_5);
  assign _zz_when_ArraySlice_l166_214_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_214_5 = {1'd0, _zz_when_ArraySlice_l166_214_6};
  assign _zz_when_ArraySlice_l166_214_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_215 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_215_1);
  assign _zz_when_ArraySlice_l158_215_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_215_1 = {1'd0, _zz_when_ArraySlice_l158_215_2};
  assign _zz_when_ArraySlice_l158_215_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_215_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_215 = {3'd0, _zz_when_ArraySlice_l159_215_1};
  assign _zz_when_ArraySlice_l159_215_2 = (_zz_when_ArraySlice_l159_215_3 - _zz_when_ArraySlice_l159_215_4);
  assign _zz_when_ArraySlice_l159_215_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_215_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_215_5);
  assign _zz_when_ArraySlice_l159_215_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_215_5 = {1'd0, _zz_when_ArraySlice_l159_215_6};
  assign _zz__zz_realValue_0_215 = {1'd0, wReg};
  assign _zz__zz_realValue_0_215_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_215_1 = (_zz_realValue_0_215_2 + _zz_realValue_0_215_3);
  assign _zz_realValue_0_215_2 = {1'd0, wReg};
  assign _zz_realValue_0_215_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_215_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_215 = {3'd0, _zz_when_ArraySlice_l166_215_1};
  assign _zz_when_ArraySlice_l166_215_2 = (_zz_when_ArraySlice_l166_215_3 + _zz_when_ArraySlice_l166_215_7);
  assign _zz_when_ArraySlice_l166_215_3 = (realValue_0_215 - _zz_when_ArraySlice_l166_215_4);
  assign _zz_when_ArraySlice_l166_215_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_215_5);
  assign _zz_when_ArraySlice_l166_215_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_215_5 = {1'd0, _zz_when_ArraySlice_l166_215_6};
  assign _zz_when_ArraySlice_l166_215_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_1 = (_zz_when_ArraySlice_l260_2 + _zz_when_ArraySlice_l260_6);
  assign _zz_when_ArraySlice_l260_2 = (_zz_when_ArraySlice_l260_3 + 8'h01);
  assign _zz_when_ArraySlice_l260_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l260_4);
  assign _zz_when_ArraySlice_l260_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_4 = {1'd0, _zz_when_ArraySlice_l260_5};
  assign _zz_when_ArraySlice_l260_7 = 4'b0000;
  assign _zz_when_ArraySlice_l260_6 = {4'd0, _zz_when_ArraySlice_l260_7};
  assign _zz_when_ArraySlice_l263 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_1 = (_zz_when_ArraySlice_l263_2 + 8'h01);
  assign _zz_when_ArraySlice_l263_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l263_3);
  assign _zz_when_ArraySlice_l263_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_3 = {1'd0, _zz_when_ArraySlice_l263_4};
  assign _zz_selectReadFifo_0_22 = (selectReadFifo_0 + _zz_selectReadFifo_0_23);
  assign _zz_selectReadFifo_0_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_23 = {1'd0, _zz_selectReadFifo_0_24};
  assign _zz_when_ArraySlice_l270 = (_zz_when_ArraySlice_l270_1 % aReg);
  assign _zz_when_ArraySlice_l270_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l274_3);
  assign _zz_when_ArraySlice_l274_1 = _zz_when_ArraySlice_l274_2[6:0];
  assign _zz_when_ArraySlice_l274_4 = 4'b0000;
  assign _zz_when_ArraySlice_l274_3 = {4'd0, _zz_when_ArraySlice_l274_4};
  assign _zz_when_ArraySlice_l275_1 = (_zz_when_ArraySlice_l275_2 - _zz_when_ArraySlice_l275_3);
  assign _zz_when_ArraySlice_l275 = {5'd0, _zz_when_ArraySlice_l275_1};
  assign _zz_when_ArraySlice_l275_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_4 = 1'b1;
  assign _zz_when_ArraySlice_l275_3 = {7'd0, _zz_when_ArraySlice_l275_4};
  assign _zz__zz_realValue1_0_25 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_25_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_25_1 = (_zz_realValue1_0_25_2 + _zz_realValue1_0_25_3);
  assign _zz_realValue1_0_25_2 = {1'd0, hReg};
  assign _zz_realValue1_0_25_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l277 = {1'd0, _zz_when_ArraySlice_l277_1};
  assign _zz_when_ArraySlice_l277_2 = (realValue1_0_25 / aReg);
  assign _zz_selectReadFifo_0_25 = (selectReadFifo_0 - _zz_selectReadFifo_0_26);
  assign _zz_selectReadFifo_0_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_216 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_216_1);
  assign _zz_when_ArraySlice_l158_216_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_216_1 = {4'd0, _zz_when_ArraySlice_l158_216_2};
  assign _zz_when_ArraySlice_l158_216_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_216 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_216_1 = (_zz_when_ArraySlice_l159_216_2 - _zz_when_ArraySlice_l159_216_3);
  assign _zz_when_ArraySlice_l159_216_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_216_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_216_4);
  assign _zz_when_ArraySlice_l159_216_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_216_4 = {4'd0, _zz_when_ArraySlice_l159_216_5};
  assign _zz__zz_realValue_0_216 = {1'd0, wReg};
  assign _zz__zz_realValue_0_216_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_216_1 = (_zz_realValue_0_216_2 + _zz_realValue_0_216_3);
  assign _zz_realValue_0_216_2 = {1'd0, wReg};
  assign _zz_realValue_0_216_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_216 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_216_1 = (_zz_when_ArraySlice_l166_216_2 + _zz_when_ArraySlice_l166_216_6);
  assign _zz_when_ArraySlice_l166_216_2 = (realValue_0_216 - _zz_when_ArraySlice_l166_216_3);
  assign _zz_when_ArraySlice_l166_216_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_216_4);
  assign _zz_when_ArraySlice_l166_216_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_216_4 = {4'd0, _zz_when_ArraySlice_l166_216_5};
  assign _zz_when_ArraySlice_l166_216_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_217 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_217_1);
  assign _zz_when_ArraySlice_l158_217_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_217_1 = {3'd0, _zz_when_ArraySlice_l158_217_2};
  assign _zz_when_ArraySlice_l158_217_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_217_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_217 = {1'd0, _zz_when_ArraySlice_l159_217_1};
  assign _zz_when_ArraySlice_l159_217_2 = (_zz_when_ArraySlice_l159_217_3 - _zz_when_ArraySlice_l159_217_4);
  assign _zz_when_ArraySlice_l159_217_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_217_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_217_5);
  assign _zz_when_ArraySlice_l159_217_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_217_5 = {3'd0, _zz_when_ArraySlice_l159_217_6};
  assign _zz__zz_realValue_0_217 = {1'd0, wReg};
  assign _zz__zz_realValue_0_217_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_217_1 = (_zz_realValue_0_217_2 + _zz_realValue_0_217_3);
  assign _zz_realValue_0_217_2 = {1'd0, wReg};
  assign _zz_realValue_0_217_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_217_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_217 = {1'd0, _zz_when_ArraySlice_l166_217_1};
  assign _zz_when_ArraySlice_l166_217_2 = (_zz_when_ArraySlice_l166_217_3 + _zz_when_ArraySlice_l166_217_7);
  assign _zz_when_ArraySlice_l166_217_3 = (realValue_0_217 - _zz_when_ArraySlice_l166_217_4);
  assign _zz_when_ArraySlice_l166_217_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_217_5);
  assign _zz_when_ArraySlice_l166_217_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_217_5 = {3'd0, _zz_when_ArraySlice_l166_217_6};
  assign _zz_when_ArraySlice_l166_217_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_218 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_218_1);
  assign _zz_when_ArraySlice_l158_218_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_218_1 = {2'd0, _zz_when_ArraySlice_l158_218_2};
  assign _zz_when_ArraySlice_l158_218_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_218_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_218 = {1'd0, _zz_when_ArraySlice_l159_218_1};
  assign _zz_when_ArraySlice_l159_218_2 = (_zz_when_ArraySlice_l159_218_3 - _zz_when_ArraySlice_l159_218_4);
  assign _zz_when_ArraySlice_l159_218_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_218_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_218_5);
  assign _zz_when_ArraySlice_l159_218_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_218_5 = {2'd0, _zz_when_ArraySlice_l159_218_6};
  assign _zz__zz_realValue_0_218 = {1'd0, wReg};
  assign _zz__zz_realValue_0_218_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_218_1 = (_zz_realValue_0_218_2 + _zz_realValue_0_218_3);
  assign _zz_realValue_0_218_2 = {1'd0, wReg};
  assign _zz_realValue_0_218_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_218_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_218 = {1'd0, _zz_when_ArraySlice_l166_218_1};
  assign _zz_when_ArraySlice_l166_218_2 = (_zz_when_ArraySlice_l166_218_3 + _zz_when_ArraySlice_l166_218_7);
  assign _zz_when_ArraySlice_l166_218_3 = (realValue_0_218 - _zz_when_ArraySlice_l166_218_4);
  assign _zz_when_ArraySlice_l166_218_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_218_5);
  assign _zz_when_ArraySlice_l166_218_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_218_5 = {2'd0, _zz_when_ArraySlice_l166_218_6};
  assign _zz_when_ArraySlice_l166_218_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_219 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_219_1);
  assign _zz_when_ArraySlice_l158_219_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_219_1 = {2'd0, _zz_when_ArraySlice_l158_219_2};
  assign _zz_when_ArraySlice_l158_219_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_219_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_219 = {1'd0, _zz_when_ArraySlice_l159_219_1};
  assign _zz_when_ArraySlice_l159_219_2 = (_zz_when_ArraySlice_l159_219_3 - _zz_when_ArraySlice_l159_219_4);
  assign _zz_when_ArraySlice_l159_219_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_219_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_219_5);
  assign _zz_when_ArraySlice_l159_219_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_219_5 = {2'd0, _zz_when_ArraySlice_l159_219_6};
  assign _zz__zz_realValue_0_219 = {1'd0, wReg};
  assign _zz__zz_realValue_0_219_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_219_1 = (_zz_realValue_0_219_2 + _zz_realValue_0_219_3);
  assign _zz_realValue_0_219_2 = {1'd0, wReg};
  assign _zz_realValue_0_219_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_219_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_219 = {1'd0, _zz_when_ArraySlice_l166_219_1};
  assign _zz_when_ArraySlice_l166_219_2 = (_zz_when_ArraySlice_l166_219_3 + _zz_when_ArraySlice_l166_219_7);
  assign _zz_when_ArraySlice_l166_219_3 = (realValue_0_219 - _zz_when_ArraySlice_l166_219_4);
  assign _zz_when_ArraySlice_l166_219_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_219_5);
  assign _zz_when_ArraySlice_l166_219_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_219_5 = {2'd0, _zz_when_ArraySlice_l166_219_6};
  assign _zz_when_ArraySlice_l166_219_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_220 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_220_1);
  assign _zz_when_ArraySlice_l158_220_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_220_1 = {1'd0, _zz_when_ArraySlice_l158_220_2};
  assign _zz_when_ArraySlice_l158_220_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_220_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_220 = {1'd0, _zz_when_ArraySlice_l159_220_1};
  assign _zz_when_ArraySlice_l159_220_2 = (_zz_when_ArraySlice_l159_220_3 - _zz_when_ArraySlice_l159_220_4);
  assign _zz_when_ArraySlice_l159_220_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_220_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_220_5);
  assign _zz_when_ArraySlice_l159_220_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_220_5 = {1'd0, _zz_when_ArraySlice_l159_220_6};
  assign _zz__zz_realValue_0_220 = {1'd0, wReg};
  assign _zz__zz_realValue_0_220_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_220_1 = (_zz_realValue_0_220_2 + _zz_realValue_0_220_3);
  assign _zz_realValue_0_220_2 = {1'd0, wReg};
  assign _zz_realValue_0_220_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_220_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_220 = {1'd0, _zz_when_ArraySlice_l166_220_1};
  assign _zz_when_ArraySlice_l166_220_2 = (_zz_when_ArraySlice_l166_220_3 + _zz_when_ArraySlice_l166_220_7);
  assign _zz_when_ArraySlice_l166_220_3 = (realValue_0_220 - _zz_when_ArraySlice_l166_220_4);
  assign _zz_when_ArraySlice_l166_220_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_220_5);
  assign _zz_when_ArraySlice_l166_220_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_220_5 = {1'd0, _zz_when_ArraySlice_l166_220_6};
  assign _zz_when_ArraySlice_l166_220_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_221 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_221_1);
  assign _zz_when_ArraySlice_l158_221_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_221_1 = {1'd0, _zz_when_ArraySlice_l158_221_2};
  assign _zz_when_ArraySlice_l158_221_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_221_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_221 = {2'd0, _zz_when_ArraySlice_l159_221_1};
  assign _zz_when_ArraySlice_l159_221_2 = (_zz_when_ArraySlice_l159_221_3 - _zz_when_ArraySlice_l159_221_4);
  assign _zz_when_ArraySlice_l159_221_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_221_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_221_5);
  assign _zz_when_ArraySlice_l159_221_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_221_5 = {1'd0, _zz_when_ArraySlice_l159_221_6};
  assign _zz__zz_realValue_0_221 = {1'd0, wReg};
  assign _zz__zz_realValue_0_221_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_221_1 = (_zz_realValue_0_221_2 + _zz_realValue_0_221_3);
  assign _zz_realValue_0_221_2 = {1'd0, wReg};
  assign _zz_realValue_0_221_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_221_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_221 = {2'd0, _zz_when_ArraySlice_l166_221_1};
  assign _zz_when_ArraySlice_l166_221_2 = (_zz_when_ArraySlice_l166_221_3 + _zz_when_ArraySlice_l166_221_7);
  assign _zz_when_ArraySlice_l166_221_3 = (realValue_0_221 - _zz_when_ArraySlice_l166_221_4);
  assign _zz_when_ArraySlice_l166_221_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_221_5);
  assign _zz_when_ArraySlice_l166_221_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_221_5 = {1'd0, _zz_when_ArraySlice_l166_221_6};
  assign _zz_when_ArraySlice_l166_221_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_222 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_222_1);
  assign _zz_when_ArraySlice_l158_222_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_222_1 = {1'd0, _zz_when_ArraySlice_l158_222_2};
  assign _zz_when_ArraySlice_l158_222_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_222_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_222 = {2'd0, _zz_when_ArraySlice_l159_222_1};
  assign _zz_when_ArraySlice_l159_222_2 = (_zz_when_ArraySlice_l159_222_3 - _zz_when_ArraySlice_l159_222_4);
  assign _zz_when_ArraySlice_l159_222_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_222_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_222_5);
  assign _zz_when_ArraySlice_l159_222_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_222_5 = {1'd0, _zz_when_ArraySlice_l159_222_6};
  assign _zz__zz_realValue_0_222 = {1'd0, wReg};
  assign _zz__zz_realValue_0_222_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_222_1 = (_zz_realValue_0_222_2 + _zz_realValue_0_222_3);
  assign _zz_realValue_0_222_2 = {1'd0, wReg};
  assign _zz_realValue_0_222_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_222_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_222 = {2'd0, _zz_when_ArraySlice_l166_222_1};
  assign _zz_when_ArraySlice_l166_222_2 = (_zz_when_ArraySlice_l166_222_3 + _zz_when_ArraySlice_l166_222_7);
  assign _zz_when_ArraySlice_l166_222_3 = (realValue_0_222 - _zz_when_ArraySlice_l166_222_4);
  assign _zz_when_ArraySlice_l166_222_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_222_5);
  assign _zz_when_ArraySlice_l166_222_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_222_5 = {1'd0, _zz_when_ArraySlice_l166_222_6};
  assign _zz_when_ArraySlice_l166_222_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_223 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_223_1);
  assign _zz_when_ArraySlice_l158_223_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_223_1 = {1'd0, _zz_when_ArraySlice_l158_223_2};
  assign _zz_when_ArraySlice_l158_223_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_223_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_223 = {3'd0, _zz_when_ArraySlice_l159_223_1};
  assign _zz_when_ArraySlice_l159_223_2 = (_zz_when_ArraySlice_l159_223_3 - _zz_when_ArraySlice_l159_223_4);
  assign _zz_when_ArraySlice_l159_223_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_223_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_223_5);
  assign _zz_when_ArraySlice_l159_223_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_223_5 = {1'd0, _zz_when_ArraySlice_l159_223_6};
  assign _zz__zz_realValue_0_223 = {1'd0, wReg};
  assign _zz__zz_realValue_0_223_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_223_1 = (_zz_realValue_0_223_2 + _zz_realValue_0_223_3);
  assign _zz_realValue_0_223_2 = {1'd0, wReg};
  assign _zz_realValue_0_223_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_223_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_223 = {3'd0, _zz_when_ArraySlice_l166_223_1};
  assign _zz_when_ArraySlice_l166_223_2 = (_zz_when_ArraySlice_l166_223_3 + _zz_when_ArraySlice_l166_223_7);
  assign _zz_when_ArraySlice_l166_223_3 = (realValue_0_223 - _zz_when_ArraySlice_l166_223_4);
  assign _zz_when_ArraySlice_l166_223_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_223_5);
  assign _zz_when_ArraySlice_l166_223_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_223_5 = {1'd0, _zz_when_ArraySlice_l166_223_6};
  assign _zz_when_ArraySlice_l166_223_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_1 = (_zz_when_ArraySlice_l285_2 + _zz_when_ArraySlice_l285_6);
  assign _zz_when_ArraySlice_l285_2 = (_zz_when_ArraySlice_l285_3 + 8'h01);
  assign _zz_when_ArraySlice_l285_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l285_4);
  assign _zz_when_ArraySlice_l285_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_4 = {1'd0, _zz_when_ArraySlice_l285_5};
  assign _zz_when_ArraySlice_l285_7 = 4'b0000;
  assign _zz_when_ArraySlice_l285_6 = {4'd0, _zz_when_ArraySlice_l285_7};
  assign _zz_when_ArraySlice_l288 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_1 = (_zz_when_ArraySlice_l288_2 + 8'h01);
  assign _zz_when_ArraySlice_l288_2 = (selectReadFifo_0 + _zz_when_ArraySlice_l288_3);
  assign _zz_when_ArraySlice_l288_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_3 = {1'd0, _zz_when_ArraySlice_l288_4};
  assign _zz_selectReadFifo_0_27 = (selectReadFifo_0 + _zz_selectReadFifo_0_28);
  assign _zz_selectReadFifo_0_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_0_28 = {1'd0, _zz_selectReadFifo_0_29};
  assign _zz_when_ArraySlice_l295 = (_zz_when_ArraySlice_l295_1 % aReg);
  assign _zz_when_ArraySlice_l295_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_1 = (_zz_when_ArraySlice_l306_2 - 8'h01);
  assign _zz_when_ArraySlice_l306 = {5'd0, _zz_when_ArraySlice_l306_1};
  assign _zz_when_ArraySlice_l306_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_26 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_26_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_26_1 = (_zz_realValue1_0_26_2 + _zz_realValue1_0_26_3);
  assign _zz_realValue1_0_26_2 = {1'd0, hReg};
  assign _zz_realValue1_0_26_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_1 = (outSliceNumb_0_value + 7'h01);
  assign _zz_when_ArraySlice_l307 = {1'd0, _zz_when_ArraySlice_l307_1};
  assign _zz_when_ArraySlice_l307_2 = (realValue1_0_26 / aReg);
  assign _zz_selectReadFifo_0_30 = (selectReadFifo_0 - _zz_selectReadFifo_0_31);
  assign _zz_selectReadFifo_0_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_224 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_224_1);
  assign _zz_when_ArraySlice_l158_224_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_224_1 = {4'd0, _zz_when_ArraySlice_l158_224_2};
  assign _zz_when_ArraySlice_l158_224_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_224 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_224_1 = (_zz_when_ArraySlice_l159_224_2 - _zz_when_ArraySlice_l159_224_3);
  assign _zz_when_ArraySlice_l159_224_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_224_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_224_4);
  assign _zz_when_ArraySlice_l159_224_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_224_4 = {4'd0, _zz_when_ArraySlice_l159_224_5};
  assign _zz__zz_realValue_0_224 = {1'd0, wReg};
  assign _zz__zz_realValue_0_224_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_224_1 = (_zz_realValue_0_224_2 + _zz_realValue_0_224_3);
  assign _zz_realValue_0_224_2 = {1'd0, wReg};
  assign _zz_realValue_0_224_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_224 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_224_1 = (_zz_when_ArraySlice_l166_224_2 + _zz_when_ArraySlice_l166_224_6);
  assign _zz_when_ArraySlice_l166_224_2 = (realValue_0_224 - _zz_when_ArraySlice_l166_224_3);
  assign _zz_when_ArraySlice_l166_224_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_224_4);
  assign _zz_when_ArraySlice_l166_224_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_224_4 = {4'd0, _zz_when_ArraySlice_l166_224_5};
  assign _zz_when_ArraySlice_l166_224_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_225 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_225_1);
  assign _zz_when_ArraySlice_l158_225_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_225_1 = {3'd0, _zz_when_ArraySlice_l158_225_2};
  assign _zz_when_ArraySlice_l158_225_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_225_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_225 = {1'd0, _zz_when_ArraySlice_l159_225_1};
  assign _zz_when_ArraySlice_l159_225_2 = (_zz_when_ArraySlice_l159_225_3 - _zz_when_ArraySlice_l159_225_4);
  assign _zz_when_ArraySlice_l159_225_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_225_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_225_5);
  assign _zz_when_ArraySlice_l159_225_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_225_5 = {3'd0, _zz_when_ArraySlice_l159_225_6};
  assign _zz__zz_realValue_0_225 = {1'd0, wReg};
  assign _zz__zz_realValue_0_225_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_225_1 = (_zz_realValue_0_225_2 + _zz_realValue_0_225_3);
  assign _zz_realValue_0_225_2 = {1'd0, wReg};
  assign _zz_realValue_0_225_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_225_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_225 = {1'd0, _zz_when_ArraySlice_l166_225_1};
  assign _zz_when_ArraySlice_l166_225_2 = (_zz_when_ArraySlice_l166_225_3 + _zz_when_ArraySlice_l166_225_7);
  assign _zz_when_ArraySlice_l166_225_3 = (realValue_0_225 - _zz_when_ArraySlice_l166_225_4);
  assign _zz_when_ArraySlice_l166_225_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_225_5);
  assign _zz_when_ArraySlice_l166_225_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_225_5 = {3'd0, _zz_when_ArraySlice_l166_225_6};
  assign _zz_when_ArraySlice_l166_225_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_226 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_226_1);
  assign _zz_when_ArraySlice_l158_226_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_226_1 = {2'd0, _zz_when_ArraySlice_l158_226_2};
  assign _zz_when_ArraySlice_l158_226_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_226_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_226 = {1'd0, _zz_when_ArraySlice_l159_226_1};
  assign _zz_when_ArraySlice_l159_226_2 = (_zz_when_ArraySlice_l159_226_3 - _zz_when_ArraySlice_l159_226_4);
  assign _zz_when_ArraySlice_l159_226_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_226_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_226_5);
  assign _zz_when_ArraySlice_l159_226_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_226_5 = {2'd0, _zz_when_ArraySlice_l159_226_6};
  assign _zz__zz_realValue_0_226 = {1'd0, wReg};
  assign _zz__zz_realValue_0_226_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_226_1 = (_zz_realValue_0_226_2 + _zz_realValue_0_226_3);
  assign _zz_realValue_0_226_2 = {1'd0, wReg};
  assign _zz_realValue_0_226_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_226_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_226 = {1'd0, _zz_when_ArraySlice_l166_226_1};
  assign _zz_when_ArraySlice_l166_226_2 = (_zz_when_ArraySlice_l166_226_3 + _zz_when_ArraySlice_l166_226_7);
  assign _zz_when_ArraySlice_l166_226_3 = (realValue_0_226 - _zz_when_ArraySlice_l166_226_4);
  assign _zz_when_ArraySlice_l166_226_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_226_5);
  assign _zz_when_ArraySlice_l166_226_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_226_5 = {2'd0, _zz_when_ArraySlice_l166_226_6};
  assign _zz_when_ArraySlice_l166_226_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_227 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_227_1);
  assign _zz_when_ArraySlice_l158_227_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_227_1 = {2'd0, _zz_when_ArraySlice_l158_227_2};
  assign _zz_when_ArraySlice_l158_227_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_227_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_227 = {1'd0, _zz_when_ArraySlice_l159_227_1};
  assign _zz_when_ArraySlice_l159_227_2 = (_zz_when_ArraySlice_l159_227_3 - _zz_when_ArraySlice_l159_227_4);
  assign _zz_when_ArraySlice_l159_227_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_227_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_227_5);
  assign _zz_when_ArraySlice_l159_227_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_227_5 = {2'd0, _zz_when_ArraySlice_l159_227_6};
  assign _zz__zz_realValue_0_227 = {1'd0, wReg};
  assign _zz__zz_realValue_0_227_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_227_1 = (_zz_realValue_0_227_2 + _zz_realValue_0_227_3);
  assign _zz_realValue_0_227_2 = {1'd0, wReg};
  assign _zz_realValue_0_227_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_227_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_227 = {1'd0, _zz_when_ArraySlice_l166_227_1};
  assign _zz_when_ArraySlice_l166_227_2 = (_zz_when_ArraySlice_l166_227_3 + _zz_when_ArraySlice_l166_227_7);
  assign _zz_when_ArraySlice_l166_227_3 = (realValue_0_227 - _zz_when_ArraySlice_l166_227_4);
  assign _zz_when_ArraySlice_l166_227_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_227_5);
  assign _zz_when_ArraySlice_l166_227_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_227_5 = {2'd0, _zz_when_ArraySlice_l166_227_6};
  assign _zz_when_ArraySlice_l166_227_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_228 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_228_1);
  assign _zz_when_ArraySlice_l158_228_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_228_1 = {1'd0, _zz_when_ArraySlice_l158_228_2};
  assign _zz_when_ArraySlice_l158_228_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_228_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_228 = {1'd0, _zz_when_ArraySlice_l159_228_1};
  assign _zz_when_ArraySlice_l159_228_2 = (_zz_when_ArraySlice_l159_228_3 - _zz_when_ArraySlice_l159_228_4);
  assign _zz_when_ArraySlice_l159_228_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_228_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_228_5);
  assign _zz_when_ArraySlice_l159_228_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_228_5 = {1'd0, _zz_when_ArraySlice_l159_228_6};
  assign _zz__zz_realValue_0_228 = {1'd0, wReg};
  assign _zz__zz_realValue_0_228_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_228_1 = (_zz_realValue_0_228_2 + _zz_realValue_0_228_3);
  assign _zz_realValue_0_228_2 = {1'd0, wReg};
  assign _zz_realValue_0_228_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_228_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_228 = {1'd0, _zz_when_ArraySlice_l166_228_1};
  assign _zz_when_ArraySlice_l166_228_2 = (_zz_when_ArraySlice_l166_228_3 + _zz_when_ArraySlice_l166_228_7);
  assign _zz_when_ArraySlice_l166_228_3 = (realValue_0_228 - _zz_when_ArraySlice_l166_228_4);
  assign _zz_when_ArraySlice_l166_228_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_228_5);
  assign _zz_when_ArraySlice_l166_228_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_228_5 = {1'd0, _zz_when_ArraySlice_l166_228_6};
  assign _zz_when_ArraySlice_l166_228_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_229 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_229_1);
  assign _zz_when_ArraySlice_l158_229_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_229_1 = {1'd0, _zz_when_ArraySlice_l158_229_2};
  assign _zz_when_ArraySlice_l158_229_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_229_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_229 = {2'd0, _zz_when_ArraySlice_l159_229_1};
  assign _zz_when_ArraySlice_l159_229_2 = (_zz_when_ArraySlice_l159_229_3 - _zz_when_ArraySlice_l159_229_4);
  assign _zz_when_ArraySlice_l159_229_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_229_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_229_5);
  assign _zz_when_ArraySlice_l159_229_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_229_5 = {1'd0, _zz_when_ArraySlice_l159_229_6};
  assign _zz__zz_realValue_0_229 = {1'd0, wReg};
  assign _zz__zz_realValue_0_229_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_229_1 = (_zz_realValue_0_229_2 + _zz_realValue_0_229_3);
  assign _zz_realValue_0_229_2 = {1'd0, wReg};
  assign _zz_realValue_0_229_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_229_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_229 = {2'd0, _zz_when_ArraySlice_l166_229_1};
  assign _zz_when_ArraySlice_l166_229_2 = (_zz_when_ArraySlice_l166_229_3 + _zz_when_ArraySlice_l166_229_7);
  assign _zz_when_ArraySlice_l166_229_3 = (realValue_0_229 - _zz_when_ArraySlice_l166_229_4);
  assign _zz_when_ArraySlice_l166_229_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_229_5);
  assign _zz_when_ArraySlice_l166_229_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_229_5 = {1'd0, _zz_when_ArraySlice_l166_229_6};
  assign _zz_when_ArraySlice_l166_229_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_230 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_230_1);
  assign _zz_when_ArraySlice_l158_230_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_230_1 = {1'd0, _zz_when_ArraySlice_l158_230_2};
  assign _zz_when_ArraySlice_l158_230_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_230_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_230 = {2'd0, _zz_when_ArraySlice_l159_230_1};
  assign _zz_when_ArraySlice_l159_230_2 = (_zz_when_ArraySlice_l159_230_3 - _zz_when_ArraySlice_l159_230_4);
  assign _zz_when_ArraySlice_l159_230_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_230_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_230_5);
  assign _zz_when_ArraySlice_l159_230_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_230_5 = {1'd0, _zz_when_ArraySlice_l159_230_6};
  assign _zz__zz_realValue_0_230 = {1'd0, wReg};
  assign _zz__zz_realValue_0_230_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_230_1 = (_zz_realValue_0_230_2 + _zz_realValue_0_230_3);
  assign _zz_realValue_0_230_2 = {1'd0, wReg};
  assign _zz_realValue_0_230_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_230_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_230 = {2'd0, _zz_when_ArraySlice_l166_230_1};
  assign _zz_when_ArraySlice_l166_230_2 = (_zz_when_ArraySlice_l166_230_3 + _zz_when_ArraySlice_l166_230_7);
  assign _zz_when_ArraySlice_l166_230_3 = (realValue_0_230 - _zz_when_ArraySlice_l166_230_4);
  assign _zz_when_ArraySlice_l166_230_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_230_5);
  assign _zz_when_ArraySlice_l166_230_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_230_5 = {1'd0, _zz_when_ArraySlice_l166_230_6};
  assign _zz_when_ArraySlice_l166_230_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_231 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_231_1);
  assign _zz_when_ArraySlice_l158_231_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_231_1 = {1'd0, _zz_when_ArraySlice_l158_231_2};
  assign _zz_when_ArraySlice_l158_231_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_231_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_231 = {3'd0, _zz_when_ArraySlice_l159_231_1};
  assign _zz_when_ArraySlice_l159_231_2 = (_zz_when_ArraySlice_l159_231_3 - _zz_when_ArraySlice_l159_231_4);
  assign _zz_when_ArraySlice_l159_231_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_231_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_231_5);
  assign _zz_when_ArraySlice_l159_231_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_231_5 = {1'd0, _zz_when_ArraySlice_l159_231_6};
  assign _zz__zz_realValue_0_231 = {1'd0, wReg};
  assign _zz__zz_realValue_0_231_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_231_1 = (_zz_realValue_0_231_2 + _zz_realValue_0_231_3);
  assign _zz_realValue_0_231_2 = {1'd0, wReg};
  assign _zz_realValue_0_231_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_231_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_231 = {3'd0, _zz_when_ArraySlice_l166_231_1};
  assign _zz_when_ArraySlice_l166_231_2 = (_zz_when_ArraySlice_l166_231_3 + _zz_when_ArraySlice_l166_231_7);
  assign _zz_when_ArraySlice_l166_231_3 = (realValue_0_231 - _zz_when_ArraySlice_l166_231_4);
  assign _zz_when_ArraySlice_l166_231_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_231_5);
  assign _zz_when_ArraySlice_l166_231_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_231_5 = {1'd0, _zz_when_ArraySlice_l166_231_6};
  assign _zz_when_ArraySlice_l166_231_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318 = (_zz_when_ArraySlice_l318_1 % aReg);
  assign _zz_when_ArraySlice_l318_1 = (handshakeTimes_0_value + 13'h0001);
  assign _zz_when_ArraySlice_l304 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_1 = (selectReadFifo_0 + _zz_when_ArraySlice_l304_2);
  assign _zz_when_ArraySlice_l304_3 = 4'b0000;
  assign _zz_when_ArraySlice_l304_2 = {4'd0, _zz_when_ArraySlice_l304_3};
  assign _zz_when_ArraySlice_l325_1 = (_zz_when_ArraySlice_l325_2 - 8'h01);
  assign _zz_when_ArraySlice_l325 = {5'd0, _zz_when_ArraySlice_l325_1};
  assign _zz_when_ArraySlice_l325_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_1_1 = (selectReadFifo_1 + _zz_when_ArraySlice_l233_1_2);
  assign _zz_when_ArraySlice_l233_1_3 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l233_1_2 = {3'd0, _zz_when_ArraySlice_l233_1_3};
  assign _zz_when_ArraySlice_l233_1_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l234_1_4);
  assign _zz_when_ArraySlice_l234_1_2 = _zz_when_ArraySlice_l234_1_3[6:0];
  assign _zz_when_ArraySlice_l234_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l234_1_4 = {3'd0, _zz_when_ArraySlice_l234_1_5};
  assign _zz__zz_outputStreamArrayData_1_valid_1_2 = (bReg * 1'b1);
  assign _zz__zz_outputStreamArrayData_1_valid_1_1 = {3'd0, _zz__zz_outputStreamArrayData_1_valid_1_2};
  assign _zz__zz_12 = _zz_outputStreamArrayData_1_valid_1[6:0];
  assign _zz_outputStreamArrayData_1_valid_5 = _zz_outputStreamArrayData_1_valid_1[6:0];
  assign _zz_outputStreamArrayData_1_payload_3 = _zz_outputStreamArrayData_1_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l240_1_4);
  assign _zz_when_ArraySlice_l240_1_2 = _zz_when_ArraySlice_l240_1_3[6:0];
  assign _zz_when_ArraySlice_l240_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l240_1_4 = {3'd0, _zz_when_ArraySlice_l240_1_5};
  assign _zz_when_ArraySlice_l241_1_2 = (_zz_when_ArraySlice_l241_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l241_1_1 = {5'd0, _zz_when_ArraySlice_l241_1_2};
  assign _zz_when_ArraySlice_l241_1_3 = (bReg * aReg);
  assign _zz_selectReadFifo_1_16 = (selectReadFifo_1 - _zz_selectReadFifo_1_17);
  assign _zz_selectReadFifo_1_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_1_1 = (_zz_when_ArraySlice_l244_1_2 % aReg);
  assign _zz_when_ArraySlice_l244_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l249_1_4);
  assign _zz_when_ArraySlice_l249_1_2 = _zz_when_ArraySlice_l249_1_3[6:0];
  assign _zz_when_ArraySlice_l249_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l249_1_4 = {3'd0, _zz_when_ArraySlice_l249_1_5};
  assign _zz_when_ArraySlice_l250_1_2 = (_zz_when_ArraySlice_l250_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l250_1_1 = {5'd0, _zz_when_ArraySlice_l250_1_2};
  assign _zz_when_ArraySlice_l250_1_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_27 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_27_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_27_1 = (_zz_realValue1_0_27_2 + _zz_realValue1_0_27_3);
  assign _zz_realValue1_0_27_2 = {1'd0, hReg};
  assign _zz_realValue1_0_27_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l252_1_1 = {1'd0, _zz_when_ArraySlice_l252_1_2};
  assign _zz_when_ArraySlice_l252_1_3 = (realValue1_0_27 / aReg);
  assign _zz_selectReadFifo_1_18 = (selectReadFifo_1 - _zz_selectReadFifo_1_19);
  assign _zz_selectReadFifo_1_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_1_21 = 1'b1;
  assign _zz_selectReadFifo_1_20 = {7'd0, _zz_selectReadFifo_1_21};
  assign _zz_when_ArraySlice_l158_232 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_232_1);
  assign _zz_when_ArraySlice_l158_232_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_232_1 = {4'd0, _zz_when_ArraySlice_l158_232_2};
  assign _zz_when_ArraySlice_l158_232_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_232 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_232_1 = (_zz_when_ArraySlice_l159_232_2 - _zz_when_ArraySlice_l159_232_3);
  assign _zz_when_ArraySlice_l159_232_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_232_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_232_4);
  assign _zz_when_ArraySlice_l159_232_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_232_4 = {4'd0, _zz_when_ArraySlice_l159_232_5};
  assign _zz__zz_realValue_0_232 = {1'd0, wReg};
  assign _zz__zz_realValue_0_232_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_232_1 = (_zz_realValue_0_232_2 + _zz_realValue_0_232_3);
  assign _zz_realValue_0_232_2 = {1'd0, wReg};
  assign _zz_realValue_0_232_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_232 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_232_1 = (_zz_when_ArraySlice_l166_232_2 + _zz_when_ArraySlice_l166_232_6);
  assign _zz_when_ArraySlice_l166_232_2 = (realValue_0_232 - _zz_when_ArraySlice_l166_232_3);
  assign _zz_when_ArraySlice_l166_232_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_232_4);
  assign _zz_when_ArraySlice_l166_232_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_232_4 = {4'd0, _zz_when_ArraySlice_l166_232_5};
  assign _zz_when_ArraySlice_l166_232_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_233 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_233_1);
  assign _zz_when_ArraySlice_l158_233_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_233_1 = {3'd0, _zz_when_ArraySlice_l158_233_2};
  assign _zz_when_ArraySlice_l158_233_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_233_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_233 = {1'd0, _zz_when_ArraySlice_l159_233_1};
  assign _zz_when_ArraySlice_l159_233_2 = (_zz_when_ArraySlice_l159_233_3 - _zz_when_ArraySlice_l159_233_4);
  assign _zz_when_ArraySlice_l159_233_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_233_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_233_5);
  assign _zz_when_ArraySlice_l159_233_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_233_5 = {3'd0, _zz_when_ArraySlice_l159_233_6};
  assign _zz__zz_realValue_0_233 = {1'd0, wReg};
  assign _zz__zz_realValue_0_233_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_233_1 = (_zz_realValue_0_233_2 + _zz_realValue_0_233_3);
  assign _zz_realValue_0_233_2 = {1'd0, wReg};
  assign _zz_realValue_0_233_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_233_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_233 = {1'd0, _zz_when_ArraySlice_l166_233_1};
  assign _zz_when_ArraySlice_l166_233_2 = (_zz_when_ArraySlice_l166_233_3 + _zz_when_ArraySlice_l166_233_7);
  assign _zz_when_ArraySlice_l166_233_3 = (realValue_0_233 - _zz_when_ArraySlice_l166_233_4);
  assign _zz_when_ArraySlice_l166_233_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_233_5);
  assign _zz_when_ArraySlice_l166_233_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_233_5 = {3'd0, _zz_when_ArraySlice_l166_233_6};
  assign _zz_when_ArraySlice_l166_233_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_234 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_234_1);
  assign _zz_when_ArraySlice_l158_234_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_234_1 = {2'd0, _zz_when_ArraySlice_l158_234_2};
  assign _zz_when_ArraySlice_l158_234_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_234_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_234 = {1'd0, _zz_when_ArraySlice_l159_234_1};
  assign _zz_when_ArraySlice_l159_234_2 = (_zz_when_ArraySlice_l159_234_3 - _zz_when_ArraySlice_l159_234_4);
  assign _zz_when_ArraySlice_l159_234_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_234_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_234_5);
  assign _zz_when_ArraySlice_l159_234_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_234_5 = {2'd0, _zz_when_ArraySlice_l159_234_6};
  assign _zz__zz_realValue_0_234 = {1'd0, wReg};
  assign _zz__zz_realValue_0_234_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_234_1 = (_zz_realValue_0_234_2 + _zz_realValue_0_234_3);
  assign _zz_realValue_0_234_2 = {1'd0, wReg};
  assign _zz_realValue_0_234_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_234_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_234 = {1'd0, _zz_when_ArraySlice_l166_234_1};
  assign _zz_when_ArraySlice_l166_234_2 = (_zz_when_ArraySlice_l166_234_3 + _zz_when_ArraySlice_l166_234_7);
  assign _zz_when_ArraySlice_l166_234_3 = (realValue_0_234 - _zz_when_ArraySlice_l166_234_4);
  assign _zz_when_ArraySlice_l166_234_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_234_5);
  assign _zz_when_ArraySlice_l166_234_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_234_5 = {2'd0, _zz_when_ArraySlice_l166_234_6};
  assign _zz_when_ArraySlice_l166_234_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_235 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_235_1);
  assign _zz_when_ArraySlice_l158_235_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_235_1 = {2'd0, _zz_when_ArraySlice_l158_235_2};
  assign _zz_when_ArraySlice_l158_235_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_235_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_235 = {1'd0, _zz_when_ArraySlice_l159_235_1};
  assign _zz_when_ArraySlice_l159_235_2 = (_zz_when_ArraySlice_l159_235_3 - _zz_when_ArraySlice_l159_235_4);
  assign _zz_when_ArraySlice_l159_235_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_235_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_235_5);
  assign _zz_when_ArraySlice_l159_235_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_235_5 = {2'd0, _zz_when_ArraySlice_l159_235_6};
  assign _zz__zz_realValue_0_235 = {1'd0, wReg};
  assign _zz__zz_realValue_0_235_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_235_1 = (_zz_realValue_0_235_2 + _zz_realValue_0_235_3);
  assign _zz_realValue_0_235_2 = {1'd0, wReg};
  assign _zz_realValue_0_235_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_235_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_235 = {1'd0, _zz_when_ArraySlice_l166_235_1};
  assign _zz_when_ArraySlice_l166_235_2 = (_zz_when_ArraySlice_l166_235_3 + _zz_when_ArraySlice_l166_235_7);
  assign _zz_when_ArraySlice_l166_235_3 = (realValue_0_235 - _zz_when_ArraySlice_l166_235_4);
  assign _zz_when_ArraySlice_l166_235_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_235_5);
  assign _zz_when_ArraySlice_l166_235_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_235_5 = {2'd0, _zz_when_ArraySlice_l166_235_6};
  assign _zz_when_ArraySlice_l166_235_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_236 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_236_1);
  assign _zz_when_ArraySlice_l158_236_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_236_1 = {1'd0, _zz_when_ArraySlice_l158_236_2};
  assign _zz_when_ArraySlice_l158_236_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_236_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_236 = {1'd0, _zz_when_ArraySlice_l159_236_1};
  assign _zz_when_ArraySlice_l159_236_2 = (_zz_when_ArraySlice_l159_236_3 - _zz_when_ArraySlice_l159_236_4);
  assign _zz_when_ArraySlice_l159_236_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_236_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_236_5);
  assign _zz_when_ArraySlice_l159_236_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_236_5 = {1'd0, _zz_when_ArraySlice_l159_236_6};
  assign _zz__zz_realValue_0_236 = {1'd0, wReg};
  assign _zz__zz_realValue_0_236_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_236_1 = (_zz_realValue_0_236_2 + _zz_realValue_0_236_3);
  assign _zz_realValue_0_236_2 = {1'd0, wReg};
  assign _zz_realValue_0_236_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_236_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_236 = {1'd0, _zz_when_ArraySlice_l166_236_1};
  assign _zz_when_ArraySlice_l166_236_2 = (_zz_when_ArraySlice_l166_236_3 + _zz_when_ArraySlice_l166_236_7);
  assign _zz_when_ArraySlice_l166_236_3 = (realValue_0_236 - _zz_when_ArraySlice_l166_236_4);
  assign _zz_when_ArraySlice_l166_236_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_236_5);
  assign _zz_when_ArraySlice_l166_236_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_236_5 = {1'd0, _zz_when_ArraySlice_l166_236_6};
  assign _zz_when_ArraySlice_l166_236_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_237 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_237_1);
  assign _zz_when_ArraySlice_l158_237_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_237_1 = {1'd0, _zz_when_ArraySlice_l158_237_2};
  assign _zz_when_ArraySlice_l158_237_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_237_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_237 = {2'd0, _zz_when_ArraySlice_l159_237_1};
  assign _zz_when_ArraySlice_l159_237_2 = (_zz_when_ArraySlice_l159_237_3 - _zz_when_ArraySlice_l159_237_4);
  assign _zz_when_ArraySlice_l159_237_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_237_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_237_5);
  assign _zz_when_ArraySlice_l159_237_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_237_5 = {1'd0, _zz_when_ArraySlice_l159_237_6};
  assign _zz__zz_realValue_0_237 = {1'd0, wReg};
  assign _zz__zz_realValue_0_237_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_237_1 = (_zz_realValue_0_237_2 + _zz_realValue_0_237_3);
  assign _zz_realValue_0_237_2 = {1'd0, wReg};
  assign _zz_realValue_0_237_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_237_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_237 = {2'd0, _zz_when_ArraySlice_l166_237_1};
  assign _zz_when_ArraySlice_l166_237_2 = (_zz_when_ArraySlice_l166_237_3 + _zz_when_ArraySlice_l166_237_7);
  assign _zz_when_ArraySlice_l166_237_3 = (realValue_0_237 - _zz_when_ArraySlice_l166_237_4);
  assign _zz_when_ArraySlice_l166_237_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_237_5);
  assign _zz_when_ArraySlice_l166_237_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_237_5 = {1'd0, _zz_when_ArraySlice_l166_237_6};
  assign _zz_when_ArraySlice_l166_237_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_238 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_238_1);
  assign _zz_when_ArraySlice_l158_238_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_238_1 = {1'd0, _zz_when_ArraySlice_l158_238_2};
  assign _zz_when_ArraySlice_l158_238_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_238_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_238 = {2'd0, _zz_when_ArraySlice_l159_238_1};
  assign _zz_when_ArraySlice_l159_238_2 = (_zz_when_ArraySlice_l159_238_3 - _zz_when_ArraySlice_l159_238_4);
  assign _zz_when_ArraySlice_l159_238_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_238_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_238_5);
  assign _zz_when_ArraySlice_l159_238_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_238_5 = {1'd0, _zz_when_ArraySlice_l159_238_6};
  assign _zz__zz_realValue_0_238 = {1'd0, wReg};
  assign _zz__zz_realValue_0_238_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_238_1 = (_zz_realValue_0_238_2 + _zz_realValue_0_238_3);
  assign _zz_realValue_0_238_2 = {1'd0, wReg};
  assign _zz_realValue_0_238_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_238_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_238 = {2'd0, _zz_when_ArraySlice_l166_238_1};
  assign _zz_when_ArraySlice_l166_238_2 = (_zz_when_ArraySlice_l166_238_3 + _zz_when_ArraySlice_l166_238_7);
  assign _zz_when_ArraySlice_l166_238_3 = (realValue_0_238 - _zz_when_ArraySlice_l166_238_4);
  assign _zz_when_ArraySlice_l166_238_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_238_5);
  assign _zz_when_ArraySlice_l166_238_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_238_5 = {1'd0, _zz_when_ArraySlice_l166_238_6};
  assign _zz_when_ArraySlice_l166_238_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_239 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_239_1);
  assign _zz_when_ArraySlice_l158_239_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_239_1 = {1'd0, _zz_when_ArraySlice_l158_239_2};
  assign _zz_when_ArraySlice_l158_239_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_239_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_239 = {3'd0, _zz_when_ArraySlice_l159_239_1};
  assign _zz_when_ArraySlice_l159_239_2 = (_zz_when_ArraySlice_l159_239_3 - _zz_when_ArraySlice_l159_239_4);
  assign _zz_when_ArraySlice_l159_239_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_239_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_239_5);
  assign _zz_when_ArraySlice_l159_239_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_239_5 = {1'd0, _zz_when_ArraySlice_l159_239_6};
  assign _zz__zz_realValue_0_239 = {1'd0, wReg};
  assign _zz__zz_realValue_0_239_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_239_1 = (_zz_realValue_0_239_2 + _zz_realValue_0_239_3);
  assign _zz_realValue_0_239_2 = {1'd0, wReg};
  assign _zz_realValue_0_239_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_239_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_239 = {3'd0, _zz_when_ArraySlice_l166_239_1};
  assign _zz_when_ArraySlice_l166_239_2 = (_zz_when_ArraySlice_l166_239_3 + _zz_when_ArraySlice_l166_239_7);
  assign _zz_when_ArraySlice_l166_239_3 = (realValue_0_239 - _zz_when_ArraySlice_l166_239_4);
  assign _zz_when_ArraySlice_l166_239_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_239_5);
  assign _zz_when_ArraySlice_l166_239_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_239_5 = {1'd0, _zz_when_ArraySlice_l166_239_6};
  assign _zz_when_ArraySlice_l166_239_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_1_2 = (_zz_when_ArraySlice_l260_1_3 + _zz_when_ArraySlice_l260_1_7);
  assign _zz_when_ArraySlice_l260_1_3 = (_zz_when_ArraySlice_l260_1_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l260_1_5);
  assign _zz_when_ArraySlice_l260_1_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_1_5 = {1'd0, _zz_when_ArraySlice_l260_1_6};
  assign _zz_when_ArraySlice_l260_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l260_1_7 = {3'd0, _zz_when_ArraySlice_l260_1_8};
  assign _zz_when_ArraySlice_l263_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_1_2 = (_zz_when_ArraySlice_l263_1_3 + 8'h01);
  assign _zz_when_ArraySlice_l263_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l263_1_4);
  assign _zz_when_ArraySlice_l263_1_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_1_4 = {1'd0, _zz_when_ArraySlice_l263_1_5};
  assign _zz_selectReadFifo_1_22 = (selectReadFifo_1 + _zz_selectReadFifo_1_23);
  assign _zz_selectReadFifo_1_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_23 = {1'd0, _zz_selectReadFifo_1_24};
  assign _zz_when_ArraySlice_l270_1_1 = (_zz_when_ArraySlice_l270_1_2 % aReg);
  assign _zz_when_ArraySlice_l270_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l274_1_4);
  assign _zz_when_ArraySlice_l274_1_2 = _zz_when_ArraySlice_l274_1_3[6:0];
  assign _zz_when_ArraySlice_l274_1_5 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l274_1_4 = {3'd0, _zz_when_ArraySlice_l274_1_5};
  assign _zz_when_ArraySlice_l275_1_2 = (_zz_when_ArraySlice_l275_1_3 - _zz_when_ArraySlice_l275_1_4);
  assign _zz_when_ArraySlice_l275_1_1 = {5'd0, _zz_when_ArraySlice_l275_1_2};
  assign _zz_when_ArraySlice_l275_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_1_5 = 1'b1;
  assign _zz_when_ArraySlice_l275_1_4 = {7'd0, _zz_when_ArraySlice_l275_1_5};
  assign _zz__zz_realValue1_0_28 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_28_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_28_1 = (_zz_realValue1_0_28_2 + _zz_realValue1_0_28_3);
  assign _zz_realValue1_0_28_2 = {1'd0, hReg};
  assign _zz_realValue1_0_28_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l277_1_1 = {1'd0, _zz_when_ArraySlice_l277_1_2};
  assign _zz_when_ArraySlice_l277_1_3 = (realValue1_0_28 / aReg);
  assign _zz_selectReadFifo_1_25 = (selectReadFifo_1 - _zz_selectReadFifo_1_26);
  assign _zz_selectReadFifo_1_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_240 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_240_1);
  assign _zz_when_ArraySlice_l158_240_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_240_1 = {4'd0, _zz_when_ArraySlice_l158_240_2};
  assign _zz_when_ArraySlice_l158_240_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_240 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_240_1 = (_zz_when_ArraySlice_l159_240_2 - _zz_when_ArraySlice_l159_240_3);
  assign _zz_when_ArraySlice_l159_240_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_240_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_240_4);
  assign _zz_when_ArraySlice_l159_240_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_240_4 = {4'd0, _zz_when_ArraySlice_l159_240_5};
  assign _zz__zz_realValue_0_240 = {1'd0, wReg};
  assign _zz__zz_realValue_0_240_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_240_1 = (_zz_realValue_0_240_2 + _zz_realValue_0_240_3);
  assign _zz_realValue_0_240_2 = {1'd0, wReg};
  assign _zz_realValue_0_240_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_240 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_240_1 = (_zz_when_ArraySlice_l166_240_2 + _zz_when_ArraySlice_l166_240_6);
  assign _zz_when_ArraySlice_l166_240_2 = (realValue_0_240 - _zz_when_ArraySlice_l166_240_3);
  assign _zz_when_ArraySlice_l166_240_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_240_4);
  assign _zz_when_ArraySlice_l166_240_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_240_4 = {4'd0, _zz_when_ArraySlice_l166_240_5};
  assign _zz_when_ArraySlice_l166_240_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_241 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_241_1);
  assign _zz_when_ArraySlice_l158_241_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_241_1 = {3'd0, _zz_when_ArraySlice_l158_241_2};
  assign _zz_when_ArraySlice_l158_241_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_241_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_241 = {1'd0, _zz_when_ArraySlice_l159_241_1};
  assign _zz_when_ArraySlice_l159_241_2 = (_zz_when_ArraySlice_l159_241_3 - _zz_when_ArraySlice_l159_241_4);
  assign _zz_when_ArraySlice_l159_241_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_241_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_241_5);
  assign _zz_when_ArraySlice_l159_241_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_241_5 = {3'd0, _zz_when_ArraySlice_l159_241_6};
  assign _zz__zz_realValue_0_241 = {1'd0, wReg};
  assign _zz__zz_realValue_0_241_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_241_1 = (_zz_realValue_0_241_2 + _zz_realValue_0_241_3);
  assign _zz_realValue_0_241_2 = {1'd0, wReg};
  assign _zz_realValue_0_241_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_241_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_241 = {1'd0, _zz_when_ArraySlice_l166_241_1};
  assign _zz_when_ArraySlice_l166_241_2 = (_zz_when_ArraySlice_l166_241_3 + _zz_when_ArraySlice_l166_241_7);
  assign _zz_when_ArraySlice_l166_241_3 = (realValue_0_241 - _zz_when_ArraySlice_l166_241_4);
  assign _zz_when_ArraySlice_l166_241_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_241_5);
  assign _zz_when_ArraySlice_l166_241_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_241_5 = {3'd0, _zz_when_ArraySlice_l166_241_6};
  assign _zz_when_ArraySlice_l166_241_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_242 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_242_1);
  assign _zz_when_ArraySlice_l158_242_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_242_1 = {2'd0, _zz_when_ArraySlice_l158_242_2};
  assign _zz_when_ArraySlice_l158_242_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_242_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_242 = {1'd0, _zz_when_ArraySlice_l159_242_1};
  assign _zz_when_ArraySlice_l159_242_2 = (_zz_when_ArraySlice_l159_242_3 - _zz_when_ArraySlice_l159_242_4);
  assign _zz_when_ArraySlice_l159_242_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_242_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_242_5);
  assign _zz_when_ArraySlice_l159_242_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_242_5 = {2'd0, _zz_when_ArraySlice_l159_242_6};
  assign _zz__zz_realValue_0_242 = {1'd0, wReg};
  assign _zz__zz_realValue_0_242_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_242_1 = (_zz_realValue_0_242_2 + _zz_realValue_0_242_3);
  assign _zz_realValue_0_242_2 = {1'd0, wReg};
  assign _zz_realValue_0_242_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_242_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_242 = {1'd0, _zz_when_ArraySlice_l166_242_1};
  assign _zz_when_ArraySlice_l166_242_2 = (_zz_when_ArraySlice_l166_242_3 + _zz_when_ArraySlice_l166_242_7);
  assign _zz_when_ArraySlice_l166_242_3 = (realValue_0_242 - _zz_when_ArraySlice_l166_242_4);
  assign _zz_when_ArraySlice_l166_242_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_242_5);
  assign _zz_when_ArraySlice_l166_242_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_242_5 = {2'd0, _zz_when_ArraySlice_l166_242_6};
  assign _zz_when_ArraySlice_l166_242_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_243 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_243_1);
  assign _zz_when_ArraySlice_l158_243_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_243_1 = {2'd0, _zz_when_ArraySlice_l158_243_2};
  assign _zz_when_ArraySlice_l158_243_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_243_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_243 = {1'd0, _zz_when_ArraySlice_l159_243_1};
  assign _zz_when_ArraySlice_l159_243_2 = (_zz_when_ArraySlice_l159_243_3 - _zz_when_ArraySlice_l159_243_4);
  assign _zz_when_ArraySlice_l159_243_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_243_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_243_5);
  assign _zz_when_ArraySlice_l159_243_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_243_5 = {2'd0, _zz_when_ArraySlice_l159_243_6};
  assign _zz__zz_realValue_0_243 = {1'd0, wReg};
  assign _zz__zz_realValue_0_243_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_243_1 = (_zz_realValue_0_243_2 + _zz_realValue_0_243_3);
  assign _zz_realValue_0_243_2 = {1'd0, wReg};
  assign _zz_realValue_0_243_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_243_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_243 = {1'd0, _zz_when_ArraySlice_l166_243_1};
  assign _zz_when_ArraySlice_l166_243_2 = (_zz_when_ArraySlice_l166_243_3 + _zz_when_ArraySlice_l166_243_7);
  assign _zz_when_ArraySlice_l166_243_3 = (realValue_0_243 - _zz_when_ArraySlice_l166_243_4);
  assign _zz_when_ArraySlice_l166_243_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_243_5);
  assign _zz_when_ArraySlice_l166_243_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_243_5 = {2'd0, _zz_when_ArraySlice_l166_243_6};
  assign _zz_when_ArraySlice_l166_243_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_244 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_244_1);
  assign _zz_when_ArraySlice_l158_244_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_244_1 = {1'd0, _zz_when_ArraySlice_l158_244_2};
  assign _zz_when_ArraySlice_l158_244_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_244_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_244 = {1'd0, _zz_when_ArraySlice_l159_244_1};
  assign _zz_when_ArraySlice_l159_244_2 = (_zz_when_ArraySlice_l159_244_3 - _zz_when_ArraySlice_l159_244_4);
  assign _zz_when_ArraySlice_l159_244_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_244_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_244_5);
  assign _zz_when_ArraySlice_l159_244_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_244_5 = {1'd0, _zz_when_ArraySlice_l159_244_6};
  assign _zz__zz_realValue_0_244 = {1'd0, wReg};
  assign _zz__zz_realValue_0_244_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_244_1 = (_zz_realValue_0_244_2 + _zz_realValue_0_244_3);
  assign _zz_realValue_0_244_2 = {1'd0, wReg};
  assign _zz_realValue_0_244_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_244_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_244 = {1'd0, _zz_when_ArraySlice_l166_244_1};
  assign _zz_when_ArraySlice_l166_244_2 = (_zz_when_ArraySlice_l166_244_3 + _zz_when_ArraySlice_l166_244_7);
  assign _zz_when_ArraySlice_l166_244_3 = (realValue_0_244 - _zz_when_ArraySlice_l166_244_4);
  assign _zz_when_ArraySlice_l166_244_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_244_5);
  assign _zz_when_ArraySlice_l166_244_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_244_5 = {1'd0, _zz_when_ArraySlice_l166_244_6};
  assign _zz_when_ArraySlice_l166_244_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_245 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_245_1);
  assign _zz_when_ArraySlice_l158_245_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_245_1 = {1'd0, _zz_when_ArraySlice_l158_245_2};
  assign _zz_when_ArraySlice_l158_245_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_245_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_245 = {2'd0, _zz_when_ArraySlice_l159_245_1};
  assign _zz_when_ArraySlice_l159_245_2 = (_zz_when_ArraySlice_l159_245_3 - _zz_when_ArraySlice_l159_245_4);
  assign _zz_when_ArraySlice_l159_245_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_245_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_245_5);
  assign _zz_when_ArraySlice_l159_245_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_245_5 = {1'd0, _zz_when_ArraySlice_l159_245_6};
  assign _zz__zz_realValue_0_245 = {1'd0, wReg};
  assign _zz__zz_realValue_0_245_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_245_1 = (_zz_realValue_0_245_2 + _zz_realValue_0_245_3);
  assign _zz_realValue_0_245_2 = {1'd0, wReg};
  assign _zz_realValue_0_245_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_245_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_245 = {2'd0, _zz_when_ArraySlice_l166_245_1};
  assign _zz_when_ArraySlice_l166_245_2 = (_zz_when_ArraySlice_l166_245_3 + _zz_when_ArraySlice_l166_245_7);
  assign _zz_when_ArraySlice_l166_245_3 = (realValue_0_245 - _zz_when_ArraySlice_l166_245_4);
  assign _zz_when_ArraySlice_l166_245_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_245_5);
  assign _zz_when_ArraySlice_l166_245_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_245_5 = {1'd0, _zz_when_ArraySlice_l166_245_6};
  assign _zz_when_ArraySlice_l166_245_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_246 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_246_1);
  assign _zz_when_ArraySlice_l158_246_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_246_1 = {1'd0, _zz_when_ArraySlice_l158_246_2};
  assign _zz_when_ArraySlice_l158_246_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_246_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_246 = {2'd0, _zz_when_ArraySlice_l159_246_1};
  assign _zz_when_ArraySlice_l159_246_2 = (_zz_when_ArraySlice_l159_246_3 - _zz_when_ArraySlice_l159_246_4);
  assign _zz_when_ArraySlice_l159_246_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_246_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_246_5);
  assign _zz_when_ArraySlice_l159_246_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_246_5 = {1'd0, _zz_when_ArraySlice_l159_246_6};
  assign _zz__zz_realValue_0_246 = {1'd0, wReg};
  assign _zz__zz_realValue_0_246_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_246_1 = (_zz_realValue_0_246_2 + _zz_realValue_0_246_3);
  assign _zz_realValue_0_246_2 = {1'd0, wReg};
  assign _zz_realValue_0_246_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_246_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_246 = {2'd0, _zz_when_ArraySlice_l166_246_1};
  assign _zz_when_ArraySlice_l166_246_2 = (_zz_when_ArraySlice_l166_246_3 + _zz_when_ArraySlice_l166_246_7);
  assign _zz_when_ArraySlice_l166_246_3 = (realValue_0_246 - _zz_when_ArraySlice_l166_246_4);
  assign _zz_when_ArraySlice_l166_246_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_246_5);
  assign _zz_when_ArraySlice_l166_246_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_246_5 = {1'd0, _zz_when_ArraySlice_l166_246_6};
  assign _zz_when_ArraySlice_l166_246_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_247 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_247_1);
  assign _zz_when_ArraySlice_l158_247_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_247_1 = {1'd0, _zz_when_ArraySlice_l158_247_2};
  assign _zz_when_ArraySlice_l158_247_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_247_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_247 = {3'd0, _zz_when_ArraySlice_l159_247_1};
  assign _zz_when_ArraySlice_l159_247_2 = (_zz_when_ArraySlice_l159_247_3 - _zz_when_ArraySlice_l159_247_4);
  assign _zz_when_ArraySlice_l159_247_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_247_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_247_5);
  assign _zz_when_ArraySlice_l159_247_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_247_5 = {1'd0, _zz_when_ArraySlice_l159_247_6};
  assign _zz__zz_realValue_0_247 = {1'd0, wReg};
  assign _zz__zz_realValue_0_247_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_247_1 = (_zz_realValue_0_247_2 + _zz_realValue_0_247_3);
  assign _zz_realValue_0_247_2 = {1'd0, wReg};
  assign _zz_realValue_0_247_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_247_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_247 = {3'd0, _zz_when_ArraySlice_l166_247_1};
  assign _zz_when_ArraySlice_l166_247_2 = (_zz_when_ArraySlice_l166_247_3 + _zz_when_ArraySlice_l166_247_7);
  assign _zz_when_ArraySlice_l166_247_3 = (realValue_0_247 - _zz_when_ArraySlice_l166_247_4);
  assign _zz_when_ArraySlice_l166_247_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_247_5);
  assign _zz_when_ArraySlice_l166_247_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_247_5 = {1'd0, _zz_when_ArraySlice_l166_247_6};
  assign _zz_when_ArraySlice_l166_247_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_1_2 = (_zz_when_ArraySlice_l285_1_3 + _zz_when_ArraySlice_l285_1_7);
  assign _zz_when_ArraySlice_l285_1_3 = (_zz_when_ArraySlice_l285_1_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_1_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l285_1_5);
  assign _zz_when_ArraySlice_l285_1_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_1_5 = {1'd0, _zz_when_ArraySlice_l285_1_6};
  assign _zz_when_ArraySlice_l285_1_8 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l285_1_7 = {3'd0, _zz_when_ArraySlice_l285_1_8};
  assign _zz_when_ArraySlice_l288_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_1_2 = (_zz_when_ArraySlice_l288_1_3 + 8'h01);
  assign _zz_when_ArraySlice_l288_1_3 = (selectReadFifo_1 + _zz_when_ArraySlice_l288_1_4);
  assign _zz_when_ArraySlice_l288_1_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_1_4 = {1'd0, _zz_when_ArraySlice_l288_1_5};
  assign _zz_selectReadFifo_1_27 = (selectReadFifo_1 + _zz_selectReadFifo_1_28);
  assign _zz_selectReadFifo_1_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_1_28 = {1'd0, _zz_selectReadFifo_1_29};
  assign _zz_when_ArraySlice_l295_1_1 = (_zz_when_ArraySlice_l295_1_2 % aReg);
  assign _zz_when_ArraySlice_l295_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_1_2 = (_zz_when_ArraySlice_l306_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l306_1_1 = {5'd0, _zz_when_ArraySlice_l306_1_2};
  assign _zz_when_ArraySlice_l306_1_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_29 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_29_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_29_1 = (_zz_realValue1_0_29_2 + _zz_realValue1_0_29_3);
  assign _zz_realValue1_0_29_2 = {1'd0, hReg};
  assign _zz_realValue1_0_29_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_1_2 = (outSliceNumb_1_value + 7'h01);
  assign _zz_when_ArraySlice_l307_1_1 = {1'd0, _zz_when_ArraySlice_l307_1_2};
  assign _zz_when_ArraySlice_l307_1_3 = (realValue1_0_29 / aReg);
  assign _zz_selectReadFifo_1_30 = (selectReadFifo_1 - _zz_selectReadFifo_1_31);
  assign _zz_selectReadFifo_1_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_248 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_248_1);
  assign _zz_when_ArraySlice_l158_248_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_248_1 = {4'd0, _zz_when_ArraySlice_l158_248_2};
  assign _zz_when_ArraySlice_l158_248_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_248 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_248_1 = (_zz_when_ArraySlice_l159_248_2 - _zz_when_ArraySlice_l159_248_3);
  assign _zz_when_ArraySlice_l159_248_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_248_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_248_4);
  assign _zz_when_ArraySlice_l159_248_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_248_4 = {4'd0, _zz_when_ArraySlice_l159_248_5};
  assign _zz__zz_realValue_0_248 = {1'd0, wReg};
  assign _zz__zz_realValue_0_248_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_248_1 = (_zz_realValue_0_248_2 + _zz_realValue_0_248_3);
  assign _zz_realValue_0_248_2 = {1'd0, wReg};
  assign _zz_realValue_0_248_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_248 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_248_1 = (_zz_when_ArraySlice_l166_248_2 + _zz_when_ArraySlice_l166_248_6);
  assign _zz_when_ArraySlice_l166_248_2 = (realValue_0_248 - _zz_when_ArraySlice_l166_248_3);
  assign _zz_when_ArraySlice_l166_248_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_248_4);
  assign _zz_when_ArraySlice_l166_248_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_248_4 = {4'd0, _zz_when_ArraySlice_l166_248_5};
  assign _zz_when_ArraySlice_l166_248_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_249 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_249_1);
  assign _zz_when_ArraySlice_l158_249_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_249_1 = {3'd0, _zz_when_ArraySlice_l158_249_2};
  assign _zz_when_ArraySlice_l158_249_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_249_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_249 = {1'd0, _zz_when_ArraySlice_l159_249_1};
  assign _zz_when_ArraySlice_l159_249_2 = (_zz_when_ArraySlice_l159_249_3 - _zz_when_ArraySlice_l159_249_4);
  assign _zz_when_ArraySlice_l159_249_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_249_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_249_5);
  assign _zz_when_ArraySlice_l159_249_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_249_5 = {3'd0, _zz_when_ArraySlice_l159_249_6};
  assign _zz__zz_realValue_0_249 = {1'd0, wReg};
  assign _zz__zz_realValue_0_249_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_249_1 = (_zz_realValue_0_249_2 + _zz_realValue_0_249_3);
  assign _zz_realValue_0_249_2 = {1'd0, wReg};
  assign _zz_realValue_0_249_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_249_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_249 = {1'd0, _zz_when_ArraySlice_l166_249_1};
  assign _zz_when_ArraySlice_l166_249_2 = (_zz_when_ArraySlice_l166_249_3 + _zz_when_ArraySlice_l166_249_7);
  assign _zz_when_ArraySlice_l166_249_3 = (realValue_0_249 - _zz_when_ArraySlice_l166_249_4);
  assign _zz_when_ArraySlice_l166_249_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_249_5);
  assign _zz_when_ArraySlice_l166_249_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_249_5 = {3'd0, _zz_when_ArraySlice_l166_249_6};
  assign _zz_when_ArraySlice_l166_249_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_250 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_250_1);
  assign _zz_when_ArraySlice_l158_250_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_250_1 = {2'd0, _zz_when_ArraySlice_l158_250_2};
  assign _zz_when_ArraySlice_l158_250_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_250_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_250 = {1'd0, _zz_when_ArraySlice_l159_250_1};
  assign _zz_when_ArraySlice_l159_250_2 = (_zz_when_ArraySlice_l159_250_3 - _zz_when_ArraySlice_l159_250_4);
  assign _zz_when_ArraySlice_l159_250_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_250_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_250_5);
  assign _zz_when_ArraySlice_l159_250_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_250_5 = {2'd0, _zz_when_ArraySlice_l159_250_6};
  assign _zz__zz_realValue_0_250 = {1'd0, wReg};
  assign _zz__zz_realValue_0_250_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_250_1 = (_zz_realValue_0_250_2 + _zz_realValue_0_250_3);
  assign _zz_realValue_0_250_2 = {1'd0, wReg};
  assign _zz_realValue_0_250_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_250_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_250 = {1'd0, _zz_when_ArraySlice_l166_250_1};
  assign _zz_when_ArraySlice_l166_250_2 = (_zz_when_ArraySlice_l166_250_3 + _zz_when_ArraySlice_l166_250_7);
  assign _zz_when_ArraySlice_l166_250_3 = (realValue_0_250 - _zz_when_ArraySlice_l166_250_4);
  assign _zz_when_ArraySlice_l166_250_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_250_5);
  assign _zz_when_ArraySlice_l166_250_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_250_5 = {2'd0, _zz_when_ArraySlice_l166_250_6};
  assign _zz_when_ArraySlice_l166_250_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_251 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_251_1);
  assign _zz_when_ArraySlice_l158_251_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_251_1 = {2'd0, _zz_when_ArraySlice_l158_251_2};
  assign _zz_when_ArraySlice_l158_251_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_251_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_251 = {1'd0, _zz_when_ArraySlice_l159_251_1};
  assign _zz_when_ArraySlice_l159_251_2 = (_zz_when_ArraySlice_l159_251_3 - _zz_when_ArraySlice_l159_251_4);
  assign _zz_when_ArraySlice_l159_251_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_251_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_251_5);
  assign _zz_when_ArraySlice_l159_251_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_251_5 = {2'd0, _zz_when_ArraySlice_l159_251_6};
  assign _zz__zz_realValue_0_251 = {1'd0, wReg};
  assign _zz__zz_realValue_0_251_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_251_1 = (_zz_realValue_0_251_2 + _zz_realValue_0_251_3);
  assign _zz_realValue_0_251_2 = {1'd0, wReg};
  assign _zz_realValue_0_251_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_251_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_251 = {1'd0, _zz_when_ArraySlice_l166_251_1};
  assign _zz_when_ArraySlice_l166_251_2 = (_zz_when_ArraySlice_l166_251_3 + _zz_when_ArraySlice_l166_251_7);
  assign _zz_when_ArraySlice_l166_251_3 = (realValue_0_251 - _zz_when_ArraySlice_l166_251_4);
  assign _zz_when_ArraySlice_l166_251_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_251_5);
  assign _zz_when_ArraySlice_l166_251_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_251_5 = {2'd0, _zz_when_ArraySlice_l166_251_6};
  assign _zz_when_ArraySlice_l166_251_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_252 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_252_1);
  assign _zz_when_ArraySlice_l158_252_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_252_1 = {1'd0, _zz_when_ArraySlice_l158_252_2};
  assign _zz_when_ArraySlice_l158_252_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_252_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_252 = {1'd0, _zz_when_ArraySlice_l159_252_1};
  assign _zz_when_ArraySlice_l159_252_2 = (_zz_when_ArraySlice_l159_252_3 - _zz_when_ArraySlice_l159_252_4);
  assign _zz_when_ArraySlice_l159_252_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_252_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_252_5);
  assign _zz_when_ArraySlice_l159_252_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_252_5 = {1'd0, _zz_when_ArraySlice_l159_252_6};
  assign _zz__zz_realValue_0_252 = {1'd0, wReg};
  assign _zz__zz_realValue_0_252_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_252_1 = (_zz_realValue_0_252_2 + _zz_realValue_0_252_3);
  assign _zz_realValue_0_252_2 = {1'd0, wReg};
  assign _zz_realValue_0_252_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_252_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_252 = {1'd0, _zz_when_ArraySlice_l166_252_1};
  assign _zz_when_ArraySlice_l166_252_2 = (_zz_when_ArraySlice_l166_252_3 + _zz_when_ArraySlice_l166_252_7);
  assign _zz_when_ArraySlice_l166_252_3 = (realValue_0_252 - _zz_when_ArraySlice_l166_252_4);
  assign _zz_when_ArraySlice_l166_252_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_252_5);
  assign _zz_when_ArraySlice_l166_252_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_252_5 = {1'd0, _zz_when_ArraySlice_l166_252_6};
  assign _zz_when_ArraySlice_l166_252_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_253 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_253_1);
  assign _zz_when_ArraySlice_l158_253_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_253_1 = {1'd0, _zz_when_ArraySlice_l158_253_2};
  assign _zz_when_ArraySlice_l158_253_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_253_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_253 = {2'd0, _zz_when_ArraySlice_l159_253_1};
  assign _zz_when_ArraySlice_l159_253_2 = (_zz_when_ArraySlice_l159_253_3 - _zz_when_ArraySlice_l159_253_4);
  assign _zz_when_ArraySlice_l159_253_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_253_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_253_5);
  assign _zz_when_ArraySlice_l159_253_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_253_5 = {1'd0, _zz_when_ArraySlice_l159_253_6};
  assign _zz__zz_realValue_0_253 = {1'd0, wReg};
  assign _zz__zz_realValue_0_253_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_253_1 = (_zz_realValue_0_253_2 + _zz_realValue_0_253_3);
  assign _zz_realValue_0_253_2 = {1'd0, wReg};
  assign _zz_realValue_0_253_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_253_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_253 = {2'd0, _zz_when_ArraySlice_l166_253_1};
  assign _zz_when_ArraySlice_l166_253_2 = (_zz_when_ArraySlice_l166_253_3 + _zz_when_ArraySlice_l166_253_7);
  assign _zz_when_ArraySlice_l166_253_3 = (realValue_0_253 - _zz_when_ArraySlice_l166_253_4);
  assign _zz_when_ArraySlice_l166_253_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_253_5);
  assign _zz_when_ArraySlice_l166_253_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_253_5 = {1'd0, _zz_when_ArraySlice_l166_253_6};
  assign _zz_when_ArraySlice_l166_253_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_254 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_254_1);
  assign _zz_when_ArraySlice_l158_254_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_254_1 = {1'd0, _zz_when_ArraySlice_l158_254_2};
  assign _zz_when_ArraySlice_l158_254_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_254_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_254 = {2'd0, _zz_when_ArraySlice_l159_254_1};
  assign _zz_when_ArraySlice_l159_254_2 = (_zz_when_ArraySlice_l159_254_3 - _zz_when_ArraySlice_l159_254_4);
  assign _zz_when_ArraySlice_l159_254_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_254_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_254_5);
  assign _zz_when_ArraySlice_l159_254_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_254_5 = {1'd0, _zz_when_ArraySlice_l159_254_6};
  assign _zz__zz_realValue_0_254 = {1'd0, wReg};
  assign _zz__zz_realValue_0_254_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_254_1 = (_zz_realValue_0_254_2 + _zz_realValue_0_254_3);
  assign _zz_realValue_0_254_2 = {1'd0, wReg};
  assign _zz_realValue_0_254_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_254_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_254 = {2'd0, _zz_when_ArraySlice_l166_254_1};
  assign _zz_when_ArraySlice_l166_254_2 = (_zz_when_ArraySlice_l166_254_3 + _zz_when_ArraySlice_l166_254_7);
  assign _zz_when_ArraySlice_l166_254_3 = (realValue_0_254 - _zz_when_ArraySlice_l166_254_4);
  assign _zz_when_ArraySlice_l166_254_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_254_5);
  assign _zz_when_ArraySlice_l166_254_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_254_5 = {1'd0, _zz_when_ArraySlice_l166_254_6};
  assign _zz_when_ArraySlice_l166_254_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_255 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_255_1);
  assign _zz_when_ArraySlice_l158_255_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_255_1 = {1'd0, _zz_when_ArraySlice_l158_255_2};
  assign _zz_when_ArraySlice_l158_255_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_255_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_255 = {3'd0, _zz_when_ArraySlice_l159_255_1};
  assign _zz_when_ArraySlice_l159_255_2 = (_zz_when_ArraySlice_l159_255_3 - _zz_when_ArraySlice_l159_255_4);
  assign _zz_when_ArraySlice_l159_255_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_255_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_255_5);
  assign _zz_when_ArraySlice_l159_255_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_255_5 = {1'd0, _zz_when_ArraySlice_l159_255_6};
  assign _zz__zz_realValue_0_255 = {1'd0, wReg};
  assign _zz__zz_realValue_0_255_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_255_1 = (_zz_realValue_0_255_2 + _zz_realValue_0_255_3);
  assign _zz_realValue_0_255_2 = {1'd0, wReg};
  assign _zz_realValue_0_255_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_255_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_255 = {3'd0, _zz_when_ArraySlice_l166_255_1};
  assign _zz_when_ArraySlice_l166_255_2 = (_zz_when_ArraySlice_l166_255_3 + _zz_when_ArraySlice_l166_255_7);
  assign _zz_when_ArraySlice_l166_255_3 = (realValue_0_255 - _zz_when_ArraySlice_l166_255_4);
  assign _zz_when_ArraySlice_l166_255_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_255_5);
  assign _zz_when_ArraySlice_l166_255_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_255_5 = {1'd0, _zz_when_ArraySlice_l166_255_6};
  assign _zz_when_ArraySlice_l166_255_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_1_1 = (_zz_when_ArraySlice_l318_1_2 % aReg);
  assign _zz_when_ArraySlice_l318_1_2 = (handshakeTimes_1_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_1_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_1_2 = (selectReadFifo_1 + _zz_when_ArraySlice_l304_1_3);
  assign _zz_when_ArraySlice_l304_1_4 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l304_1_3 = {3'd0, _zz_when_ArraySlice_l304_1_4};
  assign _zz_when_ArraySlice_l325_1_2 = (_zz_when_ArraySlice_l325_1_3 - 8'h01);
  assign _zz_when_ArraySlice_l325_1_1 = {5'd0, _zz_when_ArraySlice_l325_1_2};
  assign _zz_when_ArraySlice_l325_1_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_2_1 = (selectReadFifo_2 + _zz_when_ArraySlice_l233_2_2);
  assign _zz_when_ArraySlice_l233_2_3 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l233_2_2 = {2'd0, _zz_when_ArraySlice_l233_2_3};
  assign _zz_when_ArraySlice_l233_2_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l234_2_4);
  assign _zz_when_ArraySlice_l234_2_2 = _zz_when_ArraySlice_l234_2_3[6:0];
  assign _zz_when_ArraySlice_l234_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l234_2_4 = {2'd0, _zz_when_ArraySlice_l234_2_5};
  assign _zz__zz_outputStreamArrayData_2_valid_1_2 = (bReg * 2'b10);
  assign _zz__zz_outputStreamArrayData_2_valid_1_1 = {2'd0, _zz__zz_outputStreamArrayData_2_valid_1_2};
  assign _zz__zz_13 = _zz_outputStreamArrayData_2_valid_1[6:0];
  assign _zz_outputStreamArrayData_2_valid_5 = _zz_outputStreamArrayData_2_valid_1[6:0];
  assign _zz_outputStreamArrayData_2_payload_3 = _zz_outputStreamArrayData_2_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l240_2_4);
  assign _zz_when_ArraySlice_l240_2_2 = _zz_when_ArraySlice_l240_2_3[6:0];
  assign _zz_when_ArraySlice_l240_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l240_2_4 = {2'd0, _zz_when_ArraySlice_l240_2_5};
  assign _zz_when_ArraySlice_l241_2_2 = (_zz_when_ArraySlice_l241_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l241_2_1 = {5'd0, _zz_when_ArraySlice_l241_2_2};
  assign _zz_when_ArraySlice_l241_2_3 = (bReg * aReg);
  assign _zz_selectReadFifo_2_16 = (selectReadFifo_2 - _zz_selectReadFifo_2_17);
  assign _zz_selectReadFifo_2_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_2 = (_zz_when_ArraySlice_l244_2_1 % aReg);
  assign _zz_when_ArraySlice_l244_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l249_2_4);
  assign _zz_when_ArraySlice_l249_2_2 = _zz_when_ArraySlice_l249_2_3[6:0];
  assign _zz_when_ArraySlice_l249_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l249_2_4 = {2'd0, _zz_when_ArraySlice_l249_2_5};
  assign _zz_when_ArraySlice_l250_2_2 = (_zz_when_ArraySlice_l250_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l250_2_1 = {5'd0, _zz_when_ArraySlice_l250_2_2};
  assign _zz_when_ArraySlice_l250_2_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_30 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_30_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_30_1 = (_zz_realValue1_0_30_2 + _zz_realValue1_0_30_3);
  assign _zz_realValue1_0_30_2 = {1'd0, hReg};
  assign _zz_realValue1_0_30_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l252_2_1 = {1'd0, _zz_when_ArraySlice_l252_2_2};
  assign _zz_when_ArraySlice_l252_2_3 = (realValue1_0_30 / aReg);
  assign _zz_selectReadFifo_2_18 = (selectReadFifo_2 - _zz_selectReadFifo_2_19);
  assign _zz_selectReadFifo_2_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_2_21 = 1'b1;
  assign _zz_selectReadFifo_2_20 = {7'd0, _zz_selectReadFifo_2_21};
  assign _zz_when_ArraySlice_l158_256 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_256_1);
  assign _zz_when_ArraySlice_l158_256_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_256_1 = {4'd0, _zz_when_ArraySlice_l158_256_2};
  assign _zz_when_ArraySlice_l158_256_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_256 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_256_1 = (_zz_when_ArraySlice_l159_256_2 - _zz_when_ArraySlice_l159_256_3);
  assign _zz_when_ArraySlice_l159_256_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_256_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_256_4);
  assign _zz_when_ArraySlice_l159_256_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_256_4 = {4'd0, _zz_when_ArraySlice_l159_256_5};
  assign _zz__zz_realValue_0_256 = {1'd0, wReg};
  assign _zz__zz_realValue_0_256_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_256_1 = (_zz_realValue_0_256_2 + _zz_realValue_0_256_3);
  assign _zz_realValue_0_256_2 = {1'd0, wReg};
  assign _zz_realValue_0_256_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_256 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_256_1 = (_zz_when_ArraySlice_l166_256_2 + _zz_when_ArraySlice_l166_256_6);
  assign _zz_when_ArraySlice_l166_256_2 = (realValue_0_256 - _zz_when_ArraySlice_l166_256_3);
  assign _zz_when_ArraySlice_l166_256_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_256_4);
  assign _zz_when_ArraySlice_l166_256_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_256_4 = {4'd0, _zz_when_ArraySlice_l166_256_5};
  assign _zz_when_ArraySlice_l166_256_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_257 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_257_1);
  assign _zz_when_ArraySlice_l158_257_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_257_1 = {3'd0, _zz_when_ArraySlice_l158_257_2};
  assign _zz_when_ArraySlice_l158_257_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_257_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_257 = {1'd0, _zz_when_ArraySlice_l159_257_1};
  assign _zz_when_ArraySlice_l159_257_2 = (_zz_when_ArraySlice_l159_257_3 - _zz_when_ArraySlice_l159_257_4);
  assign _zz_when_ArraySlice_l159_257_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_257_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_257_5);
  assign _zz_when_ArraySlice_l159_257_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_257_5 = {3'd0, _zz_when_ArraySlice_l159_257_6};
  assign _zz__zz_realValue_0_257 = {1'd0, wReg};
  assign _zz__zz_realValue_0_257_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_257_1 = (_zz_realValue_0_257_2 + _zz_realValue_0_257_3);
  assign _zz_realValue_0_257_2 = {1'd0, wReg};
  assign _zz_realValue_0_257_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_257_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_257 = {1'd0, _zz_when_ArraySlice_l166_257_1};
  assign _zz_when_ArraySlice_l166_257_2 = (_zz_when_ArraySlice_l166_257_3 + _zz_when_ArraySlice_l166_257_7);
  assign _zz_when_ArraySlice_l166_257_3 = (realValue_0_257 - _zz_when_ArraySlice_l166_257_4);
  assign _zz_when_ArraySlice_l166_257_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_257_5);
  assign _zz_when_ArraySlice_l166_257_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_257_5 = {3'd0, _zz_when_ArraySlice_l166_257_6};
  assign _zz_when_ArraySlice_l166_257_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_258 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_258_1);
  assign _zz_when_ArraySlice_l158_258_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_258_1 = {2'd0, _zz_when_ArraySlice_l158_258_2};
  assign _zz_when_ArraySlice_l158_258_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_258_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_258 = {1'd0, _zz_when_ArraySlice_l159_258_1};
  assign _zz_when_ArraySlice_l159_258_2 = (_zz_when_ArraySlice_l159_258_3 - _zz_when_ArraySlice_l159_258_4);
  assign _zz_when_ArraySlice_l159_258_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_258_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_258_5);
  assign _zz_when_ArraySlice_l159_258_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_258_5 = {2'd0, _zz_when_ArraySlice_l159_258_6};
  assign _zz__zz_realValue_0_258 = {1'd0, wReg};
  assign _zz__zz_realValue_0_258_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_258_1 = (_zz_realValue_0_258_2 + _zz_realValue_0_258_3);
  assign _zz_realValue_0_258_2 = {1'd0, wReg};
  assign _zz_realValue_0_258_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_258_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_258 = {1'd0, _zz_when_ArraySlice_l166_258_1};
  assign _zz_when_ArraySlice_l166_258_2 = (_zz_when_ArraySlice_l166_258_3 + _zz_when_ArraySlice_l166_258_7);
  assign _zz_when_ArraySlice_l166_258_3 = (realValue_0_258 - _zz_when_ArraySlice_l166_258_4);
  assign _zz_when_ArraySlice_l166_258_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_258_5);
  assign _zz_when_ArraySlice_l166_258_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_258_5 = {2'd0, _zz_when_ArraySlice_l166_258_6};
  assign _zz_when_ArraySlice_l166_258_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_259 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_259_1);
  assign _zz_when_ArraySlice_l158_259_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_259_1 = {2'd0, _zz_when_ArraySlice_l158_259_2};
  assign _zz_when_ArraySlice_l158_259_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_259_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_259 = {1'd0, _zz_when_ArraySlice_l159_259_1};
  assign _zz_when_ArraySlice_l159_259_2 = (_zz_when_ArraySlice_l159_259_3 - _zz_when_ArraySlice_l159_259_4);
  assign _zz_when_ArraySlice_l159_259_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_259_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_259_5);
  assign _zz_when_ArraySlice_l159_259_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_259_5 = {2'd0, _zz_when_ArraySlice_l159_259_6};
  assign _zz__zz_realValue_0_259 = {1'd0, wReg};
  assign _zz__zz_realValue_0_259_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_259_1 = (_zz_realValue_0_259_2 + _zz_realValue_0_259_3);
  assign _zz_realValue_0_259_2 = {1'd0, wReg};
  assign _zz_realValue_0_259_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_259_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_259 = {1'd0, _zz_when_ArraySlice_l166_259_1};
  assign _zz_when_ArraySlice_l166_259_2 = (_zz_when_ArraySlice_l166_259_3 + _zz_when_ArraySlice_l166_259_7);
  assign _zz_when_ArraySlice_l166_259_3 = (realValue_0_259 - _zz_when_ArraySlice_l166_259_4);
  assign _zz_when_ArraySlice_l166_259_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_259_5);
  assign _zz_when_ArraySlice_l166_259_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_259_5 = {2'd0, _zz_when_ArraySlice_l166_259_6};
  assign _zz_when_ArraySlice_l166_259_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_260 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_260_1);
  assign _zz_when_ArraySlice_l158_260_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_260_1 = {1'd0, _zz_when_ArraySlice_l158_260_2};
  assign _zz_when_ArraySlice_l158_260_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_260_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_260 = {1'd0, _zz_when_ArraySlice_l159_260_1};
  assign _zz_when_ArraySlice_l159_260_2 = (_zz_when_ArraySlice_l159_260_3 - _zz_when_ArraySlice_l159_260_4);
  assign _zz_when_ArraySlice_l159_260_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_260_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_260_5);
  assign _zz_when_ArraySlice_l159_260_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_260_5 = {1'd0, _zz_when_ArraySlice_l159_260_6};
  assign _zz__zz_realValue_0_260 = {1'd0, wReg};
  assign _zz__zz_realValue_0_260_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_260_1 = (_zz_realValue_0_260_2 + _zz_realValue_0_260_3);
  assign _zz_realValue_0_260_2 = {1'd0, wReg};
  assign _zz_realValue_0_260_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_260_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_260 = {1'd0, _zz_when_ArraySlice_l166_260_1};
  assign _zz_when_ArraySlice_l166_260_2 = (_zz_when_ArraySlice_l166_260_3 + _zz_when_ArraySlice_l166_260_7);
  assign _zz_when_ArraySlice_l166_260_3 = (realValue_0_260 - _zz_when_ArraySlice_l166_260_4);
  assign _zz_when_ArraySlice_l166_260_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_260_5);
  assign _zz_when_ArraySlice_l166_260_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_260_5 = {1'd0, _zz_when_ArraySlice_l166_260_6};
  assign _zz_when_ArraySlice_l166_260_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_261 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_261_1);
  assign _zz_when_ArraySlice_l158_261_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_261_1 = {1'd0, _zz_when_ArraySlice_l158_261_2};
  assign _zz_when_ArraySlice_l158_261_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_261_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_261 = {2'd0, _zz_when_ArraySlice_l159_261_1};
  assign _zz_when_ArraySlice_l159_261_2 = (_zz_when_ArraySlice_l159_261_3 - _zz_when_ArraySlice_l159_261_4);
  assign _zz_when_ArraySlice_l159_261_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_261_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_261_5);
  assign _zz_when_ArraySlice_l159_261_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_261_5 = {1'd0, _zz_when_ArraySlice_l159_261_6};
  assign _zz__zz_realValue_0_261 = {1'd0, wReg};
  assign _zz__zz_realValue_0_261_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_261_1 = (_zz_realValue_0_261_2 + _zz_realValue_0_261_3);
  assign _zz_realValue_0_261_2 = {1'd0, wReg};
  assign _zz_realValue_0_261_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_261_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_261 = {2'd0, _zz_when_ArraySlice_l166_261_1};
  assign _zz_when_ArraySlice_l166_261_2 = (_zz_when_ArraySlice_l166_261_3 + _zz_when_ArraySlice_l166_261_7);
  assign _zz_when_ArraySlice_l166_261_3 = (realValue_0_261 - _zz_when_ArraySlice_l166_261_4);
  assign _zz_when_ArraySlice_l166_261_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_261_5);
  assign _zz_when_ArraySlice_l166_261_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_261_5 = {1'd0, _zz_when_ArraySlice_l166_261_6};
  assign _zz_when_ArraySlice_l166_261_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_262 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_262_1);
  assign _zz_when_ArraySlice_l158_262_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_262_1 = {1'd0, _zz_when_ArraySlice_l158_262_2};
  assign _zz_when_ArraySlice_l158_262_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_262_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_262 = {2'd0, _zz_when_ArraySlice_l159_262_1};
  assign _zz_when_ArraySlice_l159_262_2 = (_zz_when_ArraySlice_l159_262_3 - _zz_when_ArraySlice_l159_262_4);
  assign _zz_when_ArraySlice_l159_262_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_262_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_262_5);
  assign _zz_when_ArraySlice_l159_262_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_262_5 = {1'd0, _zz_when_ArraySlice_l159_262_6};
  assign _zz__zz_realValue_0_262 = {1'd0, wReg};
  assign _zz__zz_realValue_0_262_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_262_1 = (_zz_realValue_0_262_2 + _zz_realValue_0_262_3);
  assign _zz_realValue_0_262_2 = {1'd0, wReg};
  assign _zz_realValue_0_262_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_262_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_262 = {2'd0, _zz_when_ArraySlice_l166_262_1};
  assign _zz_when_ArraySlice_l166_262_2 = (_zz_when_ArraySlice_l166_262_3 + _zz_when_ArraySlice_l166_262_7);
  assign _zz_when_ArraySlice_l166_262_3 = (realValue_0_262 - _zz_when_ArraySlice_l166_262_4);
  assign _zz_when_ArraySlice_l166_262_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_262_5);
  assign _zz_when_ArraySlice_l166_262_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_262_5 = {1'd0, _zz_when_ArraySlice_l166_262_6};
  assign _zz_when_ArraySlice_l166_262_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_263 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_263_1);
  assign _zz_when_ArraySlice_l158_263_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_263_1 = {1'd0, _zz_when_ArraySlice_l158_263_2};
  assign _zz_when_ArraySlice_l158_263_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_263_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_263 = {3'd0, _zz_when_ArraySlice_l159_263_1};
  assign _zz_when_ArraySlice_l159_263_2 = (_zz_when_ArraySlice_l159_263_3 - _zz_when_ArraySlice_l159_263_4);
  assign _zz_when_ArraySlice_l159_263_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_263_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_263_5);
  assign _zz_when_ArraySlice_l159_263_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_263_5 = {1'd0, _zz_when_ArraySlice_l159_263_6};
  assign _zz__zz_realValue_0_263 = {1'd0, wReg};
  assign _zz__zz_realValue_0_263_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_263_1 = (_zz_realValue_0_263_2 + _zz_realValue_0_263_3);
  assign _zz_realValue_0_263_2 = {1'd0, wReg};
  assign _zz_realValue_0_263_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_263_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_263 = {3'd0, _zz_when_ArraySlice_l166_263_1};
  assign _zz_when_ArraySlice_l166_263_2 = (_zz_when_ArraySlice_l166_263_3 + _zz_when_ArraySlice_l166_263_7);
  assign _zz_when_ArraySlice_l166_263_3 = (realValue_0_263 - _zz_when_ArraySlice_l166_263_4);
  assign _zz_when_ArraySlice_l166_263_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_263_5);
  assign _zz_when_ArraySlice_l166_263_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_263_5 = {1'd0, _zz_when_ArraySlice_l166_263_6};
  assign _zz_when_ArraySlice_l166_263_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_2_2 = (_zz_when_ArraySlice_l260_2_3 + _zz_when_ArraySlice_l260_2_7);
  assign _zz_when_ArraySlice_l260_2_3 = (_zz_when_ArraySlice_l260_2_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l260_2_5);
  assign _zz_when_ArraySlice_l260_2_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_2_5 = {1'd0, _zz_when_ArraySlice_l260_2_6};
  assign _zz_when_ArraySlice_l260_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l260_2_7 = {2'd0, _zz_when_ArraySlice_l260_2_8};
  assign _zz_when_ArraySlice_l263_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_2_2 = (_zz_when_ArraySlice_l263_2_3 + 8'h01);
  assign _zz_when_ArraySlice_l263_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l263_2_4);
  assign _zz_when_ArraySlice_l263_2_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_2_4 = {1'd0, _zz_when_ArraySlice_l263_2_5};
  assign _zz_selectReadFifo_2_22 = (selectReadFifo_2 + _zz_selectReadFifo_2_23);
  assign _zz_selectReadFifo_2_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_23 = {1'd0, _zz_selectReadFifo_2_24};
  assign _zz_when_ArraySlice_l270_2 = (_zz_when_ArraySlice_l270_2_1 % aReg);
  assign _zz_when_ArraySlice_l270_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l274_2_4);
  assign _zz_when_ArraySlice_l274_2_2 = _zz_when_ArraySlice_l274_2_3[6:0];
  assign _zz_when_ArraySlice_l274_2_5 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l274_2_4 = {2'd0, _zz_when_ArraySlice_l274_2_5};
  assign _zz_when_ArraySlice_l275_2_2 = (_zz_when_ArraySlice_l275_2_3 - _zz_when_ArraySlice_l275_2_4);
  assign _zz_when_ArraySlice_l275_2_1 = {5'd0, _zz_when_ArraySlice_l275_2_2};
  assign _zz_when_ArraySlice_l275_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_2_5 = 1'b1;
  assign _zz_when_ArraySlice_l275_2_4 = {7'd0, _zz_when_ArraySlice_l275_2_5};
  assign _zz__zz_realValue1_0_31 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_31_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_31_1 = (_zz_realValue1_0_31_2 + _zz_realValue1_0_31_3);
  assign _zz_realValue1_0_31_2 = {1'd0, hReg};
  assign _zz_realValue1_0_31_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l277_2_1 = {1'd0, _zz_when_ArraySlice_l277_2_2};
  assign _zz_when_ArraySlice_l277_2_3 = (realValue1_0_31 / aReg);
  assign _zz_selectReadFifo_2_25 = (selectReadFifo_2 - _zz_selectReadFifo_2_26);
  assign _zz_selectReadFifo_2_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_264 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_264_1);
  assign _zz_when_ArraySlice_l158_264_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_264_1 = {4'd0, _zz_when_ArraySlice_l158_264_2};
  assign _zz_when_ArraySlice_l158_264_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_264 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_264_1 = (_zz_when_ArraySlice_l159_264_2 - _zz_when_ArraySlice_l159_264_3);
  assign _zz_when_ArraySlice_l159_264_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_264_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_264_4);
  assign _zz_when_ArraySlice_l159_264_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_264_4 = {4'd0, _zz_when_ArraySlice_l159_264_5};
  assign _zz__zz_realValue_0_264 = {1'd0, wReg};
  assign _zz__zz_realValue_0_264_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_264_1 = (_zz_realValue_0_264_2 + _zz_realValue_0_264_3);
  assign _zz_realValue_0_264_2 = {1'd0, wReg};
  assign _zz_realValue_0_264_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_264 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_264_1 = (_zz_when_ArraySlice_l166_264_2 + _zz_when_ArraySlice_l166_264_6);
  assign _zz_when_ArraySlice_l166_264_2 = (realValue_0_264 - _zz_when_ArraySlice_l166_264_3);
  assign _zz_when_ArraySlice_l166_264_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_264_4);
  assign _zz_when_ArraySlice_l166_264_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_264_4 = {4'd0, _zz_when_ArraySlice_l166_264_5};
  assign _zz_when_ArraySlice_l166_264_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_265 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_265_1);
  assign _zz_when_ArraySlice_l158_265_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_265_1 = {3'd0, _zz_when_ArraySlice_l158_265_2};
  assign _zz_when_ArraySlice_l158_265_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_265_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_265 = {1'd0, _zz_when_ArraySlice_l159_265_1};
  assign _zz_when_ArraySlice_l159_265_2 = (_zz_when_ArraySlice_l159_265_3 - _zz_when_ArraySlice_l159_265_4);
  assign _zz_when_ArraySlice_l159_265_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_265_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_265_5);
  assign _zz_when_ArraySlice_l159_265_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_265_5 = {3'd0, _zz_when_ArraySlice_l159_265_6};
  assign _zz__zz_realValue_0_265 = {1'd0, wReg};
  assign _zz__zz_realValue_0_265_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_265_1 = (_zz_realValue_0_265_2 + _zz_realValue_0_265_3);
  assign _zz_realValue_0_265_2 = {1'd0, wReg};
  assign _zz_realValue_0_265_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_265_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_265 = {1'd0, _zz_when_ArraySlice_l166_265_1};
  assign _zz_when_ArraySlice_l166_265_2 = (_zz_when_ArraySlice_l166_265_3 + _zz_when_ArraySlice_l166_265_7);
  assign _zz_when_ArraySlice_l166_265_3 = (realValue_0_265 - _zz_when_ArraySlice_l166_265_4);
  assign _zz_when_ArraySlice_l166_265_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_265_5);
  assign _zz_when_ArraySlice_l166_265_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_265_5 = {3'd0, _zz_when_ArraySlice_l166_265_6};
  assign _zz_when_ArraySlice_l166_265_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_266 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_266_1);
  assign _zz_when_ArraySlice_l158_266_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_266_1 = {2'd0, _zz_when_ArraySlice_l158_266_2};
  assign _zz_when_ArraySlice_l158_266_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_266_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_266 = {1'd0, _zz_when_ArraySlice_l159_266_1};
  assign _zz_when_ArraySlice_l159_266_2 = (_zz_when_ArraySlice_l159_266_3 - _zz_when_ArraySlice_l159_266_4);
  assign _zz_when_ArraySlice_l159_266_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_266_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_266_5);
  assign _zz_when_ArraySlice_l159_266_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_266_5 = {2'd0, _zz_when_ArraySlice_l159_266_6};
  assign _zz__zz_realValue_0_266 = {1'd0, wReg};
  assign _zz__zz_realValue_0_266_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_266_1 = (_zz_realValue_0_266_2 + _zz_realValue_0_266_3);
  assign _zz_realValue_0_266_2 = {1'd0, wReg};
  assign _zz_realValue_0_266_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_266_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_266 = {1'd0, _zz_when_ArraySlice_l166_266_1};
  assign _zz_when_ArraySlice_l166_266_2 = (_zz_when_ArraySlice_l166_266_3 + _zz_when_ArraySlice_l166_266_7);
  assign _zz_when_ArraySlice_l166_266_3 = (realValue_0_266 - _zz_when_ArraySlice_l166_266_4);
  assign _zz_when_ArraySlice_l166_266_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_266_5);
  assign _zz_when_ArraySlice_l166_266_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_266_5 = {2'd0, _zz_when_ArraySlice_l166_266_6};
  assign _zz_when_ArraySlice_l166_266_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_267 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_267_1);
  assign _zz_when_ArraySlice_l158_267_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_267_1 = {2'd0, _zz_when_ArraySlice_l158_267_2};
  assign _zz_when_ArraySlice_l158_267_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_267_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_267 = {1'd0, _zz_when_ArraySlice_l159_267_1};
  assign _zz_when_ArraySlice_l159_267_2 = (_zz_when_ArraySlice_l159_267_3 - _zz_when_ArraySlice_l159_267_4);
  assign _zz_when_ArraySlice_l159_267_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_267_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_267_5);
  assign _zz_when_ArraySlice_l159_267_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_267_5 = {2'd0, _zz_when_ArraySlice_l159_267_6};
  assign _zz__zz_realValue_0_267 = {1'd0, wReg};
  assign _zz__zz_realValue_0_267_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_267_1 = (_zz_realValue_0_267_2 + _zz_realValue_0_267_3);
  assign _zz_realValue_0_267_2 = {1'd0, wReg};
  assign _zz_realValue_0_267_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_267_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_267 = {1'd0, _zz_when_ArraySlice_l166_267_1};
  assign _zz_when_ArraySlice_l166_267_2 = (_zz_when_ArraySlice_l166_267_3 + _zz_when_ArraySlice_l166_267_7);
  assign _zz_when_ArraySlice_l166_267_3 = (realValue_0_267 - _zz_when_ArraySlice_l166_267_4);
  assign _zz_when_ArraySlice_l166_267_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_267_5);
  assign _zz_when_ArraySlice_l166_267_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_267_5 = {2'd0, _zz_when_ArraySlice_l166_267_6};
  assign _zz_when_ArraySlice_l166_267_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_268 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_268_1);
  assign _zz_when_ArraySlice_l158_268_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_268_1 = {1'd0, _zz_when_ArraySlice_l158_268_2};
  assign _zz_when_ArraySlice_l158_268_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_268_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_268 = {1'd0, _zz_when_ArraySlice_l159_268_1};
  assign _zz_when_ArraySlice_l159_268_2 = (_zz_when_ArraySlice_l159_268_3 - _zz_when_ArraySlice_l159_268_4);
  assign _zz_when_ArraySlice_l159_268_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_268_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_268_5);
  assign _zz_when_ArraySlice_l159_268_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_268_5 = {1'd0, _zz_when_ArraySlice_l159_268_6};
  assign _zz__zz_realValue_0_268 = {1'd0, wReg};
  assign _zz__zz_realValue_0_268_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_268_1 = (_zz_realValue_0_268_2 + _zz_realValue_0_268_3);
  assign _zz_realValue_0_268_2 = {1'd0, wReg};
  assign _zz_realValue_0_268_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_268_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_268 = {1'd0, _zz_when_ArraySlice_l166_268_1};
  assign _zz_when_ArraySlice_l166_268_2 = (_zz_when_ArraySlice_l166_268_3 + _zz_when_ArraySlice_l166_268_7);
  assign _zz_when_ArraySlice_l166_268_3 = (realValue_0_268 - _zz_when_ArraySlice_l166_268_4);
  assign _zz_when_ArraySlice_l166_268_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_268_5);
  assign _zz_when_ArraySlice_l166_268_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_268_5 = {1'd0, _zz_when_ArraySlice_l166_268_6};
  assign _zz_when_ArraySlice_l166_268_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_269 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_269_1);
  assign _zz_when_ArraySlice_l158_269_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_269_1 = {1'd0, _zz_when_ArraySlice_l158_269_2};
  assign _zz_when_ArraySlice_l158_269_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_269_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_269 = {2'd0, _zz_when_ArraySlice_l159_269_1};
  assign _zz_when_ArraySlice_l159_269_2 = (_zz_when_ArraySlice_l159_269_3 - _zz_when_ArraySlice_l159_269_4);
  assign _zz_when_ArraySlice_l159_269_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_269_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_269_5);
  assign _zz_when_ArraySlice_l159_269_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_269_5 = {1'd0, _zz_when_ArraySlice_l159_269_6};
  assign _zz__zz_realValue_0_269 = {1'd0, wReg};
  assign _zz__zz_realValue_0_269_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_269_1 = (_zz_realValue_0_269_2 + _zz_realValue_0_269_3);
  assign _zz_realValue_0_269_2 = {1'd0, wReg};
  assign _zz_realValue_0_269_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_269_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_269 = {2'd0, _zz_when_ArraySlice_l166_269_1};
  assign _zz_when_ArraySlice_l166_269_2 = (_zz_when_ArraySlice_l166_269_3 + _zz_when_ArraySlice_l166_269_7);
  assign _zz_when_ArraySlice_l166_269_3 = (realValue_0_269 - _zz_when_ArraySlice_l166_269_4);
  assign _zz_when_ArraySlice_l166_269_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_269_5);
  assign _zz_when_ArraySlice_l166_269_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_269_5 = {1'd0, _zz_when_ArraySlice_l166_269_6};
  assign _zz_when_ArraySlice_l166_269_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_270 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_270_1);
  assign _zz_when_ArraySlice_l158_270_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_270_1 = {1'd0, _zz_when_ArraySlice_l158_270_2};
  assign _zz_when_ArraySlice_l158_270_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_270_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_270 = {2'd0, _zz_when_ArraySlice_l159_270_1};
  assign _zz_when_ArraySlice_l159_270_2 = (_zz_when_ArraySlice_l159_270_3 - _zz_when_ArraySlice_l159_270_4);
  assign _zz_when_ArraySlice_l159_270_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_270_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_270_5);
  assign _zz_when_ArraySlice_l159_270_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_270_5 = {1'd0, _zz_when_ArraySlice_l159_270_6};
  assign _zz__zz_realValue_0_270 = {1'd0, wReg};
  assign _zz__zz_realValue_0_270_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_270_1 = (_zz_realValue_0_270_2 + _zz_realValue_0_270_3);
  assign _zz_realValue_0_270_2 = {1'd0, wReg};
  assign _zz_realValue_0_270_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_270_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_270 = {2'd0, _zz_when_ArraySlice_l166_270_1};
  assign _zz_when_ArraySlice_l166_270_2 = (_zz_when_ArraySlice_l166_270_3 + _zz_when_ArraySlice_l166_270_7);
  assign _zz_when_ArraySlice_l166_270_3 = (realValue_0_270 - _zz_when_ArraySlice_l166_270_4);
  assign _zz_when_ArraySlice_l166_270_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_270_5);
  assign _zz_when_ArraySlice_l166_270_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_270_5 = {1'd0, _zz_when_ArraySlice_l166_270_6};
  assign _zz_when_ArraySlice_l166_270_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_271 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_271_1);
  assign _zz_when_ArraySlice_l158_271_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_271_1 = {1'd0, _zz_when_ArraySlice_l158_271_2};
  assign _zz_when_ArraySlice_l158_271_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_271_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_271 = {3'd0, _zz_when_ArraySlice_l159_271_1};
  assign _zz_when_ArraySlice_l159_271_2 = (_zz_when_ArraySlice_l159_271_3 - _zz_when_ArraySlice_l159_271_4);
  assign _zz_when_ArraySlice_l159_271_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_271_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_271_5);
  assign _zz_when_ArraySlice_l159_271_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_271_5 = {1'd0, _zz_when_ArraySlice_l159_271_6};
  assign _zz__zz_realValue_0_271 = {1'd0, wReg};
  assign _zz__zz_realValue_0_271_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_271_1 = (_zz_realValue_0_271_2 + _zz_realValue_0_271_3);
  assign _zz_realValue_0_271_2 = {1'd0, wReg};
  assign _zz_realValue_0_271_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_271_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_271 = {3'd0, _zz_when_ArraySlice_l166_271_1};
  assign _zz_when_ArraySlice_l166_271_2 = (_zz_when_ArraySlice_l166_271_3 + _zz_when_ArraySlice_l166_271_7);
  assign _zz_when_ArraySlice_l166_271_3 = (realValue_0_271 - _zz_when_ArraySlice_l166_271_4);
  assign _zz_when_ArraySlice_l166_271_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_271_5);
  assign _zz_when_ArraySlice_l166_271_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_271_5 = {1'd0, _zz_when_ArraySlice_l166_271_6};
  assign _zz_when_ArraySlice_l166_271_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_2_2 = (_zz_when_ArraySlice_l285_2_3 + _zz_when_ArraySlice_l285_2_7);
  assign _zz_when_ArraySlice_l285_2_3 = (_zz_when_ArraySlice_l285_2_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_2_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l285_2_5);
  assign _zz_when_ArraySlice_l285_2_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_2_5 = {1'd0, _zz_when_ArraySlice_l285_2_6};
  assign _zz_when_ArraySlice_l285_2_8 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l285_2_7 = {2'd0, _zz_when_ArraySlice_l285_2_8};
  assign _zz_when_ArraySlice_l288_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_2_2 = (_zz_when_ArraySlice_l288_2_3 + 8'h01);
  assign _zz_when_ArraySlice_l288_2_3 = (selectReadFifo_2 + _zz_when_ArraySlice_l288_2_4);
  assign _zz_when_ArraySlice_l288_2_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_2_4 = {1'd0, _zz_when_ArraySlice_l288_2_5};
  assign _zz_selectReadFifo_2_27 = (selectReadFifo_2 + _zz_selectReadFifo_2_28);
  assign _zz_selectReadFifo_2_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_2_28 = {1'd0, _zz_selectReadFifo_2_29};
  assign _zz_when_ArraySlice_l295_2 = (_zz_when_ArraySlice_l295_2_1 % aReg);
  assign _zz_when_ArraySlice_l295_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_2_2 = (_zz_when_ArraySlice_l306_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l306_2_1 = {5'd0, _zz_when_ArraySlice_l306_2_2};
  assign _zz_when_ArraySlice_l306_2_3 = (bReg * aReg);
  assign _zz__zz_realValue1_0_32 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_32_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_32_1 = (_zz_realValue1_0_32_2 + _zz_realValue1_0_32_3);
  assign _zz_realValue1_0_32_2 = {1'd0, hReg};
  assign _zz_realValue1_0_32_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_2_2 = (outSliceNumb_2_value + 7'h01);
  assign _zz_when_ArraySlice_l307_2_1 = {1'd0, _zz_when_ArraySlice_l307_2_2};
  assign _zz_when_ArraySlice_l307_2_3 = (realValue1_0_32 / aReg);
  assign _zz_selectReadFifo_2_30 = (selectReadFifo_2 - _zz_selectReadFifo_2_31);
  assign _zz_selectReadFifo_2_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_272 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_272_1);
  assign _zz_when_ArraySlice_l158_272_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_272_1 = {4'd0, _zz_when_ArraySlice_l158_272_2};
  assign _zz_when_ArraySlice_l158_272_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_272 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_272_1 = (_zz_when_ArraySlice_l159_272_2 - _zz_when_ArraySlice_l159_272_3);
  assign _zz_when_ArraySlice_l159_272_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_272_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_272_4);
  assign _zz_when_ArraySlice_l159_272_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_272_4 = {4'd0, _zz_when_ArraySlice_l159_272_5};
  assign _zz__zz_realValue_0_272 = {1'd0, wReg};
  assign _zz__zz_realValue_0_272_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_272_1 = (_zz_realValue_0_272_2 + _zz_realValue_0_272_3);
  assign _zz_realValue_0_272_2 = {1'd0, wReg};
  assign _zz_realValue_0_272_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_272 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_272_1 = (_zz_when_ArraySlice_l166_272_2 + _zz_when_ArraySlice_l166_272_6);
  assign _zz_when_ArraySlice_l166_272_2 = (realValue_0_272 - _zz_when_ArraySlice_l166_272_3);
  assign _zz_when_ArraySlice_l166_272_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_272_4);
  assign _zz_when_ArraySlice_l166_272_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_272_4 = {4'd0, _zz_when_ArraySlice_l166_272_5};
  assign _zz_when_ArraySlice_l166_272_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_273 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_273_1);
  assign _zz_when_ArraySlice_l158_273_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_273_1 = {3'd0, _zz_when_ArraySlice_l158_273_2};
  assign _zz_when_ArraySlice_l158_273_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_273_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_273 = {1'd0, _zz_when_ArraySlice_l159_273_1};
  assign _zz_when_ArraySlice_l159_273_2 = (_zz_when_ArraySlice_l159_273_3 - _zz_when_ArraySlice_l159_273_4);
  assign _zz_when_ArraySlice_l159_273_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_273_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_273_5);
  assign _zz_when_ArraySlice_l159_273_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_273_5 = {3'd0, _zz_when_ArraySlice_l159_273_6};
  assign _zz__zz_realValue_0_273 = {1'd0, wReg};
  assign _zz__zz_realValue_0_273_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_273_1 = (_zz_realValue_0_273_2 + _zz_realValue_0_273_3);
  assign _zz_realValue_0_273_2 = {1'd0, wReg};
  assign _zz_realValue_0_273_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_273_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_273 = {1'd0, _zz_when_ArraySlice_l166_273_1};
  assign _zz_when_ArraySlice_l166_273_2 = (_zz_when_ArraySlice_l166_273_3 + _zz_when_ArraySlice_l166_273_7);
  assign _zz_when_ArraySlice_l166_273_3 = (realValue_0_273 - _zz_when_ArraySlice_l166_273_4);
  assign _zz_when_ArraySlice_l166_273_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_273_5);
  assign _zz_when_ArraySlice_l166_273_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_273_5 = {3'd0, _zz_when_ArraySlice_l166_273_6};
  assign _zz_when_ArraySlice_l166_273_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_274 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_274_1);
  assign _zz_when_ArraySlice_l158_274_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_274_1 = {2'd0, _zz_when_ArraySlice_l158_274_2};
  assign _zz_when_ArraySlice_l158_274_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_274_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_274 = {1'd0, _zz_when_ArraySlice_l159_274_1};
  assign _zz_when_ArraySlice_l159_274_2 = (_zz_when_ArraySlice_l159_274_3 - _zz_when_ArraySlice_l159_274_4);
  assign _zz_when_ArraySlice_l159_274_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_274_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_274_5);
  assign _zz_when_ArraySlice_l159_274_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_274_5 = {2'd0, _zz_when_ArraySlice_l159_274_6};
  assign _zz__zz_realValue_0_274 = {1'd0, wReg};
  assign _zz__zz_realValue_0_274_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_274_1 = (_zz_realValue_0_274_2 + _zz_realValue_0_274_3);
  assign _zz_realValue_0_274_2 = {1'd0, wReg};
  assign _zz_realValue_0_274_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_274_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_274 = {1'd0, _zz_when_ArraySlice_l166_274_1};
  assign _zz_when_ArraySlice_l166_274_2 = (_zz_when_ArraySlice_l166_274_3 + _zz_when_ArraySlice_l166_274_7);
  assign _zz_when_ArraySlice_l166_274_3 = (realValue_0_274 - _zz_when_ArraySlice_l166_274_4);
  assign _zz_when_ArraySlice_l166_274_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_274_5);
  assign _zz_when_ArraySlice_l166_274_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_274_5 = {2'd0, _zz_when_ArraySlice_l166_274_6};
  assign _zz_when_ArraySlice_l166_274_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_275 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_275_1);
  assign _zz_when_ArraySlice_l158_275_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_275_1 = {2'd0, _zz_when_ArraySlice_l158_275_2};
  assign _zz_when_ArraySlice_l158_275_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_275_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_275 = {1'd0, _zz_when_ArraySlice_l159_275_1};
  assign _zz_when_ArraySlice_l159_275_2 = (_zz_when_ArraySlice_l159_275_3 - _zz_when_ArraySlice_l159_275_4);
  assign _zz_when_ArraySlice_l159_275_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_275_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_275_5);
  assign _zz_when_ArraySlice_l159_275_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_275_5 = {2'd0, _zz_when_ArraySlice_l159_275_6};
  assign _zz__zz_realValue_0_275 = {1'd0, wReg};
  assign _zz__zz_realValue_0_275_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_275_1 = (_zz_realValue_0_275_2 + _zz_realValue_0_275_3);
  assign _zz_realValue_0_275_2 = {1'd0, wReg};
  assign _zz_realValue_0_275_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_275_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_275 = {1'd0, _zz_when_ArraySlice_l166_275_1};
  assign _zz_when_ArraySlice_l166_275_2 = (_zz_when_ArraySlice_l166_275_3 + _zz_when_ArraySlice_l166_275_7);
  assign _zz_when_ArraySlice_l166_275_3 = (realValue_0_275 - _zz_when_ArraySlice_l166_275_4);
  assign _zz_when_ArraySlice_l166_275_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_275_5);
  assign _zz_when_ArraySlice_l166_275_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_275_5 = {2'd0, _zz_when_ArraySlice_l166_275_6};
  assign _zz_when_ArraySlice_l166_275_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_276 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_276_1);
  assign _zz_when_ArraySlice_l158_276_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_276_1 = {1'd0, _zz_when_ArraySlice_l158_276_2};
  assign _zz_when_ArraySlice_l158_276_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_276_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_276 = {1'd0, _zz_when_ArraySlice_l159_276_1};
  assign _zz_when_ArraySlice_l159_276_2 = (_zz_when_ArraySlice_l159_276_3 - _zz_when_ArraySlice_l159_276_4);
  assign _zz_when_ArraySlice_l159_276_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_276_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_276_5);
  assign _zz_when_ArraySlice_l159_276_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_276_5 = {1'd0, _zz_when_ArraySlice_l159_276_6};
  assign _zz__zz_realValue_0_276 = {1'd0, wReg};
  assign _zz__zz_realValue_0_276_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_276_1 = (_zz_realValue_0_276_2 + _zz_realValue_0_276_3);
  assign _zz_realValue_0_276_2 = {1'd0, wReg};
  assign _zz_realValue_0_276_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_276_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_276 = {1'd0, _zz_when_ArraySlice_l166_276_1};
  assign _zz_when_ArraySlice_l166_276_2 = (_zz_when_ArraySlice_l166_276_3 + _zz_when_ArraySlice_l166_276_7);
  assign _zz_when_ArraySlice_l166_276_3 = (realValue_0_276 - _zz_when_ArraySlice_l166_276_4);
  assign _zz_when_ArraySlice_l166_276_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_276_5);
  assign _zz_when_ArraySlice_l166_276_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_276_5 = {1'd0, _zz_when_ArraySlice_l166_276_6};
  assign _zz_when_ArraySlice_l166_276_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_277 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_277_1);
  assign _zz_when_ArraySlice_l158_277_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_277_1 = {1'd0, _zz_when_ArraySlice_l158_277_2};
  assign _zz_when_ArraySlice_l158_277_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_277_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_277 = {2'd0, _zz_when_ArraySlice_l159_277_1};
  assign _zz_when_ArraySlice_l159_277_2 = (_zz_when_ArraySlice_l159_277_3 - _zz_when_ArraySlice_l159_277_4);
  assign _zz_when_ArraySlice_l159_277_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_277_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_277_5);
  assign _zz_when_ArraySlice_l159_277_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_277_5 = {1'd0, _zz_when_ArraySlice_l159_277_6};
  assign _zz__zz_realValue_0_277 = {1'd0, wReg};
  assign _zz__zz_realValue_0_277_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_277_1 = (_zz_realValue_0_277_2 + _zz_realValue_0_277_3);
  assign _zz_realValue_0_277_2 = {1'd0, wReg};
  assign _zz_realValue_0_277_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_277_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_277 = {2'd0, _zz_when_ArraySlice_l166_277_1};
  assign _zz_when_ArraySlice_l166_277_2 = (_zz_when_ArraySlice_l166_277_3 + _zz_when_ArraySlice_l166_277_7);
  assign _zz_when_ArraySlice_l166_277_3 = (realValue_0_277 - _zz_when_ArraySlice_l166_277_4);
  assign _zz_when_ArraySlice_l166_277_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_277_5);
  assign _zz_when_ArraySlice_l166_277_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_277_5 = {1'd0, _zz_when_ArraySlice_l166_277_6};
  assign _zz_when_ArraySlice_l166_277_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_278 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_278_1);
  assign _zz_when_ArraySlice_l158_278_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_278_1 = {1'd0, _zz_when_ArraySlice_l158_278_2};
  assign _zz_when_ArraySlice_l158_278_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_278_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_278 = {2'd0, _zz_when_ArraySlice_l159_278_1};
  assign _zz_when_ArraySlice_l159_278_2 = (_zz_when_ArraySlice_l159_278_3 - _zz_when_ArraySlice_l159_278_4);
  assign _zz_when_ArraySlice_l159_278_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_278_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_278_5);
  assign _zz_when_ArraySlice_l159_278_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_278_5 = {1'd0, _zz_when_ArraySlice_l159_278_6};
  assign _zz__zz_realValue_0_278 = {1'd0, wReg};
  assign _zz__zz_realValue_0_278_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_278_1 = (_zz_realValue_0_278_2 + _zz_realValue_0_278_3);
  assign _zz_realValue_0_278_2 = {1'd0, wReg};
  assign _zz_realValue_0_278_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_278_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_278 = {2'd0, _zz_when_ArraySlice_l166_278_1};
  assign _zz_when_ArraySlice_l166_278_2 = (_zz_when_ArraySlice_l166_278_3 + _zz_when_ArraySlice_l166_278_7);
  assign _zz_when_ArraySlice_l166_278_3 = (realValue_0_278 - _zz_when_ArraySlice_l166_278_4);
  assign _zz_when_ArraySlice_l166_278_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_278_5);
  assign _zz_when_ArraySlice_l166_278_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_278_5 = {1'd0, _zz_when_ArraySlice_l166_278_6};
  assign _zz_when_ArraySlice_l166_278_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_279 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_279_1);
  assign _zz_when_ArraySlice_l158_279_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_279_1 = {1'd0, _zz_when_ArraySlice_l158_279_2};
  assign _zz_when_ArraySlice_l158_279_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_279_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_279 = {3'd0, _zz_when_ArraySlice_l159_279_1};
  assign _zz_when_ArraySlice_l159_279_2 = (_zz_when_ArraySlice_l159_279_3 - _zz_when_ArraySlice_l159_279_4);
  assign _zz_when_ArraySlice_l159_279_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_279_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_279_5);
  assign _zz_when_ArraySlice_l159_279_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_279_5 = {1'd0, _zz_when_ArraySlice_l159_279_6};
  assign _zz__zz_realValue_0_279 = {1'd0, wReg};
  assign _zz__zz_realValue_0_279_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_279_1 = (_zz_realValue_0_279_2 + _zz_realValue_0_279_3);
  assign _zz_realValue_0_279_2 = {1'd0, wReg};
  assign _zz_realValue_0_279_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_279_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_279 = {3'd0, _zz_when_ArraySlice_l166_279_1};
  assign _zz_when_ArraySlice_l166_279_2 = (_zz_when_ArraySlice_l166_279_3 + _zz_when_ArraySlice_l166_279_7);
  assign _zz_when_ArraySlice_l166_279_3 = (realValue_0_279 - _zz_when_ArraySlice_l166_279_4);
  assign _zz_when_ArraySlice_l166_279_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_279_5);
  assign _zz_when_ArraySlice_l166_279_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_279_5 = {1'd0, _zz_when_ArraySlice_l166_279_6};
  assign _zz_when_ArraySlice_l166_279_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_2 = (_zz_when_ArraySlice_l318_2_1 % aReg);
  assign _zz_when_ArraySlice_l318_2_1 = (handshakeTimes_2_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_2_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_2_2 = (selectReadFifo_2 + _zz_when_ArraySlice_l304_2_3);
  assign _zz_when_ArraySlice_l304_2_4 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l304_2_3 = {2'd0, _zz_when_ArraySlice_l304_2_4};
  assign _zz_when_ArraySlice_l325_2_2 = (_zz_when_ArraySlice_l325_2_3 - 8'h01);
  assign _zz_when_ArraySlice_l325_2_1 = {5'd0, _zz_when_ArraySlice_l325_2_2};
  assign _zz_when_ArraySlice_l325_2_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_3_1 = (selectReadFifo_3 + _zz_when_ArraySlice_l233_3_2);
  assign _zz_when_ArraySlice_l233_3_3 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l233_3_2 = {2'd0, _zz_when_ArraySlice_l233_3_3};
  assign _zz_when_ArraySlice_l233_3_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l234_3_4);
  assign _zz_when_ArraySlice_l234_3_2 = _zz_when_ArraySlice_l234_3_3[6:0];
  assign _zz_when_ArraySlice_l234_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l234_3_4 = {2'd0, _zz_when_ArraySlice_l234_3_5};
  assign _zz__zz_outputStreamArrayData_3_valid_1_2 = (bReg * 2'b11);
  assign _zz__zz_outputStreamArrayData_3_valid_1_1 = {2'd0, _zz__zz_outputStreamArrayData_3_valid_1_2};
  assign _zz__zz_14 = _zz_outputStreamArrayData_3_valid_1[6:0];
  assign _zz_outputStreamArrayData_3_valid_5 = _zz_outputStreamArrayData_3_valid_1[6:0];
  assign _zz_outputStreamArrayData_3_payload_3 = _zz_outputStreamArrayData_3_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l240_3_4);
  assign _zz_when_ArraySlice_l240_3_2 = _zz_when_ArraySlice_l240_3_3[6:0];
  assign _zz_when_ArraySlice_l240_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l240_3_4 = {2'd0, _zz_when_ArraySlice_l240_3_5};
  assign _zz_when_ArraySlice_l241_3_1 = (_zz_when_ArraySlice_l241_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l241_3 = {5'd0, _zz_when_ArraySlice_l241_3_1};
  assign _zz_when_ArraySlice_l241_3_2 = (bReg * aReg);
  assign _zz_selectReadFifo_3_16 = (selectReadFifo_3 - _zz_selectReadFifo_3_17);
  assign _zz_selectReadFifo_3_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_3 = (_zz_when_ArraySlice_l244_3_1 % aReg);
  assign _zz_when_ArraySlice_l244_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l249_3_4);
  assign _zz_when_ArraySlice_l249_3_2 = _zz_when_ArraySlice_l249_3_3[6:0];
  assign _zz_when_ArraySlice_l249_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l249_3_4 = {2'd0, _zz_when_ArraySlice_l249_3_5};
  assign _zz_when_ArraySlice_l250_3_1 = (_zz_when_ArraySlice_l250_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l250_3 = {5'd0, _zz_when_ArraySlice_l250_3_1};
  assign _zz_when_ArraySlice_l250_3_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_33 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_33_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_33_1 = (_zz_realValue1_0_33_2 + _zz_realValue1_0_33_3);
  assign _zz_realValue1_0_33_2 = {1'd0, hReg};
  assign _zz_realValue1_0_33_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l252_3 = {1'd0, _zz_when_ArraySlice_l252_3_1};
  assign _zz_when_ArraySlice_l252_3_2 = (realValue1_0_33 / aReg);
  assign _zz_selectReadFifo_3_18 = (selectReadFifo_3 - _zz_selectReadFifo_3_19);
  assign _zz_selectReadFifo_3_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_3_21 = 1'b1;
  assign _zz_selectReadFifo_3_20 = {7'd0, _zz_selectReadFifo_3_21};
  assign _zz_when_ArraySlice_l158_280 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_280_1);
  assign _zz_when_ArraySlice_l158_280_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_280_1 = {4'd0, _zz_when_ArraySlice_l158_280_2};
  assign _zz_when_ArraySlice_l158_280_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_280 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_280_1 = (_zz_when_ArraySlice_l159_280_2 - _zz_when_ArraySlice_l159_280_3);
  assign _zz_when_ArraySlice_l159_280_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_280_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_280_4);
  assign _zz_when_ArraySlice_l159_280_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_280_4 = {4'd0, _zz_when_ArraySlice_l159_280_5};
  assign _zz__zz_realValue_0_280 = {1'd0, wReg};
  assign _zz__zz_realValue_0_280_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_280_1 = (_zz_realValue_0_280_2 + _zz_realValue_0_280_3);
  assign _zz_realValue_0_280_2 = {1'd0, wReg};
  assign _zz_realValue_0_280_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_280 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_280_1 = (_zz_when_ArraySlice_l166_280_2 + _zz_when_ArraySlice_l166_280_6);
  assign _zz_when_ArraySlice_l166_280_2 = (realValue_0_280 - _zz_when_ArraySlice_l166_280_3);
  assign _zz_when_ArraySlice_l166_280_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_280_4);
  assign _zz_when_ArraySlice_l166_280_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_280_4 = {4'd0, _zz_when_ArraySlice_l166_280_5};
  assign _zz_when_ArraySlice_l166_280_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_281 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_281_1);
  assign _zz_when_ArraySlice_l158_281_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_281_1 = {3'd0, _zz_when_ArraySlice_l158_281_2};
  assign _zz_when_ArraySlice_l158_281_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_281_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_281 = {1'd0, _zz_when_ArraySlice_l159_281_1};
  assign _zz_when_ArraySlice_l159_281_2 = (_zz_when_ArraySlice_l159_281_3 - _zz_when_ArraySlice_l159_281_4);
  assign _zz_when_ArraySlice_l159_281_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_281_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_281_5);
  assign _zz_when_ArraySlice_l159_281_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_281_5 = {3'd0, _zz_when_ArraySlice_l159_281_6};
  assign _zz__zz_realValue_0_281 = {1'd0, wReg};
  assign _zz__zz_realValue_0_281_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_281_1 = (_zz_realValue_0_281_2 + _zz_realValue_0_281_3);
  assign _zz_realValue_0_281_2 = {1'd0, wReg};
  assign _zz_realValue_0_281_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_281_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_281 = {1'd0, _zz_when_ArraySlice_l166_281_1};
  assign _zz_when_ArraySlice_l166_281_2 = (_zz_when_ArraySlice_l166_281_3 + _zz_when_ArraySlice_l166_281_7);
  assign _zz_when_ArraySlice_l166_281_3 = (realValue_0_281 - _zz_when_ArraySlice_l166_281_4);
  assign _zz_when_ArraySlice_l166_281_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_281_5);
  assign _zz_when_ArraySlice_l166_281_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_281_5 = {3'd0, _zz_when_ArraySlice_l166_281_6};
  assign _zz_when_ArraySlice_l166_281_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_282 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_282_1);
  assign _zz_when_ArraySlice_l158_282_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_282_1 = {2'd0, _zz_when_ArraySlice_l158_282_2};
  assign _zz_when_ArraySlice_l158_282_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_282_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_282 = {1'd0, _zz_when_ArraySlice_l159_282_1};
  assign _zz_when_ArraySlice_l159_282_2 = (_zz_when_ArraySlice_l159_282_3 - _zz_when_ArraySlice_l159_282_4);
  assign _zz_when_ArraySlice_l159_282_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_282_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_282_5);
  assign _zz_when_ArraySlice_l159_282_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_282_5 = {2'd0, _zz_when_ArraySlice_l159_282_6};
  assign _zz__zz_realValue_0_282 = {1'd0, wReg};
  assign _zz__zz_realValue_0_282_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_282_1 = (_zz_realValue_0_282_2 + _zz_realValue_0_282_3);
  assign _zz_realValue_0_282_2 = {1'd0, wReg};
  assign _zz_realValue_0_282_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_282_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_282 = {1'd0, _zz_when_ArraySlice_l166_282_1};
  assign _zz_when_ArraySlice_l166_282_2 = (_zz_when_ArraySlice_l166_282_3 + _zz_when_ArraySlice_l166_282_7);
  assign _zz_when_ArraySlice_l166_282_3 = (realValue_0_282 - _zz_when_ArraySlice_l166_282_4);
  assign _zz_when_ArraySlice_l166_282_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_282_5);
  assign _zz_when_ArraySlice_l166_282_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_282_5 = {2'd0, _zz_when_ArraySlice_l166_282_6};
  assign _zz_when_ArraySlice_l166_282_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_283 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_283_1);
  assign _zz_when_ArraySlice_l158_283_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_283_1 = {2'd0, _zz_when_ArraySlice_l158_283_2};
  assign _zz_when_ArraySlice_l158_283_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_283_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_283 = {1'd0, _zz_when_ArraySlice_l159_283_1};
  assign _zz_when_ArraySlice_l159_283_2 = (_zz_when_ArraySlice_l159_283_3 - _zz_when_ArraySlice_l159_283_4);
  assign _zz_when_ArraySlice_l159_283_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_283_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_283_5);
  assign _zz_when_ArraySlice_l159_283_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_283_5 = {2'd0, _zz_when_ArraySlice_l159_283_6};
  assign _zz__zz_realValue_0_283 = {1'd0, wReg};
  assign _zz__zz_realValue_0_283_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_283_1 = (_zz_realValue_0_283_2 + _zz_realValue_0_283_3);
  assign _zz_realValue_0_283_2 = {1'd0, wReg};
  assign _zz_realValue_0_283_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_283_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_283 = {1'd0, _zz_when_ArraySlice_l166_283_1};
  assign _zz_when_ArraySlice_l166_283_2 = (_zz_when_ArraySlice_l166_283_3 + _zz_when_ArraySlice_l166_283_7);
  assign _zz_when_ArraySlice_l166_283_3 = (realValue_0_283 - _zz_when_ArraySlice_l166_283_4);
  assign _zz_when_ArraySlice_l166_283_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_283_5);
  assign _zz_when_ArraySlice_l166_283_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_283_5 = {2'd0, _zz_when_ArraySlice_l166_283_6};
  assign _zz_when_ArraySlice_l166_283_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_284 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_284_1);
  assign _zz_when_ArraySlice_l158_284_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_284_1 = {1'd0, _zz_when_ArraySlice_l158_284_2};
  assign _zz_when_ArraySlice_l158_284_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_284_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_284 = {1'd0, _zz_when_ArraySlice_l159_284_1};
  assign _zz_when_ArraySlice_l159_284_2 = (_zz_when_ArraySlice_l159_284_3 - _zz_when_ArraySlice_l159_284_4);
  assign _zz_when_ArraySlice_l159_284_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_284_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_284_5);
  assign _zz_when_ArraySlice_l159_284_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_284_5 = {1'd0, _zz_when_ArraySlice_l159_284_6};
  assign _zz__zz_realValue_0_284 = {1'd0, wReg};
  assign _zz__zz_realValue_0_284_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_284_1 = (_zz_realValue_0_284_2 + _zz_realValue_0_284_3);
  assign _zz_realValue_0_284_2 = {1'd0, wReg};
  assign _zz_realValue_0_284_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_284_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_284 = {1'd0, _zz_when_ArraySlice_l166_284_1};
  assign _zz_when_ArraySlice_l166_284_2 = (_zz_when_ArraySlice_l166_284_3 + _zz_when_ArraySlice_l166_284_7);
  assign _zz_when_ArraySlice_l166_284_3 = (realValue_0_284 - _zz_when_ArraySlice_l166_284_4);
  assign _zz_when_ArraySlice_l166_284_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_284_5);
  assign _zz_when_ArraySlice_l166_284_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_284_5 = {1'd0, _zz_when_ArraySlice_l166_284_6};
  assign _zz_when_ArraySlice_l166_284_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_285 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_285_1);
  assign _zz_when_ArraySlice_l158_285_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_285_1 = {1'd0, _zz_when_ArraySlice_l158_285_2};
  assign _zz_when_ArraySlice_l158_285_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_285_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_285 = {2'd0, _zz_when_ArraySlice_l159_285_1};
  assign _zz_when_ArraySlice_l159_285_2 = (_zz_when_ArraySlice_l159_285_3 - _zz_when_ArraySlice_l159_285_4);
  assign _zz_when_ArraySlice_l159_285_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_285_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_285_5);
  assign _zz_when_ArraySlice_l159_285_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_285_5 = {1'd0, _zz_when_ArraySlice_l159_285_6};
  assign _zz__zz_realValue_0_285 = {1'd0, wReg};
  assign _zz__zz_realValue_0_285_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_285_1 = (_zz_realValue_0_285_2 + _zz_realValue_0_285_3);
  assign _zz_realValue_0_285_2 = {1'd0, wReg};
  assign _zz_realValue_0_285_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_285_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_285 = {2'd0, _zz_when_ArraySlice_l166_285_1};
  assign _zz_when_ArraySlice_l166_285_2 = (_zz_when_ArraySlice_l166_285_3 + _zz_when_ArraySlice_l166_285_7);
  assign _zz_when_ArraySlice_l166_285_3 = (realValue_0_285 - _zz_when_ArraySlice_l166_285_4);
  assign _zz_when_ArraySlice_l166_285_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_285_5);
  assign _zz_when_ArraySlice_l166_285_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_285_5 = {1'd0, _zz_when_ArraySlice_l166_285_6};
  assign _zz_when_ArraySlice_l166_285_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_286 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_286_1);
  assign _zz_when_ArraySlice_l158_286_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_286_1 = {1'd0, _zz_when_ArraySlice_l158_286_2};
  assign _zz_when_ArraySlice_l158_286_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_286_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_286 = {2'd0, _zz_when_ArraySlice_l159_286_1};
  assign _zz_when_ArraySlice_l159_286_2 = (_zz_when_ArraySlice_l159_286_3 - _zz_when_ArraySlice_l159_286_4);
  assign _zz_when_ArraySlice_l159_286_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_286_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_286_5);
  assign _zz_when_ArraySlice_l159_286_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_286_5 = {1'd0, _zz_when_ArraySlice_l159_286_6};
  assign _zz__zz_realValue_0_286 = {1'd0, wReg};
  assign _zz__zz_realValue_0_286_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_286_1 = (_zz_realValue_0_286_2 + _zz_realValue_0_286_3);
  assign _zz_realValue_0_286_2 = {1'd0, wReg};
  assign _zz_realValue_0_286_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_286_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_286 = {2'd0, _zz_when_ArraySlice_l166_286_1};
  assign _zz_when_ArraySlice_l166_286_2 = (_zz_when_ArraySlice_l166_286_3 + _zz_when_ArraySlice_l166_286_7);
  assign _zz_when_ArraySlice_l166_286_3 = (realValue_0_286 - _zz_when_ArraySlice_l166_286_4);
  assign _zz_when_ArraySlice_l166_286_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_286_5);
  assign _zz_when_ArraySlice_l166_286_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_286_5 = {1'd0, _zz_when_ArraySlice_l166_286_6};
  assign _zz_when_ArraySlice_l166_286_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_287 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_287_1);
  assign _zz_when_ArraySlice_l158_287_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_287_1 = {1'd0, _zz_when_ArraySlice_l158_287_2};
  assign _zz_when_ArraySlice_l158_287_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_287_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_287 = {3'd0, _zz_when_ArraySlice_l159_287_1};
  assign _zz_when_ArraySlice_l159_287_2 = (_zz_when_ArraySlice_l159_287_3 - _zz_when_ArraySlice_l159_287_4);
  assign _zz_when_ArraySlice_l159_287_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_287_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_287_5);
  assign _zz_when_ArraySlice_l159_287_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_287_5 = {1'd0, _zz_when_ArraySlice_l159_287_6};
  assign _zz__zz_realValue_0_287 = {1'd0, wReg};
  assign _zz__zz_realValue_0_287_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_287_1 = (_zz_realValue_0_287_2 + _zz_realValue_0_287_3);
  assign _zz_realValue_0_287_2 = {1'd0, wReg};
  assign _zz_realValue_0_287_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_287_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_287 = {3'd0, _zz_when_ArraySlice_l166_287_1};
  assign _zz_when_ArraySlice_l166_287_2 = (_zz_when_ArraySlice_l166_287_3 + _zz_when_ArraySlice_l166_287_7);
  assign _zz_when_ArraySlice_l166_287_3 = (realValue_0_287 - _zz_when_ArraySlice_l166_287_4);
  assign _zz_when_ArraySlice_l166_287_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_287_5);
  assign _zz_when_ArraySlice_l166_287_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_287_5 = {1'd0, _zz_when_ArraySlice_l166_287_6};
  assign _zz_when_ArraySlice_l166_287_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_3_2 = (_zz_when_ArraySlice_l260_3_3 + _zz_when_ArraySlice_l260_3_7);
  assign _zz_when_ArraySlice_l260_3_3 = (_zz_when_ArraySlice_l260_3_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l260_3_5);
  assign _zz_when_ArraySlice_l260_3_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_3_5 = {1'd0, _zz_when_ArraySlice_l260_3_6};
  assign _zz_when_ArraySlice_l260_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l260_3_7 = {2'd0, _zz_when_ArraySlice_l260_3_8};
  assign _zz_when_ArraySlice_l263_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_3_2 = (_zz_when_ArraySlice_l263_3_3 + 8'h01);
  assign _zz_when_ArraySlice_l263_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l263_3_4);
  assign _zz_when_ArraySlice_l263_3_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_3_4 = {1'd0, _zz_when_ArraySlice_l263_3_5};
  assign _zz_selectReadFifo_3_22 = (selectReadFifo_3 + _zz_selectReadFifo_3_23);
  assign _zz_selectReadFifo_3_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_23 = {1'd0, _zz_selectReadFifo_3_24};
  assign _zz_when_ArraySlice_l270_3 = (_zz_when_ArraySlice_l270_3_1 % aReg);
  assign _zz_when_ArraySlice_l270_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l274_3_4);
  assign _zz_when_ArraySlice_l274_3_2 = _zz_when_ArraySlice_l274_3_3[6:0];
  assign _zz_when_ArraySlice_l274_3_5 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l274_3_4 = {2'd0, _zz_when_ArraySlice_l274_3_5};
  assign _zz_when_ArraySlice_l275_3_2 = (_zz_when_ArraySlice_l275_3_3 - _zz_when_ArraySlice_l275_3_4);
  assign _zz_when_ArraySlice_l275_3_1 = {5'd0, _zz_when_ArraySlice_l275_3_2};
  assign _zz_when_ArraySlice_l275_3_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_3_5 = 1'b1;
  assign _zz_when_ArraySlice_l275_3_4 = {7'd0, _zz_when_ArraySlice_l275_3_5};
  assign _zz__zz_realValue1_0_34 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_34_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_34_1 = (_zz_realValue1_0_34_2 + _zz_realValue1_0_34_3);
  assign _zz_realValue1_0_34_2 = {1'd0, hReg};
  assign _zz_realValue1_0_34_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l277_3 = {1'd0, _zz_when_ArraySlice_l277_3_1};
  assign _zz_when_ArraySlice_l277_3_2 = (realValue1_0_34 / aReg);
  assign _zz_selectReadFifo_3_25 = (selectReadFifo_3 - _zz_selectReadFifo_3_26);
  assign _zz_selectReadFifo_3_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_288 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_288_1);
  assign _zz_when_ArraySlice_l158_288_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_288_1 = {4'd0, _zz_when_ArraySlice_l158_288_2};
  assign _zz_when_ArraySlice_l158_288_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_288 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_288_1 = (_zz_when_ArraySlice_l159_288_2 - _zz_when_ArraySlice_l159_288_3);
  assign _zz_when_ArraySlice_l159_288_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_288_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_288_4);
  assign _zz_when_ArraySlice_l159_288_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_288_4 = {4'd0, _zz_when_ArraySlice_l159_288_5};
  assign _zz__zz_realValue_0_288 = {1'd0, wReg};
  assign _zz__zz_realValue_0_288_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_288_1 = (_zz_realValue_0_288_2 + _zz_realValue_0_288_3);
  assign _zz_realValue_0_288_2 = {1'd0, wReg};
  assign _zz_realValue_0_288_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_288 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_288_1 = (_zz_when_ArraySlice_l166_288_2 + _zz_when_ArraySlice_l166_288_6);
  assign _zz_when_ArraySlice_l166_288_2 = (realValue_0_288 - _zz_when_ArraySlice_l166_288_3);
  assign _zz_when_ArraySlice_l166_288_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_288_4);
  assign _zz_when_ArraySlice_l166_288_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_288_4 = {4'd0, _zz_when_ArraySlice_l166_288_5};
  assign _zz_when_ArraySlice_l166_288_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_289 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_289_1);
  assign _zz_when_ArraySlice_l158_289_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_289_1 = {3'd0, _zz_when_ArraySlice_l158_289_2};
  assign _zz_when_ArraySlice_l158_289_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_289_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_289 = {1'd0, _zz_when_ArraySlice_l159_289_1};
  assign _zz_when_ArraySlice_l159_289_2 = (_zz_when_ArraySlice_l159_289_3 - _zz_when_ArraySlice_l159_289_4);
  assign _zz_when_ArraySlice_l159_289_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_289_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_289_5);
  assign _zz_when_ArraySlice_l159_289_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_289_5 = {3'd0, _zz_when_ArraySlice_l159_289_6};
  assign _zz__zz_realValue_0_289 = {1'd0, wReg};
  assign _zz__zz_realValue_0_289_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_289_1 = (_zz_realValue_0_289_2 + _zz_realValue_0_289_3);
  assign _zz_realValue_0_289_2 = {1'd0, wReg};
  assign _zz_realValue_0_289_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_289_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_289 = {1'd0, _zz_when_ArraySlice_l166_289_1};
  assign _zz_when_ArraySlice_l166_289_2 = (_zz_when_ArraySlice_l166_289_3 + _zz_when_ArraySlice_l166_289_7);
  assign _zz_when_ArraySlice_l166_289_3 = (realValue_0_289 - _zz_when_ArraySlice_l166_289_4);
  assign _zz_when_ArraySlice_l166_289_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_289_5);
  assign _zz_when_ArraySlice_l166_289_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_289_5 = {3'd0, _zz_when_ArraySlice_l166_289_6};
  assign _zz_when_ArraySlice_l166_289_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_290 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_290_1);
  assign _zz_when_ArraySlice_l158_290_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_290_1 = {2'd0, _zz_when_ArraySlice_l158_290_2};
  assign _zz_when_ArraySlice_l158_290_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_290_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_290 = {1'd0, _zz_when_ArraySlice_l159_290_1};
  assign _zz_when_ArraySlice_l159_290_2 = (_zz_when_ArraySlice_l159_290_3 - _zz_when_ArraySlice_l159_290_4);
  assign _zz_when_ArraySlice_l159_290_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_290_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_290_5);
  assign _zz_when_ArraySlice_l159_290_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_290_5 = {2'd0, _zz_when_ArraySlice_l159_290_6};
  assign _zz__zz_realValue_0_290 = {1'd0, wReg};
  assign _zz__zz_realValue_0_290_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_290_1 = (_zz_realValue_0_290_2 + _zz_realValue_0_290_3);
  assign _zz_realValue_0_290_2 = {1'd0, wReg};
  assign _zz_realValue_0_290_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_290_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_290 = {1'd0, _zz_when_ArraySlice_l166_290_1};
  assign _zz_when_ArraySlice_l166_290_2 = (_zz_when_ArraySlice_l166_290_3 + _zz_when_ArraySlice_l166_290_7);
  assign _zz_when_ArraySlice_l166_290_3 = (realValue_0_290 - _zz_when_ArraySlice_l166_290_4);
  assign _zz_when_ArraySlice_l166_290_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_290_5);
  assign _zz_when_ArraySlice_l166_290_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_290_5 = {2'd0, _zz_when_ArraySlice_l166_290_6};
  assign _zz_when_ArraySlice_l166_290_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_291 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_291_1);
  assign _zz_when_ArraySlice_l158_291_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_291_1 = {2'd0, _zz_when_ArraySlice_l158_291_2};
  assign _zz_when_ArraySlice_l158_291_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_291_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_291 = {1'd0, _zz_when_ArraySlice_l159_291_1};
  assign _zz_when_ArraySlice_l159_291_2 = (_zz_when_ArraySlice_l159_291_3 - _zz_when_ArraySlice_l159_291_4);
  assign _zz_when_ArraySlice_l159_291_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_291_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_291_5);
  assign _zz_when_ArraySlice_l159_291_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_291_5 = {2'd0, _zz_when_ArraySlice_l159_291_6};
  assign _zz__zz_realValue_0_291 = {1'd0, wReg};
  assign _zz__zz_realValue_0_291_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_291_1 = (_zz_realValue_0_291_2 + _zz_realValue_0_291_3);
  assign _zz_realValue_0_291_2 = {1'd0, wReg};
  assign _zz_realValue_0_291_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_291_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_291 = {1'd0, _zz_when_ArraySlice_l166_291_1};
  assign _zz_when_ArraySlice_l166_291_2 = (_zz_when_ArraySlice_l166_291_3 + _zz_when_ArraySlice_l166_291_7);
  assign _zz_when_ArraySlice_l166_291_3 = (realValue_0_291 - _zz_when_ArraySlice_l166_291_4);
  assign _zz_when_ArraySlice_l166_291_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_291_5);
  assign _zz_when_ArraySlice_l166_291_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_291_5 = {2'd0, _zz_when_ArraySlice_l166_291_6};
  assign _zz_when_ArraySlice_l166_291_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_292 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_292_1);
  assign _zz_when_ArraySlice_l158_292_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_292_1 = {1'd0, _zz_when_ArraySlice_l158_292_2};
  assign _zz_when_ArraySlice_l158_292_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_292_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_292 = {1'd0, _zz_when_ArraySlice_l159_292_1};
  assign _zz_when_ArraySlice_l159_292_2 = (_zz_when_ArraySlice_l159_292_3 - _zz_when_ArraySlice_l159_292_4);
  assign _zz_when_ArraySlice_l159_292_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_292_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_292_5);
  assign _zz_when_ArraySlice_l159_292_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_292_5 = {1'd0, _zz_when_ArraySlice_l159_292_6};
  assign _zz__zz_realValue_0_292 = {1'd0, wReg};
  assign _zz__zz_realValue_0_292_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_292_1 = (_zz_realValue_0_292_2 + _zz_realValue_0_292_3);
  assign _zz_realValue_0_292_2 = {1'd0, wReg};
  assign _zz_realValue_0_292_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_292_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_292 = {1'd0, _zz_when_ArraySlice_l166_292_1};
  assign _zz_when_ArraySlice_l166_292_2 = (_zz_when_ArraySlice_l166_292_3 + _zz_when_ArraySlice_l166_292_7);
  assign _zz_when_ArraySlice_l166_292_3 = (realValue_0_292 - _zz_when_ArraySlice_l166_292_4);
  assign _zz_when_ArraySlice_l166_292_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_292_5);
  assign _zz_when_ArraySlice_l166_292_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_292_5 = {1'd0, _zz_when_ArraySlice_l166_292_6};
  assign _zz_when_ArraySlice_l166_292_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_293 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_293_1);
  assign _zz_when_ArraySlice_l158_293_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_293_1 = {1'd0, _zz_when_ArraySlice_l158_293_2};
  assign _zz_when_ArraySlice_l158_293_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_293_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_293 = {2'd0, _zz_when_ArraySlice_l159_293_1};
  assign _zz_when_ArraySlice_l159_293_2 = (_zz_when_ArraySlice_l159_293_3 - _zz_when_ArraySlice_l159_293_4);
  assign _zz_when_ArraySlice_l159_293_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_293_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_293_5);
  assign _zz_when_ArraySlice_l159_293_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_293_5 = {1'd0, _zz_when_ArraySlice_l159_293_6};
  assign _zz__zz_realValue_0_293 = {1'd0, wReg};
  assign _zz__zz_realValue_0_293_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_293_1 = (_zz_realValue_0_293_2 + _zz_realValue_0_293_3);
  assign _zz_realValue_0_293_2 = {1'd0, wReg};
  assign _zz_realValue_0_293_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_293_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_293 = {2'd0, _zz_when_ArraySlice_l166_293_1};
  assign _zz_when_ArraySlice_l166_293_2 = (_zz_when_ArraySlice_l166_293_3 + _zz_when_ArraySlice_l166_293_7);
  assign _zz_when_ArraySlice_l166_293_3 = (realValue_0_293 - _zz_when_ArraySlice_l166_293_4);
  assign _zz_when_ArraySlice_l166_293_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_293_5);
  assign _zz_when_ArraySlice_l166_293_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_293_5 = {1'd0, _zz_when_ArraySlice_l166_293_6};
  assign _zz_when_ArraySlice_l166_293_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_294 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_294_1);
  assign _zz_when_ArraySlice_l158_294_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_294_1 = {1'd0, _zz_when_ArraySlice_l158_294_2};
  assign _zz_when_ArraySlice_l158_294_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_294_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_294 = {2'd0, _zz_when_ArraySlice_l159_294_1};
  assign _zz_when_ArraySlice_l159_294_2 = (_zz_when_ArraySlice_l159_294_3 - _zz_when_ArraySlice_l159_294_4);
  assign _zz_when_ArraySlice_l159_294_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_294_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_294_5);
  assign _zz_when_ArraySlice_l159_294_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_294_5 = {1'd0, _zz_when_ArraySlice_l159_294_6};
  assign _zz__zz_realValue_0_294 = {1'd0, wReg};
  assign _zz__zz_realValue_0_294_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_294_1 = (_zz_realValue_0_294_2 + _zz_realValue_0_294_3);
  assign _zz_realValue_0_294_2 = {1'd0, wReg};
  assign _zz_realValue_0_294_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_294_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_294 = {2'd0, _zz_when_ArraySlice_l166_294_1};
  assign _zz_when_ArraySlice_l166_294_2 = (_zz_when_ArraySlice_l166_294_3 + _zz_when_ArraySlice_l166_294_7);
  assign _zz_when_ArraySlice_l166_294_3 = (realValue_0_294 - _zz_when_ArraySlice_l166_294_4);
  assign _zz_when_ArraySlice_l166_294_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_294_5);
  assign _zz_when_ArraySlice_l166_294_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_294_5 = {1'd0, _zz_when_ArraySlice_l166_294_6};
  assign _zz_when_ArraySlice_l166_294_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_295 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_295_1);
  assign _zz_when_ArraySlice_l158_295_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_295_1 = {1'd0, _zz_when_ArraySlice_l158_295_2};
  assign _zz_when_ArraySlice_l158_295_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_295_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_295 = {3'd0, _zz_when_ArraySlice_l159_295_1};
  assign _zz_when_ArraySlice_l159_295_2 = (_zz_when_ArraySlice_l159_295_3 - _zz_when_ArraySlice_l159_295_4);
  assign _zz_when_ArraySlice_l159_295_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_295_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_295_5);
  assign _zz_when_ArraySlice_l159_295_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_295_5 = {1'd0, _zz_when_ArraySlice_l159_295_6};
  assign _zz__zz_realValue_0_295 = {1'd0, wReg};
  assign _zz__zz_realValue_0_295_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_295_1 = (_zz_realValue_0_295_2 + _zz_realValue_0_295_3);
  assign _zz_realValue_0_295_2 = {1'd0, wReg};
  assign _zz_realValue_0_295_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_295_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_295 = {3'd0, _zz_when_ArraySlice_l166_295_1};
  assign _zz_when_ArraySlice_l166_295_2 = (_zz_when_ArraySlice_l166_295_3 + _zz_when_ArraySlice_l166_295_7);
  assign _zz_when_ArraySlice_l166_295_3 = (realValue_0_295 - _zz_when_ArraySlice_l166_295_4);
  assign _zz_when_ArraySlice_l166_295_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_295_5);
  assign _zz_when_ArraySlice_l166_295_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_295_5 = {1'd0, _zz_when_ArraySlice_l166_295_6};
  assign _zz_when_ArraySlice_l166_295_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_3_2 = (_zz_when_ArraySlice_l285_3_3 + _zz_when_ArraySlice_l285_3_7);
  assign _zz_when_ArraySlice_l285_3_3 = (_zz_when_ArraySlice_l285_3_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_3_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l285_3_5);
  assign _zz_when_ArraySlice_l285_3_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_3_5 = {1'd0, _zz_when_ArraySlice_l285_3_6};
  assign _zz_when_ArraySlice_l285_3_8 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l285_3_7 = {2'd0, _zz_when_ArraySlice_l285_3_8};
  assign _zz_when_ArraySlice_l288_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_3_2 = (_zz_when_ArraySlice_l288_3_3 + 8'h01);
  assign _zz_when_ArraySlice_l288_3_3 = (selectReadFifo_3 + _zz_when_ArraySlice_l288_3_4);
  assign _zz_when_ArraySlice_l288_3_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_3_4 = {1'd0, _zz_when_ArraySlice_l288_3_5};
  assign _zz_selectReadFifo_3_27 = (selectReadFifo_3 + _zz_selectReadFifo_3_28);
  assign _zz_selectReadFifo_3_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_3_28 = {1'd0, _zz_selectReadFifo_3_29};
  assign _zz_when_ArraySlice_l295_3 = (_zz_when_ArraySlice_l295_3_1 % aReg);
  assign _zz_when_ArraySlice_l295_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_3_1 = (_zz_when_ArraySlice_l306_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l306_3 = {5'd0, _zz_when_ArraySlice_l306_3_1};
  assign _zz_when_ArraySlice_l306_3_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_35 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_35_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_35_1 = (_zz_realValue1_0_35_2 + _zz_realValue1_0_35_3);
  assign _zz_realValue1_0_35_2 = {1'd0, hReg};
  assign _zz_realValue1_0_35_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_3_1 = (outSliceNumb_3_value + 7'h01);
  assign _zz_when_ArraySlice_l307_3 = {1'd0, _zz_when_ArraySlice_l307_3_1};
  assign _zz_when_ArraySlice_l307_3_2 = (realValue1_0_35 / aReg);
  assign _zz_selectReadFifo_3_30 = (selectReadFifo_3 - _zz_selectReadFifo_3_31);
  assign _zz_selectReadFifo_3_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_296 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_296_1);
  assign _zz_when_ArraySlice_l158_296_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_296_1 = {4'd0, _zz_when_ArraySlice_l158_296_2};
  assign _zz_when_ArraySlice_l158_296_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_296 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_296_1 = (_zz_when_ArraySlice_l159_296_2 - _zz_when_ArraySlice_l159_296_3);
  assign _zz_when_ArraySlice_l159_296_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_296_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_296_4);
  assign _zz_when_ArraySlice_l159_296_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_296_4 = {4'd0, _zz_when_ArraySlice_l159_296_5};
  assign _zz__zz_realValue_0_296 = {1'd0, wReg};
  assign _zz__zz_realValue_0_296_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_296_1 = (_zz_realValue_0_296_2 + _zz_realValue_0_296_3);
  assign _zz_realValue_0_296_2 = {1'd0, wReg};
  assign _zz_realValue_0_296_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_296 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_296_1 = (_zz_when_ArraySlice_l166_296_2 + _zz_when_ArraySlice_l166_296_6);
  assign _zz_when_ArraySlice_l166_296_2 = (realValue_0_296 - _zz_when_ArraySlice_l166_296_3);
  assign _zz_when_ArraySlice_l166_296_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_296_4);
  assign _zz_when_ArraySlice_l166_296_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_296_4 = {4'd0, _zz_when_ArraySlice_l166_296_5};
  assign _zz_when_ArraySlice_l166_296_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_297 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_297_1);
  assign _zz_when_ArraySlice_l158_297_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_297_1 = {3'd0, _zz_when_ArraySlice_l158_297_2};
  assign _zz_when_ArraySlice_l158_297_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_297_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_297 = {1'd0, _zz_when_ArraySlice_l159_297_1};
  assign _zz_when_ArraySlice_l159_297_2 = (_zz_when_ArraySlice_l159_297_3 - _zz_when_ArraySlice_l159_297_4);
  assign _zz_when_ArraySlice_l159_297_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_297_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_297_5);
  assign _zz_when_ArraySlice_l159_297_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_297_5 = {3'd0, _zz_when_ArraySlice_l159_297_6};
  assign _zz__zz_realValue_0_297 = {1'd0, wReg};
  assign _zz__zz_realValue_0_297_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_297_1 = (_zz_realValue_0_297_2 + _zz_realValue_0_297_3);
  assign _zz_realValue_0_297_2 = {1'd0, wReg};
  assign _zz_realValue_0_297_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_297_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_297 = {1'd0, _zz_when_ArraySlice_l166_297_1};
  assign _zz_when_ArraySlice_l166_297_2 = (_zz_when_ArraySlice_l166_297_3 + _zz_when_ArraySlice_l166_297_7);
  assign _zz_when_ArraySlice_l166_297_3 = (realValue_0_297 - _zz_when_ArraySlice_l166_297_4);
  assign _zz_when_ArraySlice_l166_297_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_297_5);
  assign _zz_when_ArraySlice_l166_297_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_297_5 = {3'd0, _zz_when_ArraySlice_l166_297_6};
  assign _zz_when_ArraySlice_l166_297_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_298 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_298_1);
  assign _zz_when_ArraySlice_l158_298_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_298_1 = {2'd0, _zz_when_ArraySlice_l158_298_2};
  assign _zz_when_ArraySlice_l158_298_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_298_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_298 = {1'd0, _zz_when_ArraySlice_l159_298_1};
  assign _zz_when_ArraySlice_l159_298_2 = (_zz_when_ArraySlice_l159_298_3 - _zz_when_ArraySlice_l159_298_4);
  assign _zz_when_ArraySlice_l159_298_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_298_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_298_5);
  assign _zz_when_ArraySlice_l159_298_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_298_5 = {2'd0, _zz_when_ArraySlice_l159_298_6};
  assign _zz__zz_realValue_0_298 = {1'd0, wReg};
  assign _zz__zz_realValue_0_298_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_298_1 = (_zz_realValue_0_298_2 + _zz_realValue_0_298_3);
  assign _zz_realValue_0_298_2 = {1'd0, wReg};
  assign _zz_realValue_0_298_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_298_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_298 = {1'd0, _zz_when_ArraySlice_l166_298_1};
  assign _zz_when_ArraySlice_l166_298_2 = (_zz_when_ArraySlice_l166_298_3 + _zz_when_ArraySlice_l166_298_7);
  assign _zz_when_ArraySlice_l166_298_3 = (realValue_0_298 - _zz_when_ArraySlice_l166_298_4);
  assign _zz_when_ArraySlice_l166_298_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_298_5);
  assign _zz_when_ArraySlice_l166_298_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_298_5 = {2'd0, _zz_when_ArraySlice_l166_298_6};
  assign _zz_when_ArraySlice_l166_298_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_299 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_299_1);
  assign _zz_when_ArraySlice_l158_299_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_299_1 = {2'd0, _zz_when_ArraySlice_l158_299_2};
  assign _zz_when_ArraySlice_l158_299_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_299_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_299 = {1'd0, _zz_when_ArraySlice_l159_299_1};
  assign _zz_when_ArraySlice_l159_299_2 = (_zz_when_ArraySlice_l159_299_3 - _zz_when_ArraySlice_l159_299_4);
  assign _zz_when_ArraySlice_l159_299_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_299_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_299_5);
  assign _zz_when_ArraySlice_l159_299_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_299_5 = {2'd0, _zz_when_ArraySlice_l159_299_6};
  assign _zz__zz_realValue_0_299 = {1'd0, wReg};
  assign _zz__zz_realValue_0_299_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_299_1 = (_zz_realValue_0_299_2 + _zz_realValue_0_299_3);
  assign _zz_realValue_0_299_2 = {1'd0, wReg};
  assign _zz_realValue_0_299_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_299_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_299 = {1'd0, _zz_when_ArraySlice_l166_299_1};
  assign _zz_when_ArraySlice_l166_299_2 = (_zz_when_ArraySlice_l166_299_3 + _zz_when_ArraySlice_l166_299_7);
  assign _zz_when_ArraySlice_l166_299_3 = (realValue_0_299 - _zz_when_ArraySlice_l166_299_4);
  assign _zz_when_ArraySlice_l166_299_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_299_5);
  assign _zz_when_ArraySlice_l166_299_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_299_5 = {2'd0, _zz_when_ArraySlice_l166_299_6};
  assign _zz_when_ArraySlice_l166_299_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_300 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_300_1);
  assign _zz_when_ArraySlice_l158_300_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_300_1 = {1'd0, _zz_when_ArraySlice_l158_300_2};
  assign _zz_when_ArraySlice_l158_300_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_300_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_300 = {1'd0, _zz_when_ArraySlice_l159_300_1};
  assign _zz_when_ArraySlice_l159_300_2 = (_zz_when_ArraySlice_l159_300_3 - _zz_when_ArraySlice_l159_300_4);
  assign _zz_when_ArraySlice_l159_300_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_300_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_300_5);
  assign _zz_when_ArraySlice_l159_300_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_300_5 = {1'd0, _zz_when_ArraySlice_l159_300_6};
  assign _zz__zz_realValue_0_300 = {1'd0, wReg};
  assign _zz__zz_realValue_0_300_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_300_1 = (_zz_realValue_0_300_2 + _zz_realValue_0_300_3);
  assign _zz_realValue_0_300_2 = {1'd0, wReg};
  assign _zz_realValue_0_300_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_300_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_300 = {1'd0, _zz_when_ArraySlice_l166_300_1};
  assign _zz_when_ArraySlice_l166_300_2 = (_zz_when_ArraySlice_l166_300_3 + _zz_when_ArraySlice_l166_300_7);
  assign _zz_when_ArraySlice_l166_300_3 = (realValue_0_300 - _zz_when_ArraySlice_l166_300_4);
  assign _zz_when_ArraySlice_l166_300_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_300_5);
  assign _zz_when_ArraySlice_l166_300_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_300_5 = {1'd0, _zz_when_ArraySlice_l166_300_6};
  assign _zz_when_ArraySlice_l166_300_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_301 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_301_1);
  assign _zz_when_ArraySlice_l158_301_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_301_1 = {1'd0, _zz_when_ArraySlice_l158_301_2};
  assign _zz_when_ArraySlice_l158_301_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_301_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_301 = {2'd0, _zz_when_ArraySlice_l159_301_1};
  assign _zz_when_ArraySlice_l159_301_2 = (_zz_when_ArraySlice_l159_301_3 - _zz_when_ArraySlice_l159_301_4);
  assign _zz_when_ArraySlice_l159_301_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_301_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_301_5);
  assign _zz_when_ArraySlice_l159_301_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_301_5 = {1'd0, _zz_when_ArraySlice_l159_301_6};
  assign _zz__zz_realValue_0_301 = {1'd0, wReg};
  assign _zz__zz_realValue_0_301_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_301_1 = (_zz_realValue_0_301_2 + _zz_realValue_0_301_3);
  assign _zz_realValue_0_301_2 = {1'd0, wReg};
  assign _zz_realValue_0_301_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_301_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_301 = {2'd0, _zz_when_ArraySlice_l166_301_1};
  assign _zz_when_ArraySlice_l166_301_2 = (_zz_when_ArraySlice_l166_301_3 + _zz_when_ArraySlice_l166_301_7);
  assign _zz_when_ArraySlice_l166_301_3 = (realValue_0_301 - _zz_when_ArraySlice_l166_301_4);
  assign _zz_when_ArraySlice_l166_301_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_301_5);
  assign _zz_when_ArraySlice_l166_301_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_301_5 = {1'd0, _zz_when_ArraySlice_l166_301_6};
  assign _zz_when_ArraySlice_l166_301_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_302 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_302_1);
  assign _zz_when_ArraySlice_l158_302_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_302_1 = {1'd0, _zz_when_ArraySlice_l158_302_2};
  assign _zz_when_ArraySlice_l158_302_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_302_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_302 = {2'd0, _zz_when_ArraySlice_l159_302_1};
  assign _zz_when_ArraySlice_l159_302_2 = (_zz_when_ArraySlice_l159_302_3 - _zz_when_ArraySlice_l159_302_4);
  assign _zz_when_ArraySlice_l159_302_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_302_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_302_5);
  assign _zz_when_ArraySlice_l159_302_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_302_5 = {1'd0, _zz_when_ArraySlice_l159_302_6};
  assign _zz__zz_realValue_0_302 = {1'd0, wReg};
  assign _zz__zz_realValue_0_302_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_302_1 = (_zz_realValue_0_302_2 + _zz_realValue_0_302_3);
  assign _zz_realValue_0_302_2 = {1'd0, wReg};
  assign _zz_realValue_0_302_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_302_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_302 = {2'd0, _zz_when_ArraySlice_l166_302_1};
  assign _zz_when_ArraySlice_l166_302_2 = (_zz_when_ArraySlice_l166_302_3 + _zz_when_ArraySlice_l166_302_7);
  assign _zz_when_ArraySlice_l166_302_3 = (realValue_0_302 - _zz_when_ArraySlice_l166_302_4);
  assign _zz_when_ArraySlice_l166_302_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_302_5);
  assign _zz_when_ArraySlice_l166_302_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_302_5 = {1'd0, _zz_when_ArraySlice_l166_302_6};
  assign _zz_when_ArraySlice_l166_302_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_303 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_303_1);
  assign _zz_when_ArraySlice_l158_303_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_303_1 = {1'd0, _zz_when_ArraySlice_l158_303_2};
  assign _zz_when_ArraySlice_l158_303_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_303_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_303 = {3'd0, _zz_when_ArraySlice_l159_303_1};
  assign _zz_when_ArraySlice_l159_303_2 = (_zz_when_ArraySlice_l159_303_3 - _zz_when_ArraySlice_l159_303_4);
  assign _zz_when_ArraySlice_l159_303_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_303_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_303_5);
  assign _zz_when_ArraySlice_l159_303_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_303_5 = {1'd0, _zz_when_ArraySlice_l159_303_6};
  assign _zz__zz_realValue_0_303 = {1'd0, wReg};
  assign _zz__zz_realValue_0_303_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_303_1 = (_zz_realValue_0_303_2 + _zz_realValue_0_303_3);
  assign _zz_realValue_0_303_2 = {1'd0, wReg};
  assign _zz_realValue_0_303_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_303_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_303 = {3'd0, _zz_when_ArraySlice_l166_303_1};
  assign _zz_when_ArraySlice_l166_303_2 = (_zz_when_ArraySlice_l166_303_3 + _zz_when_ArraySlice_l166_303_7);
  assign _zz_when_ArraySlice_l166_303_3 = (realValue_0_303 - _zz_when_ArraySlice_l166_303_4);
  assign _zz_when_ArraySlice_l166_303_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_303_5);
  assign _zz_when_ArraySlice_l166_303_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_303_5 = {1'd0, _zz_when_ArraySlice_l166_303_6};
  assign _zz_when_ArraySlice_l166_303_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_3 = (_zz_when_ArraySlice_l318_3_1 % aReg);
  assign _zz_when_ArraySlice_l318_3_1 = (handshakeTimes_3_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_3_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_3_2 = (selectReadFifo_3 + _zz_when_ArraySlice_l304_3_3);
  assign _zz_when_ArraySlice_l304_3_4 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l304_3_3 = {2'd0, _zz_when_ArraySlice_l304_3_4};
  assign _zz_when_ArraySlice_l325_3_1 = (_zz_when_ArraySlice_l325_3_2 - 8'h01);
  assign _zz_when_ArraySlice_l325_3 = {5'd0, _zz_when_ArraySlice_l325_3_1};
  assign _zz_when_ArraySlice_l325_3_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l233_4_1);
  assign _zz_when_ArraySlice_l233_4_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l233_4_1 = {1'd0, _zz_when_ArraySlice_l233_4_2};
  assign _zz_when_ArraySlice_l233_4_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l234_4_4);
  assign _zz_when_ArraySlice_l234_4_2 = _zz_when_ArraySlice_l234_4_3[6:0];
  assign _zz_when_ArraySlice_l234_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l234_4_4 = {1'd0, _zz_when_ArraySlice_l234_4_5};
  assign _zz__zz_outputStreamArrayData_4_valid_1_2 = (bReg * 3'b100);
  assign _zz__zz_outputStreamArrayData_4_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_4_valid_1_2};
  assign _zz__zz_15 = _zz_outputStreamArrayData_4_valid_1[6:0];
  assign _zz_outputStreamArrayData_4_valid_5 = _zz_outputStreamArrayData_4_valid_1[6:0];
  assign _zz_outputStreamArrayData_4_payload_3 = _zz_outputStreamArrayData_4_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l240_4_4);
  assign _zz_when_ArraySlice_l240_4_2 = _zz_when_ArraySlice_l240_4_3[6:0];
  assign _zz_when_ArraySlice_l240_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l240_4_4 = {1'd0, _zz_when_ArraySlice_l240_4_5};
  assign _zz_when_ArraySlice_l241_4_1 = (_zz_when_ArraySlice_l241_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l241_4 = {5'd0, _zz_when_ArraySlice_l241_4_1};
  assign _zz_when_ArraySlice_l241_4_2 = (bReg * aReg);
  assign _zz_selectReadFifo_4_16 = (selectReadFifo_4 - _zz_selectReadFifo_4_17);
  assign _zz_selectReadFifo_4_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_4 = (_zz_when_ArraySlice_l244_4_1 % aReg);
  assign _zz_when_ArraySlice_l244_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l249_4_4);
  assign _zz_when_ArraySlice_l249_4_2 = _zz_when_ArraySlice_l249_4_3[6:0];
  assign _zz_when_ArraySlice_l249_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l249_4_4 = {1'd0, _zz_when_ArraySlice_l249_4_5};
  assign _zz_when_ArraySlice_l250_4_1 = (_zz_when_ArraySlice_l250_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l250_4 = {5'd0, _zz_when_ArraySlice_l250_4_1};
  assign _zz_when_ArraySlice_l250_4_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_36 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_36_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_36_1 = (_zz_realValue1_0_36_2 + _zz_realValue1_0_36_3);
  assign _zz_realValue1_0_36_2 = {1'd0, hReg};
  assign _zz_realValue1_0_36_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l252_4 = {1'd0, _zz_when_ArraySlice_l252_4_1};
  assign _zz_when_ArraySlice_l252_4_2 = (realValue1_0_36 / aReg);
  assign _zz_selectReadFifo_4_18 = (selectReadFifo_4 - _zz_selectReadFifo_4_19);
  assign _zz_selectReadFifo_4_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_4_21 = 1'b1;
  assign _zz_selectReadFifo_4_20 = {7'd0, _zz_selectReadFifo_4_21};
  assign _zz_when_ArraySlice_l158_304 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_304_1);
  assign _zz_when_ArraySlice_l158_304_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_304_1 = {4'd0, _zz_when_ArraySlice_l158_304_2};
  assign _zz_when_ArraySlice_l158_304_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_304 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_304_1 = (_zz_when_ArraySlice_l159_304_2 - _zz_when_ArraySlice_l159_304_3);
  assign _zz_when_ArraySlice_l159_304_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_304_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_304_4);
  assign _zz_when_ArraySlice_l159_304_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_304_4 = {4'd0, _zz_when_ArraySlice_l159_304_5};
  assign _zz__zz_realValue_0_304 = {1'd0, wReg};
  assign _zz__zz_realValue_0_304_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_304_1 = (_zz_realValue_0_304_2 + _zz_realValue_0_304_3);
  assign _zz_realValue_0_304_2 = {1'd0, wReg};
  assign _zz_realValue_0_304_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_304 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_304_1 = (_zz_when_ArraySlice_l166_304_2 + _zz_when_ArraySlice_l166_304_6);
  assign _zz_when_ArraySlice_l166_304_2 = (realValue_0_304 - _zz_when_ArraySlice_l166_304_3);
  assign _zz_when_ArraySlice_l166_304_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_304_4);
  assign _zz_when_ArraySlice_l166_304_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_304_4 = {4'd0, _zz_when_ArraySlice_l166_304_5};
  assign _zz_when_ArraySlice_l166_304_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_305 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_305_1);
  assign _zz_when_ArraySlice_l158_305_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_305_1 = {3'd0, _zz_when_ArraySlice_l158_305_2};
  assign _zz_when_ArraySlice_l158_305_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_305_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_305 = {1'd0, _zz_when_ArraySlice_l159_305_1};
  assign _zz_when_ArraySlice_l159_305_2 = (_zz_when_ArraySlice_l159_305_3 - _zz_when_ArraySlice_l159_305_4);
  assign _zz_when_ArraySlice_l159_305_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_305_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_305_5);
  assign _zz_when_ArraySlice_l159_305_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_305_5 = {3'd0, _zz_when_ArraySlice_l159_305_6};
  assign _zz__zz_realValue_0_305 = {1'd0, wReg};
  assign _zz__zz_realValue_0_305_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_305_1 = (_zz_realValue_0_305_2 + _zz_realValue_0_305_3);
  assign _zz_realValue_0_305_2 = {1'd0, wReg};
  assign _zz_realValue_0_305_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_305_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_305 = {1'd0, _zz_when_ArraySlice_l166_305_1};
  assign _zz_when_ArraySlice_l166_305_2 = (_zz_when_ArraySlice_l166_305_3 + _zz_when_ArraySlice_l166_305_7);
  assign _zz_when_ArraySlice_l166_305_3 = (realValue_0_305 - _zz_when_ArraySlice_l166_305_4);
  assign _zz_when_ArraySlice_l166_305_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_305_5);
  assign _zz_when_ArraySlice_l166_305_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_305_5 = {3'd0, _zz_when_ArraySlice_l166_305_6};
  assign _zz_when_ArraySlice_l166_305_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_306 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_306_1);
  assign _zz_when_ArraySlice_l158_306_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_306_1 = {2'd0, _zz_when_ArraySlice_l158_306_2};
  assign _zz_when_ArraySlice_l158_306_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_306_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_306 = {1'd0, _zz_when_ArraySlice_l159_306_1};
  assign _zz_when_ArraySlice_l159_306_2 = (_zz_when_ArraySlice_l159_306_3 - _zz_when_ArraySlice_l159_306_4);
  assign _zz_when_ArraySlice_l159_306_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_306_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_306_5);
  assign _zz_when_ArraySlice_l159_306_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_306_5 = {2'd0, _zz_when_ArraySlice_l159_306_6};
  assign _zz__zz_realValue_0_306 = {1'd0, wReg};
  assign _zz__zz_realValue_0_306_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_306_1 = (_zz_realValue_0_306_2 + _zz_realValue_0_306_3);
  assign _zz_realValue_0_306_2 = {1'd0, wReg};
  assign _zz_realValue_0_306_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_306_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_306 = {1'd0, _zz_when_ArraySlice_l166_306_1};
  assign _zz_when_ArraySlice_l166_306_2 = (_zz_when_ArraySlice_l166_306_3 + _zz_when_ArraySlice_l166_306_7);
  assign _zz_when_ArraySlice_l166_306_3 = (realValue_0_306 - _zz_when_ArraySlice_l166_306_4);
  assign _zz_when_ArraySlice_l166_306_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_306_5);
  assign _zz_when_ArraySlice_l166_306_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_306_5 = {2'd0, _zz_when_ArraySlice_l166_306_6};
  assign _zz_when_ArraySlice_l166_306_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_307 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_307_1);
  assign _zz_when_ArraySlice_l158_307_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_307_1 = {2'd0, _zz_when_ArraySlice_l158_307_2};
  assign _zz_when_ArraySlice_l158_307_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_307_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_307 = {1'd0, _zz_when_ArraySlice_l159_307_1};
  assign _zz_when_ArraySlice_l159_307_2 = (_zz_when_ArraySlice_l159_307_3 - _zz_when_ArraySlice_l159_307_4);
  assign _zz_when_ArraySlice_l159_307_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_307_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_307_5);
  assign _zz_when_ArraySlice_l159_307_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_307_5 = {2'd0, _zz_when_ArraySlice_l159_307_6};
  assign _zz__zz_realValue_0_307 = {1'd0, wReg};
  assign _zz__zz_realValue_0_307_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_307_1 = (_zz_realValue_0_307_2 + _zz_realValue_0_307_3);
  assign _zz_realValue_0_307_2 = {1'd0, wReg};
  assign _zz_realValue_0_307_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_307_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_307 = {1'd0, _zz_when_ArraySlice_l166_307_1};
  assign _zz_when_ArraySlice_l166_307_2 = (_zz_when_ArraySlice_l166_307_3 + _zz_when_ArraySlice_l166_307_7);
  assign _zz_when_ArraySlice_l166_307_3 = (realValue_0_307 - _zz_when_ArraySlice_l166_307_4);
  assign _zz_when_ArraySlice_l166_307_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_307_5);
  assign _zz_when_ArraySlice_l166_307_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_307_5 = {2'd0, _zz_when_ArraySlice_l166_307_6};
  assign _zz_when_ArraySlice_l166_307_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_308 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_308_1);
  assign _zz_when_ArraySlice_l158_308_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_308_1 = {1'd0, _zz_when_ArraySlice_l158_308_2};
  assign _zz_when_ArraySlice_l158_308_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_308_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_308 = {1'd0, _zz_when_ArraySlice_l159_308_1};
  assign _zz_when_ArraySlice_l159_308_2 = (_zz_when_ArraySlice_l159_308_3 - _zz_when_ArraySlice_l159_308_4);
  assign _zz_when_ArraySlice_l159_308_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_308_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_308_5);
  assign _zz_when_ArraySlice_l159_308_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_308_5 = {1'd0, _zz_when_ArraySlice_l159_308_6};
  assign _zz__zz_realValue_0_308 = {1'd0, wReg};
  assign _zz__zz_realValue_0_308_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_308_1 = (_zz_realValue_0_308_2 + _zz_realValue_0_308_3);
  assign _zz_realValue_0_308_2 = {1'd0, wReg};
  assign _zz_realValue_0_308_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_308_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_308 = {1'd0, _zz_when_ArraySlice_l166_308_1};
  assign _zz_when_ArraySlice_l166_308_2 = (_zz_when_ArraySlice_l166_308_3 + _zz_when_ArraySlice_l166_308_7);
  assign _zz_when_ArraySlice_l166_308_3 = (realValue_0_308 - _zz_when_ArraySlice_l166_308_4);
  assign _zz_when_ArraySlice_l166_308_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_308_5);
  assign _zz_when_ArraySlice_l166_308_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_308_5 = {1'd0, _zz_when_ArraySlice_l166_308_6};
  assign _zz_when_ArraySlice_l166_308_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_309 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_309_1);
  assign _zz_when_ArraySlice_l158_309_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_309_1 = {1'd0, _zz_when_ArraySlice_l158_309_2};
  assign _zz_when_ArraySlice_l158_309_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_309_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_309 = {2'd0, _zz_when_ArraySlice_l159_309_1};
  assign _zz_when_ArraySlice_l159_309_2 = (_zz_when_ArraySlice_l159_309_3 - _zz_when_ArraySlice_l159_309_4);
  assign _zz_when_ArraySlice_l159_309_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_309_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_309_5);
  assign _zz_when_ArraySlice_l159_309_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_309_5 = {1'd0, _zz_when_ArraySlice_l159_309_6};
  assign _zz__zz_realValue_0_309 = {1'd0, wReg};
  assign _zz__zz_realValue_0_309_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_309_1 = (_zz_realValue_0_309_2 + _zz_realValue_0_309_3);
  assign _zz_realValue_0_309_2 = {1'd0, wReg};
  assign _zz_realValue_0_309_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_309_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_309 = {2'd0, _zz_when_ArraySlice_l166_309_1};
  assign _zz_when_ArraySlice_l166_309_2 = (_zz_when_ArraySlice_l166_309_3 + _zz_when_ArraySlice_l166_309_7);
  assign _zz_when_ArraySlice_l166_309_3 = (realValue_0_309 - _zz_when_ArraySlice_l166_309_4);
  assign _zz_when_ArraySlice_l166_309_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_309_5);
  assign _zz_when_ArraySlice_l166_309_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_309_5 = {1'd0, _zz_when_ArraySlice_l166_309_6};
  assign _zz_when_ArraySlice_l166_309_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_310 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_310_1);
  assign _zz_when_ArraySlice_l158_310_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_310_1 = {1'd0, _zz_when_ArraySlice_l158_310_2};
  assign _zz_when_ArraySlice_l158_310_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_310_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_310 = {2'd0, _zz_when_ArraySlice_l159_310_1};
  assign _zz_when_ArraySlice_l159_310_2 = (_zz_when_ArraySlice_l159_310_3 - _zz_when_ArraySlice_l159_310_4);
  assign _zz_when_ArraySlice_l159_310_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_310_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_310_5);
  assign _zz_when_ArraySlice_l159_310_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_310_5 = {1'd0, _zz_when_ArraySlice_l159_310_6};
  assign _zz__zz_realValue_0_310 = {1'd0, wReg};
  assign _zz__zz_realValue_0_310_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_310_1 = (_zz_realValue_0_310_2 + _zz_realValue_0_310_3);
  assign _zz_realValue_0_310_2 = {1'd0, wReg};
  assign _zz_realValue_0_310_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_310_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_310 = {2'd0, _zz_when_ArraySlice_l166_310_1};
  assign _zz_when_ArraySlice_l166_310_2 = (_zz_when_ArraySlice_l166_310_3 + _zz_when_ArraySlice_l166_310_7);
  assign _zz_when_ArraySlice_l166_310_3 = (realValue_0_310 - _zz_when_ArraySlice_l166_310_4);
  assign _zz_when_ArraySlice_l166_310_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_310_5);
  assign _zz_when_ArraySlice_l166_310_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_310_5 = {1'd0, _zz_when_ArraySlice_l166_310_6};
  assign _zz_when_ArraySlice_l166_310_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_311 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_311_1);
  assign _zz_when_ArraySlice_l158_311_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_311_1 = {1'd0, _zz_when_ArraySlice_l158_311_2};
  assign _zz_when_ArraySlice_l158_311_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_311_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_311 = {3'd0, _zz_when_ArraySlice_l159_311_1};
  assign _zz_when_ArraySlice_l159_311_2 = (_zz_when_ArraySlice_l159_311_3 - _zz_when_ArraySlice_l159_311_4);
  assign _zz_when_ArraySlice_l159_311_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_311_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_311_5);
  assign _zz_when_ArraySlice_l159_311_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_311_5 = {1'd0, _zz_when_ArraySlice_l159_311_6};
  assign _zz__zz_realValue_0_311 = {1'd0, wReg};
  assign _zz__zz_realValue_0_311_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_311_1 = (_zz_realValue_0_311_2 + _zz_realValue_0_311_3);
  assign _zz_realValue_0_311_2 = {1'd0, wReg};
  assign _zz_realValue_0_311_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_311_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_311 = {3'd0, _zz_when_ArraySlice_l166_311_1};
  assign _zz_when_ArraySlice_l166_311_2 = (_zz_when_ArraySlice_l166_311_3 + _zz_when_ArraySlice_l166_311_7);
  assign _zz_when_ArraySlice_l166_311_3 = (realValue_0_311 - _zz_when_ArraySlice_l166_311_4);
  assign _zz_when_ArraySlice_l166_311_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_311_5);
  assign _zz_when_ArraySlice_l166_311_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_311_5 = {1'd0, _zz_when_ArraySlice_l166_311_6};
  assign _zz_when_ArraySlice_l166_311_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_4_2 = (_zz_when_ArraySlice_l260_4_3 + _zz_when_ArraySlice_l260_4_7);
  assign _zz_when_ArraySlice_l260_4_3 = (_zz_when_ArraySlice_l260_4_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l260_4_5);
  assign _zz_when_ArraySlice_l260_4_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_4_5 = {1'd0, _zz_when_ArraySlice_l260_4_6};
  assign _zz_when_ArraySlice_l260_4_8 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l260_4_7 = {1'd0, _zz_when_ArraySlice_l260_4_8};
  assign _zz_when_ArraySlice_l263_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_4_2 = (_zz_when_ArraySlice_l263_4_3 + 8'h01);
  assign _zz_when_ArraySlice_l263_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l263_4_4);
  assign _zz_when_ArraySlice_l263_4_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_4_4 = {1'd0, _zz_when_ArraySlice_l263_4_5};
  assign _zz_selectReadFifo_4_22 = (selectReadFifo_4 + _zz_selectReadFifo_4_23);
  assign _zz_selectReadFifo_4_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_23 = {1'd0, _zz_selectReadFifo_4_24};
  assign _zz_when_ArraySlice_l270_4 = (_zz_when_ArraySlice_l270_4_1 % aReg);
  assign _zz_when_ArraySlice_l270_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l274_4_4);
  assign _zz_when_ArraySlice_l274_4_2 = _zz_when_ArraySlice_l274_4_3[6:0];
  assign _zz_when_ArraySlice_l274_4_5 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l274_4_4 = {1'd0, _zz_when_ArraySlice_l274_4_5};
  assign _zz_when_ArraySlice_l275_4_2 = (_zz_when_ArraySlice_l275_4_3 - _zz_when_ArraySlice_l275_4_4);
  assign _zz_when_ArraySlice_l275_4_1 = {5'd0, _zz_when_ArraySlice_l275_4_2};
  assign _zz_when_ArraySlice_l275_4_3 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_4_5 = 1'b1;
  assign _zz_when_ArraySlice_l275_4_4 = {7'd0, _zz_when_ArraySlice_l275_4_5};
  assign _zz__zz_realValue1_0_37 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_37_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_37_1 = (_zz_realValue1_0_37_2 + _zz_realValue1_0_37_3);
  assign _zz_realValue1_0_37_2 = {1'd0, hReg};
  assign _zz_realValue1_0_37_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l277_4 = {1'd0, _zz_when_ArraySlice_l277_4_1};
  assign _zz_when_ArraySlice_l277_4_2 = (realValue1_0_37 / aReg);
  assign _zz_selectReadFifo_4_25 = (selectReadFifo_4 - _zz_selectReadFifo_4_26);
  assign _zz_selectReadFifo_4_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_312 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_312_1);
  assign _zz_when_ArraySlice_l158_312_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_312_1 = {4'd0, _zz_when_ArraySlice_l158_312_2};
  assign _zz_when_ArraySlice_l158_312_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_312 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_312_1 = (_zz_when_ArraySlice_l159_312_2 - _zz_when_ArraySlice_l159_312_3);
  assign _zz_when_ArraySlice_l159_312_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_312_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_312_4);
  assign _zz_when_ArraySlice_l159_312_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_312_4 = {4'd0, _zz_when_ArraySlice_l159_312_5};
  assign _zz__zz_realValue_0_312 = {1'd0, wReg};
  assign _zz__zz_realValue_0_312_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_312_1 = (_zz_realValue_0_312_2 + _zz_realValue_0_312_3);
  assign _zz_realValue_0_312_2 = {1'd0, wReg};
  assign _zz_realValue_0_312_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_312 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_312_1 = (_zz_when_ArraySlice_l166_312_2 + _zz_when_ArraySlice_l166_312_6);
  assign _zz_when_ArraySlice_l166_312_2 = (realValue_0_312 - _zz_when_ArraySlice_l166_312_3);
  assign _zz_when_ArraySlice_l166_312_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_312_4);
  assign _zz_when_ArraySlice_l166_312_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_312_4 = {4'd0, _zz_when_ArraySlice_l166_312_5};
  assign _zz_when_ArraySlice_l166_312_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_313 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_313_1);
  assign _zz_when_ArraySlice_l158_313_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_313_1 = {3'd0, _zz_when_ArraySlice_l158_313_2};
  assign _zz_when_ArraySlice_l158_313_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_313_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_313 = {1'd0, _zz_when_ArraySlice_l159_313_1};
  assign _zz_when_ArraySlice_l159_313_2 = (_zz_when_ArraySlice_l159_313_3 - _zz_when_ArraySlice_l159_313_4);
  assign _zz_when_ArraySlice_l159_313_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_313_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_313_5);
  assign _zz_when_ArraySlice_l159_313_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_313_5 = {3'd0, _zz_when_ArraySlice_l159_313_6};
  assign _zz__zz_realValue_0_313 = {1'd0, wReg};
  assign _zz__zz_realValue_0_313_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_313_1 = (_zz_realValue_0_313_2 + _zz_realValue_0_313_3);
  assign _zz_realValue_0_313_2 = {1'd0, wReg};
  assign _zz_realValue_0_313_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_313_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_313 = {1'd0, _zz_when_ArraySlice_l166_313_1};
  assign _zz_when_ArraySlice_l166_313_2 = (_zz_when_ArraySlice_l166_313_3 + _zz_when_ArraySlice_l166_313_7);
  assign _zz_when_ArraySlice_l166_313_3 = (realValue_0_313 - _zz_when_ArraySlice_l166_313_4);
  assign _zz_when_ArraySlice_l166_313_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_313_5);
  assign _zz_when_ArraySlice_l166_313_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_313_5 = {3'd0, _zz_when_ArraySlice_l166_313_6};
  assign _zz_when_ArraySlice_l166_313_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_314 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_314_1);
  assign _zz_when_ArraySlice_l158_314_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_314_1 = {2'd0, _zz_when_ArraySlice_l158_314_2};
  assign _zz_when_ArraySlice_l158_314_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_314_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_314 = {1'd0, _zz_when_ArraySlice_l159_314_1};
  assign _zz_when_ArraySlice_l159_314_2 = (_zz_when_ArraySlice_l159_314_3 - _zz_when_ArraySlice_l159_314_4);
  assign _zz_when_ArraySlice_l159_314_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_314_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_314_5);
  assign _zz_when_ArraySlice_l159_314_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_314_5 = {2'd0, _zz_when_ArraySlice_l159_314_6};
  assign _zz__zz_realValue_0_314 = {1'd0, wReg};
  assign _zz__zz_realValue_0_314_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_314_1 = (_zz_realValue_0_314_2 + _zz_realValue_0_314_3);
  assign _zz_realValue_0_314_2 = {1'd0, wReg};
  assign _zz_realValue_0_314_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_314_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_314 = {1'd0, _zz_when_ArraySlice_l166_314_1};
  assign _zz_when_ArraySlice_l166_314_2 = (_zz_when_ArraySlice_l166_314_3 + _zz_when_ArraySlice_l166_314_7);
  assign _zz_when_ArraySlice_l166_314_3 = (realValue_0_314 - _zz_when_ArraySlice_l166_314_4);
  assign _zz_when_ArraySlice_l166_314_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_314_5);
  assign _zz_when_ArraySlice_l166_314_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_314_5 = {2'd0, _zz_when_ArraySlice_l166_314_6};
  assign _zz_when_ArraySlice_l166_314_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_315 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_315_1);
  assign _zz_when_ArraySlice_l158_315_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_315_1 = {2'd0, _zz_when_ArraySlice_l158_315_2};
  assign _zz_when_ArraySlice_l158_315_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_315_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_315 = {1'd0, _zz_when_ArraySlice_l159_315_1};
  assign _zz_when_ArraySlice_l159_315_2 = (_zz_when_ArraySlice_l159_315_3 - _zz_when_ArraySlice_l159_315_4);
  assign _zz_when_ArraySlice_l159_315_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_315_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_315_5);
  assign _zz_when_ArraySlice_l159_315_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_315_5 = {2'd0, _zz_when_ArraySlice_l159_315_6};
  assign _zz__zz_realValue_0_315 = {1'd0, wReg};
  assign _zz__zz_realValue_0_315_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_315_1 = (_zz_realValue_0_315_2 + _zz_realValue_0_315_3);
  assign _zz_realValue_0_315_2 = {1'd0, wReg};
  assign _zz_realValue_0_315_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_315_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_315 = {1'd0, _zz_when_ArraySlice_l166_315_1};
  assign _zz_when_ArraySlice_l166_315_2 = (_zz_when_ArraySlice_l166_315_3 + _zz_when_ArraySlice_l166_315_7);
  assign _zz_when_ArraySlice_l166_315_3 = (realValue_0_315 - _zz_when_ArraySlice_l166_315_4);
  assign _zz_when_ArraySlice_l166_315_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_315_5);
  assign _zz_when_ArraySlice_l166_315_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_315_5 = {2'd0, _zz_when_ArraySlice_l166_315_6};
  assign _zz_when_ArraySlice_l166_315_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_316 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_316_1);
  assign _zz_when_ArraySlice_l158_316_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_316_1 = {1'd0, _zz_when_ArraySlice_l158_316_2};
  assign _zz_when_ArraySlice_l158_316_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_316_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_316 = {1'd0, _zz_when_ArraySlice_l159_316_1};
  assign _zz_when_ArraySlice_l159_316_2 = (_zz_when_ArraySlice_l159_316_3 - _zz_when_ArraySlice_l159_316_4);
  assign _zz_when_ArraySlice_l159_316_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_316_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_316_5);
  assign _zz_when_ArraySlice_l159_316_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_316_5 = {1'd0, _zz_when_ArraySlice_l159_316_6};
  assign _zz__zz_realValue_0_316 = {1'd0, wReg};
  assign _zz__zz_realValue_0_316_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_316_1 = (_zz_realValue_0_316_2 + _zz_realValue_0_316_3);
  assign _zz_realValue_0_316_2 = {1'd0, wReg};
  assign _zz_realValue_0_316_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_316_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_316 = {1'd0, _zz_when_ArraySlice_l166_316_1};
  assign _zz_when_ArraySlice_l166_316_2 = (_zz_when_ArraySlice_l166_316_3 + _zz_when_ArraySlice_l166_316_7);
  assign _zz_when_ArraySlice_l166_316_3 = (realValue_0_316 - _zz_when_ArraySlice_l166_316_4);
  assign _zz_when_ArraySlice_l166_316_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_316_5);
  assign _zz_when_ArraySlice_l166_316_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_316_5 = {1'd0, _zz_when_ArraySlice_l166_316_6};
  assign _zz_when_ArraySlice_l166_316_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_317 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_317_1);
  assign _zz_when_ArraySlice_l158_317_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_317_1 = {1'd0, _zz_when_ArraySlice_l158_317_2};
  assign _zz_when_ArraySlice_l158_317_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_317_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_317 = {2'd0, _zz_when_ArraySlice_l159_317_1};
  assign _zz_when_ArraySlice_l159_317_2 = (_zz_when_ArraySlice_l159_317_3 - _zz_when_ArraySlice_l159_317_4);
  assign _zz_when_ArraySlice_l159_317_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_317_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_317_5);
  assign _zz_when_ArraySlice_l159_317_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_317_5 = {1'd0, _zz_when_ArraySlice_l159_317_6};
  assign _zz__zz_realValue_0_317 = {1'd0, wReg};
  assign _zz__zz_realValue_0_317_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_317_1 = (_zz_realValue_0_317_2 + _zz_realValue_0_317_3);
  assign _zz_realValue_0_317_2 = {1'd0, wReg};
  assign _zz_realValue_0_317_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_317_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_317 = {2'd0, _zz_when_ArraySlice_l166_317_1};
  assign _zz_when_ArraySlice_l166_317_2 = (_zz_when_ArraySlice_l166_317_3 + _zz_when_ArraySlice_l166_317_7);
  assign _zz_when_ArraySlice_l166_317_3 = (realValue_0_317 - _zz_when_ArraySlice_l166_317_4);
  assign _zz_when_ArraySlice_l166_317_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_317_5);
  assign _zz_when_ArraySlice_l166_317_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_317_5 = {1'd0, _zz_when_ArraySlice_l166_317_6};
  assign _zz_when_ArraySlice_l166_317_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_318 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_318_1);
  assign _zz_when_ArraySlice_l158_318_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_318_1 = {1'd0, _zz_when_ArraySlice_l158_318_2};
  assign _zz_when_ArraySlice_l158_318_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_318_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_318 = {2'd0, _zz_when_ArraySlice_l159_318_1};
  assign _zz_when_ArraySlice_l159_318_2 = (_zz_when_ArraySlice_l159_318_3 - _zz_when_ArraySlice_l159_318_4);
  assign _zz_when_ArraySlice_l159_318_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_318_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_318_5);
  assign _zz_when_ArraySlice_l159_318_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_318_5 = {1'd0, _zz_when_ArraySlice_l159_318_6};
  assign _zz__zz_realValue_0_318 = {1'd0, wReg};
  assign _zz__zz_realValue_0_318_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_318_1 = (_zz_realValue_0_318_2 + _zz_realValue_0_318_3);
  assign _zz_realValue_0_318_2 = {1'd0, wReg};
  assign _zz_realValue_0_318_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_318_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_318 = {2'd0, _zz_when_ArraySlice_l166_318_1};
  assign _zz_when_ArraySlice_l166_318_2 = (_zz_when_ArraySlice_l166_318_3 + _zz_when_ArraySlice_l166_318_7);
  assign _zz_when_ArraySlice_l166_318_3 = (realValue_0_318 - _zz_when_ArraySlice_l166_318_4);
  assign _zz_when_ArraySlice_l166_318_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_318_5);
  assign _zz_when_ArraySlice_l166_318_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_318_5 = {1'd0, _zz_when_ArraySlice_l166_318_6};
  assign _zz_when_ArraySlice_l166_318_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_319 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_319_1);
  assign _zz_when_ArraySlice_l158_319_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_319_1 = {1'd0, _zz_when_ArraySlice_l158_319_2};
  assign _zz_when_ArraySlice_l158_319_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_319_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_319 = {3'd0, _zz_when_ArraySlice_l159_319_1};
  assign _zz_when_ArraySlice_l159_319_2 = (_zz_when_ArraySlice_l159_319_3 - _zz_when_ArraySlice_l159_319_4);
  assign _zz_when_ArraySlice_l159_319_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_319_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_319_5);
  assign _zz_when_ArraySlice_l159_319_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_319_5 = {1'd0, _zz_when_ArraySlice_l159_319_6};
  assign _zz__zz_realValue_0_319 = {1'd0, wReg};
  assign _zz__zz_realValue_0_319_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_319_1 = (_zz_realValue_0_319_2 + _zz_realValue_0_319_3);
  assign _zz_realValue_0_319_2 = {1'd0, wReg};
  assign _zz_realValue_0_319_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_319_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_319 = {3'd0, _zz_when_ArraySlice_l166_319_1};
  assign _zz_when_ArraySlice_l166_319_2 = (_zz_when_ArraySlice_l166_319_3 + _zz_when_ArraySlice_l166_319_7);
  assign _zz_when_ArraySlice_l166_319_3 = (realValue_0_319 - _zz_when_ArraySlice_l166_319_4);
  assign _zz_when_ArraySlice_l166_319_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_319_5);
  assign _zz_when_ArraySlice_l166_319_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_319_5 = {1'd0, _zz_when_ArraySlice_l166_319_6};
  assign _zz_when_ArraySlice_l166_319_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_4_2 = (_zz_when_ArraySlice_l285_4_3 + _zz_when_ArraySlice_l285_4_7);
  assign _zz_when_ArraySlice_l285_4_3 = (_zz_when_ArraySlice_l285_4_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_4_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l285_4_5);
  assign _zz_when_ArraySlice_l285_4_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_4_5 = {1'd0, _zz_when_ArraySlice_l285_4_6};
  assign _zz_when_ArraySlice_l285_4_8 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l285_4_7 = {1'd0, _zz_when_ArraySlice_l285_4_8};
  assign _zz_when_ArraySlice_l288_4_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_4_2 = (_zz_when_ArraySlice_l288_4_3 + 8'h01);
  assign _zz_when_ArraySlice_l288_4_3 = (selectReadFifo_4 + _zz_when_ArraySlice_l288_4_4);
  assign _zz_when_ArraySlice_l288_4_5 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_4_4 = {1'd0, _zz_when_ArraySlice_l288_4_5};
  assign _zz_selectReadFifo_4_27 = (selectReadFifo_4 + _zz_selectReadFifo_4_28);
  assign _zz_selectReadFifo_4_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_4_28 = {1'd0, _zz_selectReadFifo_4_29};
  assign _zz_when_ArraySlice_l295_4 = (_zz_when_ArraySlice_l295_4_1 % aReg);
  assign _zz_when_ArraySlice_l295_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_4_1 = (_zz_when_ArraySlice_l306_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l306_4 = {5'd0, _zz_when_ArraySlice_l306_4_1};
  assign _zz_when_ArraySlice_l306_4_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_38 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_38_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_38_1 = (_zz_realValue1_0_38_2 + _zz_realValue1_0_38_3);
  assign _zz_realValue1_0_38_2 = {1'd0, hReg};
  assign _zz_realValue1_0_38_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_4_1 = (outSliceNumb_4_value + 7'h01);
  assign _zz_when_ArraySlice_l307_4 = {1'd0, _zz_when_ArraySlice_l307_4_1};
  assign _zz_when_ArraySlice_l307_4_2 = (realValue1_0_38 / aReg);
  assign _zz_selectReadFifo_4_30 = (selectReadFifo_4 - _zz_selectReadFifo_4_31);
  assign _zz_selectReadFifo_4_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_320 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_320_1);
  assign _zz_when_ArraySlice_l158_320_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_320_1 = {4'd0, _zz_when_ArraySlice_l158_320_2};
  assign _zz_when_ArraySlice_l158_320_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_320 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_320_1 = (_zz_when_ArraySlice_l159_320_2 - _zz_when_ArraySlice_l159_320_3);
  assign _zz_when_ArraySlice_l159_320_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_320_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_320_4);
  assign _zz_when_ArraySlice_l159_320_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_320_4 = {4'd0, _zz_when_ArraySlice_l159_320_5};
  assign _zz__zz_realValue_0_320 = {1'd0, wReg};
  assign _zz__zz_realValue_0_320_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_320_1 = (_zz_realValue_0_320_2 + _zz_realValue_0_320_3);
  assign _zz_realValue_0_320_2 = {1'd0, wReg};
  assign _zz_realValue_0_320_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_320 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_320_1 = (_zz_when_ArraySlice_l166_320_2 + _zz_when_ArraySlice_l166_320_6);
  assign _zz_when_ArraySlice_l166_320_2 = (realValue_0_320 - _zz_when_ArraySlice_l166_320_3);
  assign _zz_when_ArraySlice_l166_320_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_320_4);
  assign _zz_when_ArraySlice_l166_320_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_320_4 = {4'd0, _zz_when_ArraySlice_l166_320_5};
  assign _zz_when_ArraySlice_l166_320_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_321 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_321_1);
  assign _zz_when_ArraySlice_l158_321_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_321_1 = {3'd0, _zz_when_ArraySlice_l158_321_2};
  assign _zz_when_ArraySlice_l158_321_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_321_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_321 = {1'd0, _zz_when_ArraySlice_l159_321_1};
  assign _zz_when_ArraySlice_l159_321_2 = (_zz_when_ArraySlice_l159_321_3 - _zz_when_ArraySlice_l159_321_4);
  assign _zz_when_ArraySlice_l159_321_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_321_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_321_5);
  assign _zz_when_ArraySlice_l159_321_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_321_5 = {3'd0, _zz_when_ArraySlice_l159_321_6};
  assign _zz__zz_realValue_0_321 = {1'd0, wReg};
  assign _zz__zz_realValue_0_321_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_321_1 = (_zz_realValue_0_321_2 + _zz_realValue_0_321_3);
  assign _zz_realValue_0_321_2 = {1'd0, wReg};
  assign _zz_realValue_0_321_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_321_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_321 = {1'd0, _zz_when_ArraySlice_l166_321_1};
  assign _zz_when_ArraySlice_l166_321_2 = (_zz_when_ArraySlice_l166_321_3 + _zz_when_ArraySlice_l166_321_7);
  assign _zz_when_ArraySlice_l166_321_3 = (realValue_0_321 - _zz_when_ArraySlice_l166_321_4);
  assign _zz_when_ArraySlice_l166_321_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_321_5);
  assign _zz_when_ArraySlice_l166_321_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_321_5 = {3'd0, _zz_when_ArraySlice_l166_321_6};
  assign _zz_when_ArraySlice_l166_321_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_322 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_322_1);
  assign _zz_when_ArraySlice_l158_322_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_322_1 = {2'd0, _zz_when_ArraySlice_l158_322_2};
  assign _zz_when_ArraySlice_l158_322_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_322_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_322 = {1'd0, _zz_when_ArraySlice_l159_322_1};
  assign _zz_when_ArraySlice_l159_322_2 = (_zz_when_ArraySlice_l159_322_3 - _zz_when_ArraySlice_l159_322_4);
  assign _zz_when_ArraySlice_l159_322_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_322_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_322_5);
  assign _zz_when_ArraySlice_l159_322_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_322_5 = {2'd0, _zz_when_ArraySlice_l159_322_6};
  assign _zz__zz_realValue_0_322 = {1'd0, wReg};
  assign _zz__zz_realValue_0_322_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_322_1 = (_zz_realValue_0_322_2 + _zz_realValue_0_322_3);
  assign _zz_realValue_0_322_2 = {1'd0, wReg};
  assign _zz_realValue_0_322_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_322_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_322 = {1'd0, _zz_when_ArraySlice_l166_322_1};
  assign _zz_when_ArraySlice_l166_322_2 = (_zz_when_ArraySlice_l166_322_3 + _zz_when_ArraySlice_l166_322_7);
  assign _zz_when_ArraySlice_l166_322_3 = (realValue_0_322 - _zz_when_ArraySlice_l166_322_4);
  assign _zz_when_ArraySlice_l166_322_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_322_5);
  assign _zz_when_ArraySlice_l166_322_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_322_5 = {2'd0, _zz_when_ArraySlice_l166_322_6};
  assign _zz_when_ArraySlice_l166_322_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_323 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_323_1);
  assign _zz_when_ArraySlice_l158_323_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_323_1 = {2'd0, _zz_when_ArraySlice_l158_323_2};
  assign _zz_when_ArraySlice_l158_323_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_323_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_323 = {1'd0, _zz_when_ArraySlice_l159_323_1};
  assign _zz_when_ArraySlice_l159_323_2 = (_zz_when_ArraySlice_l159_323_3 - _zz_when_ArraySlice_l159_323_4);
  assign _zz_when_ArraySlice_l159_323_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_323_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_323_5);
  assign _zz_when_ArraySlice_l159_323_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_323_5 = {2'd0, _zz_when_ArraySlice_l159_323_6};
  assign _zz__zz_realValue_0_323 = {1'd0, wReg};
  assign _zz__zz_realValue_0_323_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_323_1 = (_zz_realValue_0_323_2 + _zz_realValue_0_323_3);
  assign _zz_realValue_0_323_2 = {1'd0, wReg};
  assign _zz_realValue_0_323_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_323_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_323 = {1'd0, _zz_when_ArraySlice_l166_323_1};
  assign _zz_when_ArraySlice_l166_323_2 = (_zz_when_ArraySlice_l166_323_3 + _zz_when_ArraySlice_l166_323_7);
  assign _zz_when_ArraySlice_l166_323_3 = (realValue_0_323 - _zz_when_ArraySlice_l166_323_4);
  assign _zz_when_ArraySlice_l166_323_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_323_5);
  assign _zz_when_ArraySlice_l166_323_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_323_5 = {2'd0, _zz_when_ArraySlice_l166_323_6};
  assign _zz_when_ArraySlice_l166_323_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_324 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_324_1);
  assign _zz_when_ArraySlice_l158_324_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_324_1 = {1'd0, _zz_when_ArraySlice_l158_324_2};
  assign _zz_when_ArraySlice_l158_324_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_324_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_324 = {1'd0, _zz_when_ArraySlice_l159_324_1};
  assign _zz_when_ArraySlice_l159_324_2 = (_zz_when_ArraySlice_l159_324_3 - _zz_when_ArraySlice_l159_324_4);
  assign _zz_when_ArraySlice_l159_324_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_324_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_324_5);
  assign _zz_when_ArraySlice_l159_324_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_324_5 = {1'd0, _zz_when_ArraySlice_l159_324_6};
  assign _zz__zz_realValue_0_324 = {1'd0, wReg};
  assign _zz__zz_realValue_0_324_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_324_1 = (_zz_realValue_0_324_2 + _zz_realValue_0_324_3);
  assign _zz_realValue_0_324_2 = {1'd0, wReg};
  assign _zz_realValue_0_324_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_324_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_324 = {1'd0, _zz_when_ArraySlice_l166_324_1};
  assign _zz_when_ArraySlice_l166_324_2 = (_zz_when_ArraySlice_l166_324_3 + _zz_when_ArraySlice_l166_324_7);
  assign _zz_when_ArraySlice_l166_324_3 = (realValue_0_324 - _zz_when_ArraySlice_l166_324_4);
  assign _zz_when_ArraySlice_l166_324_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_324_5);
  assign _zz_when_ArraySlice_l166_324_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_324_5 = {1'd0, _zz_when_ArraySlice_l166_324_6};
  assign _zz_when_ArraySlice_l166_324_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_325 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_325_1);
  assign _zz_when_ArraySlice_l158_325_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_325_1 = {1'd0, _zz_when_ArraySlice_l158_325_2};
  assign _zz_when_ArraySlice_l158_325_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_325_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_325 = {2'd0, _zz_when_ArraySlice_l159_325_1};
  assign _zz_when_ArraySlice_l159_325_2 = (_zz_when_ArraySlice_l159_325_3 - _zz_when_ArraySlice_l159_325_4);
  assign _zz_when_ArraySlice_l159_325_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_325_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_325_5);
  assign _zz_when_ArraySlice_l159_325_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_325_5 = {1'd0, _zz_when_ArraySlice_l159_325_6};
  assign _zz__zz_realValue_0_325 = {1'd0, wReg};
  assign _zz__zz_realValue_0_325_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_325_1 = (_zz_realValue_0_325_2 + _zz_realValue_0_325_3);
  assign _zz_realValue_0_325_2 = {1'd0, wReg};
  assign _zz_realValue_0_325_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_325_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_325 = {2'd0, _zz_when_ArraySlice_l166_325_1};
  assign _zz_when_ArraySlice_l166_325_2 = (_zz_when_ArraySlice_l166_325_3 + _zz_when_ArraySlice_l166_325_7);
  assign _zz_when_ArraySlice_l166_325_3 = (realValue_0_325 - _zz_when_ArraySlice_l166_325_4);
  assign _zz_when_ArraySlice_l166_325_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_325_5);
  assign _zz_when_ArraySlice_l166_325_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_325_5 = {1'd0, _zz_when_ArraySlice_l166_325_6};
  assign _zz_when_ArraySlice_l166_325_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_326 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_326_1);
  assign _zz_when_ArraySlice_l158_326_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_326_1 = {1'd0, _zz_when_ArraySlice_l158_326_2};
  assign _zz_when_ArraySlice_l158_326_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_326_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_326 = {2'd0, _zz_when_ArraySlice_l159_326_1};
  assign _zz_when_ArraySlice_l159_326_2 = (_zz_when_ArraySlice_l159_326_3 - _zz_when_ArraySlice_l159_326_4);
  assign _zz_when_ArraySlice_l159_326_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_326_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_326_5);
  assign _zz_when_ArraySlice_l159_326_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_326_5 = {1'd0, _zz_when_ArraySlice_l159_326_6};
  assign _zz__zz_realValue_0_326 = {1'd0, wReg};
  assign _zz__zz_realValue_0_326_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_326_1 = (_zz_realValue_0_326_2 + _zz_realValue_0_326_3);
  assign _zz_realValue_0_326_2 = {1'd0, wReg};
  assign _zz_realValue_0_326_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_326_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_326 = {2'd0, _zz_when_ArraySlice_l166_326_1};
  assign _zz_when_ArraySlice_l166_326_2 = (_zz_when_ArraySlice_l166_326_3 + _zz_when_ArraySlice_l166_326_7);
  assign _zz_when_ArraySlice_l166_326_3 = (realValue_0_326 - _zz_when_ArraySlice_l166_326_4);
  assign _zz_when_ArraySlice_l166_326_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_326_5);
  assign _zz_when_ArraySlice_l166_326_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_326_5 = {1'd0, _zz_when_ArraySlice_l166_326_6};
  assign _zz_when_ArraySlice_l166_326_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_327 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_327_1);
  assign _zz_when_ArraySlice_l158_327_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_327_1 = {1'd0, _zz_when_ArraySlice_l158_327_2};
  assign _zz_when_ArraySlice_l158_327_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_327_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_327 = {3'd0, _zz_when_ArraySlice_l159_327_1};
  assign _zz_when_ArraySlice_l159_327_2 = (_zz_when_ArraySlice_l159_327_3 - _zz_when_ArraySlice_l159_327_4);
  assign _zz_when_ArraySlice_l159_327_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_327_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_327_5);
  assign _zz_when_ArraySlice_l159_327_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_327_5 = {1'd0, _zz_when_ArraySlice_l159_327_6};
  assign _zz__zz_realValue_0_327 = {1'd0, wReg};
  assign _zz__zz_realValue_0_327_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_327_1 = (_zz_realValue_0_327_2 + _zz_realValue_0_327_3);
  assign _zz_realValue_0_327_2 = {1'd0, wReg};
  assign _zz_realValue_0_327_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_327_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_327 = {3'd0, _zz_when_ArraySlice_l166_327_1};
  assign _zz_when_ArraySlice_l166_327_2 = (_zz_when_ArraySlice_l166_327_3 + _zz_when_ArraySlice_l166_327_7);
  assign _zz_when_ArraySlice_l166_327_3 = (realValue_0_327 - _zz_when_ArraySlice_l166_327_4);
  assign _zz_when_ArraySlice_l166_327_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_327_5);
  assign _zz_when_ArraySlice_l166_327_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_327_5 = {1'd0, _zz_when_ArraySlice_l166_327_6};
  assign _zz_when_ArraySlice_l166_327_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_4 = (_zz_when_ArraySlice_l318_4_1 % aReg);
  assign _zz_when_ArraySlice_l318_4_1 = (handshakeTimes_4_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_4 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_4_1 = (selectReadFifo_4 + _zz_when_ArraySlice_l304_4_2);
  assign _zz_when_ArraySlice_l304_4_3 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l304_4_2 = {1'd0, _zz_when_ArraySlice_l304_4_3};
  assign _zz_when_ArraySlice_l325_4_1 = (_zz_when_ArraySlice_l325_4_2 - 8'h01);
  assign _zz_when_ArraySlice_l325_4 = {5'd0, _zz_when_ArraySlice_l325_4_1};
  assign _zz_when_ArraySlice_l325_4_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_5 = (selectReadFifo_5 + _zz_when_ArraySlice_l233_5_1);
  assign _zz_when_ArraySlice_l233_5_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l233_5_1 = {1'd0, _zz_when_ArraySlice_l233_5_2};
  assign _zz_when_ArraySlice_l233_5_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l234_5_3);
  assign _zz_when_ArraySlice_l234_5_1 = _zz_when_ArraySlice_l234_5_2[6:0];
  assign _zz_when_ArraySlice_l234_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l234_5_3 = {1'd0, _zz_when_ArraySlice_l234_5_4};
  assign _zz__zz_outputStreamArrayData_5_valid_1_2 = (bReg * 3'b101);
  assign _zz__zz_outputStreamArrayData_5_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_5_valid_1_2};
  assign _zz__zz_16 = _zz_outputStreamArrayData_5_valid_1[6:0];
  assign _zz_outputStreamArrayData_5_valid_5 = _zz_outputStreamArrayData_5_valid_1[6:0];
  assign _zz_outputStreamArrayData_5_payload_3 = _zz_outputStreamArrayData_5_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l240_5_3);
  assign _zz_when_ArraySlice_l240_5_1 = _zz_when_ArraySlice_l240_5_2[6:0];
  assign _zz_when_ArraySlice_l240_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l240_5_3 = {1'd0, _zz_when_ArraySlice_l240_5_4};
  assign _zz_when_ArraySlice_l241_5_1 = (_zz_when_ArraySlice_l241_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l241_5 = {5'd0, _zz_when_ArraySlice_l241_5_1};
  assign _zz_when_ArraySlice_l241_5_2 = (bReg * aReg);
  assign _zz_selectReadFifo_5_16 = (selectReadFifo_5 - _zz_selectReadFifo_5_17);
  assign _zz_selectReadFifo_5_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_5 = (_zz_when_ArraySlice_l244_5_1 % aReg);
  assign _zz_when_ArraySlice_l244_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l249_5_3);
  assign _zz_when_ArraySlice_l249_5_1 = _zz_when_ArraySlice_l249_5_2[6:0];
  assign _zz_when_ArraySlice_l249_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l249_5_3 = {1'd0, _zz_when_ArraySlice_l249_5_4};
  assign _zz_when_ArraySlice_l250_5_1 = (_zz_when_ArraySlice_l250_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l250_5 = {5'd0, _zz_when_ArraySlice_l250_5_1};
  assign _zz_when_ArraySlice_l250_5_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_39 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_39_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_39_1 = (_zz_realValue1_0_39_2 + _zz_realValue1_0_39_3);
  assign _zz_realValue1_0_39_2 = {1'd0, hReg};
  assign _zz_realValue1_0_39_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l252_5 = {1'd0, _zz_when_ArraySlice_l252_5_1};
  assign _zz_when_ArraySlice_l252_5_2 = (realValue1_0_39 / aReg);
  assign _zz_selectReadFifo_5_18 = (selectReadFifo_5 - _zz_selectReadFifo_5_19);
  assign _zz_selectReadFifo_5_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_5_21 = 1'b1;
  assign _zz_selectReadFifo_5_20 = {7'd0, _zz_selectReadFifo_5_21};
  assign _zz_when_ArraySlice_l158_328 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_328_1);
  assign _zz_when_ArraySlice_l158_328_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_328_1 = {4'd0, _zz_when_ArraySlice_l158_328_2};
  assign _zz_when_ArraySlice_l158_328_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_328 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_328_1 = (_zz_when_ArraySlice_l159_328_2 - _zz_when_ArraySlice_l159_328_3);
  assign _zz_when_ArraySlice_l159_328_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_328_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_328_4);
  assign _zz_when_ArraySlice_l159_328_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_328_4 = {4'd0, _zz_when_ArraySlice_l159_328_5};
  assign _zz__zz_realValue_0_328 = {1'd0, wReg};
  assign _zz__zz_realValue_0_328_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_328_1 = (_zz_realValue_0_328_2 + _zz_realValue_0_328_3);
  assign _zz_realValue_0_328_2 = {1'd0, wReg};
  assign _zz_realValue_0_328_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_328 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_328_1 = (_zz_when_ArraySlice_l166_328_2 + _zz_when_ArraySlice_l166_328_6);
  assign _zz_when_ArraySlice_l166_328_2 = (realValue_0_328 - _zz_when_ArraySlice_l166_328_3);
  assign _zz_when_ArraySlice_l166_328_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_328_4);
  assign _zz_when_ArraySlice_l166_328_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_328_4 = {4'd0, _zz_when_ArraySlice_l166_328_5};
  assign _zz_when_ArraySlice_l166_328_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_329 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_329_1);
  assign _zz_when_ArraySlice_l158_329_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_329_1 = {3'd0, _zz_when_ArraySlice_l158_329_2};
  assign _zz_when_ArraySlice_l158_329_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_329_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_329 = {1'd0, _zz_when_ArraySlice_l159_329_1};
  assign _zz_when_ArraySlice_l159_329_2 = (_zz_when_ArraySlice_l159_329_3 - _zz_when_ArraySlice_l159_329_4);
  assign _zz_when_ArraySlice_l159_329_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_329_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_329_5);
  assign _zz_when_ArraySlice_l159_329_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_329_5 = {3'd0, _zz_when_ArraySlice_l159_329_6};
  assign _zz__zz_realValue_0_329 = {1'd0, wReg};
  assign _zz__zz_realValue_0_329_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_329_1 = (_zz_realValue_0_329_2 + _zz_realValue_0_329_3);
  assign _zz_realValue_0_329_2 = {1'd0, wReg};
  assign _zz_realValue_0_329_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_329_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_329 = {1'd0, _zz_when_ArraySlice_l166_329_1};
  assign _zz_when_ArraySlice_l166_329_2 = (_zz_when_ArraySlice_l166_329_3 + _zz_when_ArraySlice_l166_329_7);
  assign _zz_when_ArraySlice_l166_329_3 = (realValue_0_329 - _zz_when_ArraySlice_l166_329_4);
  assign _zz_when_ArraySlice_l166_329_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_329_5);
  assign _zz_when_ArraySlice_l166_329_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_329_5 = {3'd0, _zz_when_ArraySlice_l166_329_6};
  assign _zz_when_ArraySlice_l166_329_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_330 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_330_1);
  assign _zz_when_ArraySlice_l158_330_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_330_1 = {2'd0, _zz_when_ArraySlice_l158_330_2};
  assign _zz_when_ArraySlice_l158_330_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_330_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_330 = {1'd0, _zz_when_ArraySlice_l159_330_1};
  assign _zz_when_ArraySlice_l159_330_2 = (_zz_when_ArraySlice_l159_330_3 - _zz_when_ArraySlice_l159_330_4);
  assign _zz_when_ArraySlice_l159_330_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_330_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_330_5);
  assign _zz_when_ArraySlice_l159_330_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_330_5 = {2'd0, _zz_when_ArraySlice_l159_330_6};
  assign _zz__zz_realValue_0_330 = {1'd0, wReg};
  assign _zz__zz_realValue_0_330_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_330_1 = (_zz_realValue_0_330_2 + _zz_realValue_0_330_3);
  assign _zz_realValue_0_330_2 = {1'd0, wReg};
  assign _zz_realValue_0_330_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_330_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_330 = {1'd0, _zz_when_ArraySlice_l166_330_1};
  assign _zz_when_ArraySlice_l166_330_2 = (_zz_when_ArraySlice_l166_330_3 + _zz_when_ArraySlice_l166_330_7);
  assign _zz_when_ArraySlice_l166_330_3 = (realValue_0_330 - _zz_when_ArraySlice_l166_330_4);
  assign _zz_when_ArraySlice_l166_330_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_330_5);
  assign _zz_when_ArraySlice_l166_330_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_330_5 = {2'd0, _zz_when_ArraySlice_l166_330_6};
  assign _zz_when_ArraySlice_l166_330_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_331 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_331_1);
  assign _zz_when_ArraySlice_l158_331_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_331_1 = {2'd0, _zz_when_ArraySlice_l158_331_2};
  assign _zz_when_ArraySlice_l158_331_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_331_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_331 = {1'd0, _zz_when_ArraySlice_l159_331_1};
  assign _zz_when_ArraySlice_l159_331_2 = (_zz_when_ArraySlice_l159_331_3 - _zz_when_ArraySlice_l159_331_4);
  assign _zz_when_ArraySlice_l159_331_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_331_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_331_5);
  assign _zz_when_ArraySlice_l159_331_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_331_5 = {2'd0, _zz_when_ArraySlice_l159_331_6};
  assign _zz__zz_realValue_0_331 = {1'd0, wReg};
  assign _zz__zz_realValue_0_331_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_331_1 = (_zz_realValue_0_331_2 + _zz_realValue_0_331_3);
  assign _zz_realValue_0_331_2 = {1'd0, wReg};
  assign _zz_realValue_0_331_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_331_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_331 = {1'd0, _zz_when_ArraySlice_l166_331_1};
  assign _zz_when_ArraySlice_l166_331_2 = (_zz_when_ArraySlice_l166_331_3 + _zz_when_ArraySlice_l166_331_7);
  assign _zz_when_ArraySlice_l166_331_3 = (realValue_0_331 - _zz_when_ArraySlice_l166_331_4);
  assign _zz_when_ArraySlice_l166_331_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_331_5);
  assign _zz_when_ArraySlice_l166_331_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_331_5 = {2'd0, _zz_when_ArraySlice_l166_331_6};
  assign _zz_when_ArraySlice_l166_331_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_332 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_332_1);
  assign _zz_when_ArraySlice_l158_332_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_332_1 = {1'd0, _zz_when_ArraySlice_l158_332_2};
  assign _zz_when_ArraySlice_l158_332_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_332_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_332 = {1'd0, _zz_when_ArraySlice_l159_332_1};
  assign _zz_when_ArraySlice_l159_332_2 = (_zz_when_ArraySlice_l159_332_3 - _zz_when_ArraySlice_l159_332_4);
  assign _zz_when_ArraySlice_l159_332_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_332_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_332_5);
  assign _zz_when_ArraySlice_l159_332_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_332_5 = {1'd0, _zz_when_ArraySlice_l159_332_6};
  assign _zz__zz_realValue_0_332 = {1'd0, wReg};
  assign _zz__zz_realValue_0_332_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_332_1 = (_zz_realValue_0_332_2 + _zz_realValue_0_332_3);
  assign _zz_realValue_0_332_2 = {1'd0, wReg};
  assign _zz_realValue_0_332_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_332_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_332 = {1'd0, _zz_when_ArraySlice_l166_332_1};
  assign _zz_when_ArraySlice_l166_332_2 = (_zz_when_ArraySlice_l166_332_3 + _zz_when_ArraySlice_l166_332_7);
  assign _zz_when_ArraySlice_l166_332_3 = (realValue_0_332 - _zz_when_ArraySlice_l166_332_4);
  assign _zz_when_ArraySlice_l166_332_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_332_5);
  assign _zz_when_ArraySlice_l166_332_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_332_5 = {1'd0, _zz_when_ArraySlice_l166_332_6};
  assign _zz_when_ArraySlice_l166_332_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_333 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_333_1);
  assign _zz_when_ArraySlice_l158_333_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_333_1 = {1'd0, _zz_when_ArraySlice_l158_333_2};
  assign _zz_when_ArraySlice_l158_333_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_333_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_333 = {2'd0, _zz_when_ArraySlice_l159_333_1};
  assign _zz_when_ArraySlice_l159_333_2 = (_zz_when_ArraySlice_l159_333_3 - _zz_when_ArraySlice_l159_333_4);
  assign _zz_when_ArraySlice_l159_333_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_333_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_333_5);
  assign _zz_when_ArraySlice_l159_333_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_333_5 = {1'd0, _zz_when_ArraySlice_l159_333_6};
  assign _zz__zz_realValue_0_333 = {1'd0, wReg};
  assign _zz__zz_realValue_0_333_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_333_1 = (_zz_realValue_0_333_2 + _zz_realValue_0_333_3);
  assign _zz_realValue_0_333_2 = {1'd0, wReg};
  assign _zz_realValue_0_333_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_333_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_333 = {2'd0, _zz_when_ArraySlice_l166_333_1};
  assign _zz_when_ArraySlice_l166_333_2 = (_zz_when_ArraySlice_l166_333_3 + _zz_when_ArraySlice_l166_333_7);
  assign _zz_when_ArraySlice_l166_333_3 = (realValue_0_333 - _zz_when_ArraySlice_l166_333_4);
  assign _zz_when_ArraySlice_l166_333_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_333_5);
  assign _zz_when_ArraySlice_l166_333_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_333_5 = {1'd0, _zz_when_ArraySlice_l166_333_6};
  assign _zz_when_ArraySlice_l166_333_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_334 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_334_1);
  assign _zz_when_ArraySlice_l158_334_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_334_1 = {1'd0, _zz_when_ArraySlice_l158_334_2};
  assign _zz_when_ArraySlice_l158_334_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_334_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_334 = {2'd0, _zz_when_ArraySlice_l159_334_1};
  assign _zz_when_ArraySlice_l159_334_2 = (_zz_when_ArraySlice_l159_334_3 - _zz_when_ArraySlice_l159_334_4);
  assign _zz_when_ArraySlice_l159_334_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_334_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_334_5);
  assign _zz_when_ArraySlice_l159_334_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_334_5 = {1'd0, _zz_when_ArraySlice_l159_334_6};
  assign _zz__zz_realValue_0_334 = {1'd0, wReg};
  assign _zz__zz_realValue_0_334_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_334_1 = (_zz_realValue_0_334_2 + _zz_realValue_0_334_3);
  assign _zz_realValue_0_334_2 = {1'd0, wReg};
  assign _zz_realValue_0_334_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_334_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_334 = {2'd0, _zz_when_ArraySlice_l166_334_1};
  assign _zz_when_ArraySlice_l166_334_2 = (_zz_when_ArraySlice_l166_334_3 + _zz_when_ArraySlice_l166_334_7);
  assign _zz_when_ArraySlice_l166_334_3 = (realValue_0_334 - _zz_when_ArraySlice_l166_334_4);
  assign _zz_when_ArraySlice_l166_334_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_334_5);
  assign _zz_when_ArraySlice_l166_334_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_334_5 = {1'd0, _zz_when_ArraySlice_l166_334_6};
  assign _zz_when_ArraySlice_l166_334_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_335 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_335_1);
  assign _zz_when_ArraySlice_l158_335_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_335_1 = {1'd0, _zz_when_ArraySlice_l158_335_2};
  assign _zz_when_ArraySlice_l158_335_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_335_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_335 = {3'd0, _zz_when_ArraySlice_l159_335_1};
  assign _zz_when_ArraySlice_l159_335_2 = (_zz_when_ArraySlice_l159_335_3 - _zz_when_ArraySlice_l159_335_4);
  assign _zz_when_ArraySlice_l159_335_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_335_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_335_5);
  assign _zz_when_ArraySlice_l159_335_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_335_5 = {1'd0, _zz_when_ArraySlice_l159_335_6};
  assign _zz__zz_realValue_0_335 = {1'd0, wReg};
  assign _zz__zz_realValue_0_335_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_335_1 = (_zz_realValue_0_335_2 + _zz_realValue_0_335_3);
  assign _zz_realValue_0_335_2 = {1'd0, wReg};
  assign _zz_realValue_0_335_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_335_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_335 = {3'd0, _zz_when_ArraySlice_l166_335_1};
  assign _zz_when_ArraySlice_l166_335_2 = (_zz_when_ArraySlice_l166_335_3 + _zz_when_ArraySlice_l166_335_7);
  assign _zz_when_ArraySlice_l166_335_3 = (realValue_0_335 - _zz_when_ArraySlice_l166_335_4);
  assign _zz_when_ArraySlice_l166_335_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_335_5);
  assign _zz_when_ArraySlice_l166_335_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_335_5 = {1'd0, _zz_when_ArraySlice_l166_335_6};
  assign _zz_when_ArraySlice_l166_335_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_5_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_5_2 = (_zz_when_ArraySlice_l260_5_3 + _zz_when_ArraySlice_l260_5_7);
  assign _zz_when_ArraySlice_l260_5_3 = (_zz_when_ArraySlice_l260_5_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l260_5_5);
  assign _zz_when_ArraySlice_l260_5_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_5_5 = {1'd0, _zz_when_ArraySlice_l260_5_6};
  assign _zz_when_ArraySlice_l260_5_8 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l260_5_7 = {1'd0, _zz_when_ArraySlice_l260_5_8};
  assign _zz_when_ArraySlice_l263_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_5_1 = (_zz_when_ArraySlice_l263_5_2 + 8'h01);
  assign _zz_when_ArraySlice_l263_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l263_5_3);
  assign _zz_when_ArraySlice_l263_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_5_3 = {1'd0, _zz_when_ArraySlice_l263_5_4};
  assign _zz_selectReadFifo_5_22 = (selectReadFifo_5 + _zz_selectReadFifo_5_23);
  assign _zz_selectReadFifo_5_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_23 = {1'd0, _zz_selectReadFifo_5_24};
  assign _zz_when_ArraySlice_l270_5 = (_zz_when_ArraySlice_l270_5_1 % aReg);
  assign _zz_when_ArraySlice_l270_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l274_5_3);
  assign _zz_when_ArraySlice_l274_5_1 = _zz_when_ArraySlice_l274_5_2[6:0];
  assign _zz_when_ArraySlice_l274_5_4 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l274_5_3 = {1'd0, _zz_when_ArraySlice_l274_5_4};
  assign _zz_when_ArraySlice_l275_5_1 = (_zz_when_ArraySlice_l275_5_2 - _zz_when_ArraySlice_l275_5_3);
  assign _zz_when_ArraySlice_l275_5 = {5'd0, _zz_when_ArraySlice_l275_5_1};
  assign _zz_when_ArraySlice_l275_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_5_4 = 1'b1;
  assign _zz_when_ArraySlice_l275_5_3 = {7'd0, _zz_when_ArraySlice_l275_5_4};
  assign _zz__zz_realValue1_0_40 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_40_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_40_1 = (_zz_realValue1_0_40_2 + _zz_realValue1_0_40_3);
  assign _zz_realValue1_0_40_2 = {1'd0, hReg};
  assign _zz_realValue1_0_40_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l277_5 = {1'd0, _zz_when_ArraySlice_l277_5_1};
  assign _zz_when_ArraySlice_l277_5_2 = (realValue1_0_40 / aReg);
  assign _zz_selectReadFifo_5_25 = (selectReadFifo_5 - _zz_selectReadFifo_5_26);
  assign _zz_selectReadFifo_5_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_336 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_336_1);
  assign _zz_when_ArraySlice_l158_336_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_336_1 = {4'd0, _zz_when_ArraySlice_l158_336_2};
  assign _zz_when_ArraySlice_l158_336_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_336 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_336_1 = (_zz_when_ArraySlice_l159_336_2 - _zz_when_ArraySlice_l159_336_3);
  assign _zz_when_ArraySlice_l159_336_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_336_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_336_4);
  assign _zz_when_ArraySlice_l159_336_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_336_4 = {4'd0, _zz_when_ArraySlice_l159_336_5};
  assign _zz__zz_realValue_0_336 = {1'd0, wReg};
  assign _zz__zz_realValue_0_336_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_336_1 = (_zz_realValue_0_336_2 + _zz_realValue_0_336_3);
  assign _zz_realValue_0_336_2 = {1'd0, wReg};
  assign _zz_realValue_0_336_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_336 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_336_1 = (_zz_when_ArraySlice_l166_336_2 + _zz_when_ArraySlice_l166_336_6);
  assign _zz_when_ArraySlice_l166_336_2 = (realValue_0_336 - _zz_when_ArraySlice_l166_336_3);
  assign _zz_when_ArraySlice_l166_336_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_336_4);
  assign _zz_when_ArraySlice_l166_336_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_336_4 = {4'd0, _zz_when_ArraySlice_l166_336_5};
  assign _zz_when_ArraySlice_l166_336_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_337 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_337_1);
  assign _zz_when_ArraySlice_l158_337_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_337_1 = {3'd0, _zz_when_ArraySlice_l158_337_2};
  assign _zz_when_ArraySlice_l158_337_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_337_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_337 = {1'd0, _zz_when_ArraySlice_l159_337_1};
  assign _zz_when_ArraySlice_l159_337_2 = (_zz_when_ArraySlice_l159_337_3 - _zz_when_ArraySlice_l159_337_4);
  assign _zz_when_ArraySlice_l159_337_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_337_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_337_5);
  assign _zz_when_ArraySlice_l159_337_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_337_5 = {3'd0, _zz_when_ArraySlice_l159_337_6};
  assign _zz__zz_realValue_0_337 = {1'd0, wReg};
  assign _zz__zz_realValue_0_337_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_337_1 = (_zz_realValue_0_337_2 + _zz_realValue_0_337_3);
  assign _zz_realValue_0_337_2 = {1'd0, wReg};
  assign _zz_realValue_0_337_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_337_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_337 = {1'd0, _zz_when_ArraySlice_l166_337_1};
  assign _zz_when_ArraySlice_l166_337_2 = (_zz_when_ArraySlice_l166_337_3 + _zz_when_ArraySlice_l166_337_7);
  assign _zz_when_ArraySlice_l166_337_3 = (realValue_0_337 - _zz_when_ArraySlice_l166_337_4);
  assign _zz_when_ArraySlice_l166_337_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_337_5);
  assign _zz_when_ArraySlice_l166_337_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_337_5 = {3'd0, _zz_when_ArraySlice_l166_337_6};
  assign _zz_when_ArraySlice_l166_337_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_338 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_338_1);
  assign _zz_when_ArraySlice_l158_338_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_338_1 = {2'd0, _zz_when_ArraySlice_l158_338_2};
  assign _zz_when_ArraySlice_l158_338_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_338_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_338 = {1'd0, _zz_when_ArraySlice_l159_338_1};
  assign _zz_when_ArraySlice_l159_338_2 = (_zz_when_ArraySlice_l159_338_3 - _zz_when_ArraySlice_l159_338_4);
  assign _zz_when_ArraySlice_l159_338_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_338_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_338_5);
  assign _zz_when_ArraySlice_l159_338_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_338_5 = {2'd0, _zz_when_ArraySlice_l159_338_6};
  assign _zz__zz_realValue_0_338 = {1'd0, wReg};
  assign _zz__zz_realValue_0_338_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_338_1 = (_zz_realValue_0_338_2 + _zz_realValue_0_338_3);
  assign _zz_realValue_0_338_2 = {1'd0, wReg};
  assign _zz_realValue_0_338_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_338_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_338 = {1'd0, _zz_when_ArraySlice_l166_338_1};
  assign _zz_when_ArraySlice_l166_338_2 = (_zz_when_ArraySlice_l166_338_3 + _zz_when_ArraySlice_l166_338_7);
  assign _zz_when_ArraySlice_l166_338_3 = (realValue_0_338 - _zz_when_ArraySlice_l166_338_4);
  assign _zz_when_ArraySlice_l166_338_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_338_5);
  assign _zz_when_ArraySlice_l166_338_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_338_5 = {2'd0, _zz_when_ArraySlice_l166_338_6};
  assign _zz_when_ArraySlice_l166_338_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_339 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_339_1);
  assign _zz_when_ArraySlice_l158_339_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_339_1 = {2'd0, _zz_when_ArraySlice_l158_339_2};
  assign _zz_when_ArraySlice_l158_339_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_339_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_339 = {1'd0, _zz_when_ArraySlice_l159_339_1};
  assign _zz_when_ArraySlice_l159_339_2 = (_zz_when_ArraySlice_l159_339_3 - _zz_when_ArraySlice_l159_339_4);
  assign _zz_when_ArraySlice_l159_339_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_339_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_339_5);
  assign _zz_when_ArraySlice_l159_339_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_339_5 = {2'd0, _zz_when_ArraySlice_l159_339_6};
  assign _zz__zz_realValue_0_339 = {1'd0, wReg};
  assign _zz__zz_realValue_0_339_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_339_1 = (_zz_realValue_0_339_2 + _zz_realValue_0_339_3);
  assign _zz_realValue_0_339_2 = {1'd0, wReg};
  assign _zz_realValue_0_339_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_339_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_339 = {1'd0, _zz_when_ArraySlice_l166_339_1};
  assign _zz_when_ArraySlice_l166_339_2 = (_zz_when_ArraySlice_l166_339_3 + _zz_when_ArraySlice_l166_339_7);
  assign _zz_when_ArraySlice_l166_339_3 = (realValue_0_339 - _zz_when_ArraySlice_l166_339_4);
  assign _zz_when_ArraySlice_l166_339_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_339_5);
  assign _zz_when_ArraySlice_l166_339_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_339_5 = {2'd0, _zz_when_ArraySlice_l166_339_6};
  assign _zz_when_ArraySlice_l166_339_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_340 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_340_1);
  assign _zz_when_ArraySlice_l158_340_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_340_1 = {1'd0, _zz_when_ArraySlice_l158_340_2};
  assign _zz_when_ArraySlice_l158_340_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_340_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_340 = {1'd0, _zz_when_ArraySlice_l159_340_1};
  assign _zz_when_ArraySlice_l159_340_2 = (_zz_when_ArraySlice_l159_340_3 - _zz_when_ArraySlice_l159_340_4);
  assign _zz_when_ArraySlice_l159_340_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_340_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_340_5);
  assign _zz_when_ArraySlice_l159_340_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_340_5 = {1'd0, _zz_when_ArraySlice_l159_340_6};
  assign _zz__zz_realValue_0_340 = {1'd0, wReg};
  assign _zz__zz_realValue_0_340_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_340_1 = (_zz_realValue_0_340_2 + _zz_realValue_0_340_3);
  assign _zz_realValue_0_340_2 = {1'd0, wReg};
  assign _zz_realValue_0_340_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_340_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_340 = {1'd0, _zz_when_ArraySlice_l166_340_1};
  assign _zz_when_ArraySlice_l166_340_2 = (_zz_when_ArraySlice_l166_340_3 + _zz_when_ArraySlice_l166_340_7);
  assign _zz_when_ArraySlice_l166_340_3 = (realValue_0_340 - _zz_when_ArraySlice_l166_340_4);
  assign _zz_when_ArraySlice_l166_340_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_340_5);
  assign _zz_when_ArraySlice_l166_340_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_340_5 = {1'd0, _zz_when_ArraySlice_l166_340_6};
  assign _zz_when_ArraySlice_l166_340_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_341 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_341_1);
  assign _zz_when_ArraySlice_l158_341_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_341_1 = {1'd0, _zz_when_ArraySlice_l158_341_2};
  assign _zz_when_ArraySlice_l158_341_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_341_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_341 = {2'd0, _zz_when_ArraySlice_l159_341_1};
  assign _zz_when_ArraySlice_l159_341_2 = (_zz_when_ArraySlice_l159_341_3 - _zz_when_ArraySlice_l159_341_4);
  assign _zz_when_ArraySlice_l159_341_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_341_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_341_5);
  assign _zz_when_ArraySlice_l159_341_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_341_5 = {1'd0, _zz_when_ArraySlice_l159_341_6};
  assign _zz__zz_realValue_0_341 = {1'd0, wReg};
  assign _zz__zz_realValue_0_341_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_341_1 = (_zz_realValue_0_341_2 + _zz_realValue_0_341_3);
  assign _zz_realValue_0_341_2 = {1'd0, wReg};
  assign _zz_realValue_0_341_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_341_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_341 = {2'd0, _zz_when_ArraySlice_l166_341_1};
  assign _zz_when_ArraySlice_l166_341_2 = (_zz_when_ArraySlice_l166_341_3 + _zz_when_ArraySlice_l166_341_7);
  assign _zz_when_ArraySlice_l166_341_3 = (realValue_0_341 - _zz_when_ArraySlice_l166_341_4);
  assign _zz_when_ArraySlice_l166_341_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_341_5);
  assign _zz_when_ArraySlice_l166_341_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_341_5 = {1'd0, _zz_when_ArraySlice_l166_341_6};
  assign _zz_when_ArraySlice_l166_341_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_342 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_342_1);
  assign _zz_when_ArraySlice_l158_342_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_342_1 = {1'd0, _zz_when_ArraySlice_l158_342_2};
  assign _zz_when_ArraySlice_l158_342_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_342_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_342 = {2'd0, _zz_when_ArraySlice_l159_342_1};
  assign _zz_when_ArraySlice_l159_342_2 = (_zz_when_ArraySlice_l159_342_3 - _zz_when_ArraySlice_l159_342_4);
  assign _zz_when_ArraySlice_l159_342_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_342_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_342_5);
  assign _zz_when_ArraySlice_l159_342_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_342_5 = {1'd0, _zz_when_ArraySlice_l159_342_6};
  assign _zz__zz_realValue_0_342 = {1'd0, wReg};
  assign _zz__zz_realValue_0_342_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_342_1 = (_zz_realValue_0_342_2 + _zz_realValue_0_342_3);
  assign _zz_realValue_0_342_2 = {1'd0, wReg};
  assign _zz_realValue_0_342_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_342_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_342 = {2'd0, _zz_when_ArraySlice_l166_342_1};
  assign _zz_when_ArraySlice_l166_342_2 = (_zz_when_ArraySlice_l166_342_3 + _zz_when_ArraySlice_l166_342_7);
  assign _zz_when_ArraySlice_l166_342_3 = (realValue_0_342 - _zz_when_ArraySlice_l166_342_4);
  assign _zz_when_ArraySlice_l166_342_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_342_5);
  assign _zz_when_ArraySlice_l166_342_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_342_5 = {1'd0, _zz_when_ArraySlice_l166_342_6};
  assign _zz_when_ArraySlice_l166_342_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_343 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_343_1);
  assign _zz_when_ArraySlice_l158_343_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_343_1 = {1'd0, _zz_when_ArraySlice_l158_343_2};
  assign _zz_when_ArraySlice_l158_343_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_343_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_343 = {3'd0, _zz_when_ArraySlice_l159_343_1};
  assign _zz_when_ArraySlice_l159_343_2 = (_zz_when_ArraySlice_l159_343_3 - _zz_when_ArraySlice_l159_343_4);
  assign _zz_when_ArraySlice_l159_343_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_343_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_343_5);
  assign _zz_when_ArraySlice_l159_343_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_343_5 = {1'd0, _zz_when_ArraySlice_l159_343_6};
  assign _zz__zz_realValue_0_343 = {1'd0, wReg};
  assign _zz__zz_realValue_0_343_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_343_1 = (_zz_realValue_0_343_2 + _zz_realValue_0_343_3);
  assign _zz_realValue_0_343_2 = {1'd0, wReg};
  assign _zz_realValue_0_343_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_343_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_343 = {3'd0, _zz_when_ArraySlice_l166_343_1};
  assign _zz_when_ArraySlice_l166_343_2 = (_zz_when_ArraySlice_l166_343_3 + _zz_when_ArraySlice_l166_343_7);
  assign _zz_when_ArraySlice_l166_343_3 = (realValue_0_343 - _zz_when_ArraySlice_l166_343_4);
  assign _zz_when_ArraySlice_l166_343_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_343_5);
  assign _zz_when_ArraySlice_l166_343_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_343_5 = {1'd0, _zz_when_ArraySlice_l166_343_6};
  assign _zz_when_ArraySlice_l166_343_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_5_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_5_2 = (_zz_when_ArraySlice_l285_5_3 + _zz_when_ArraySlice_l285_5_7);
  assign _zz_when_ArraySlice_l285_5_3 = (_zz_when_ArraySlice_l285_5_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_5_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l285_5_5);
  assign _zz_when_ArraySlice_l285_5_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_5_5 = {1'd0, _zz_when_ArraySlice_l285_5_6};
  assign _zz_when_ArraySlice_l285_5_8 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l285_5_7 = {1'd0, _zz_when_ArraySlice_l285_5_8};
  assign _zz_when_ArraySlice_l288_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_5_1 = (_zz_when_ArraySlice_l288_5_2 + 8'h01);
  assign _zz_when_ArraySlice_l288_5_2 = (selectReadFifo_5 + _zz_when_ArraySlice_l288_5_3);
  assign _zz_when_ArraySlice_l288_5_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_5_3 = {1'd0, _zz_when_ArraySlice_l288_5_4};
  assign _zz_selectReadFifo_5_27 = (selectReadFifo_5 + _zz_selectReadFifo_5_28);
  assign _zz_selectReadFifo_5_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_5_28 = {1'd0, _zz_selectReadFifo_5_29};
  assign _zz_when_ArraySlice_l295_5 = (_zz_when_ArraySlice_l295_5_1 % aReg);
  assign _zz_when_ArraySlice_l295_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_5_1 = (_zz_when_ArraySlice_l306_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l306_5 = {5'd0, _zz_when_ArraySlice_l306_5_1};
  assign _zz_when_ArraySlice_l306_5_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_41 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_41_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_41_1 = (_zz_realValue1_0_41_2 + _zz_realValue1_0_41_3);
  assign _zz_realValue1_0_41_2 = {1'd0, hReg};
  assign _zz_realValue1_0_41_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_5_1 = (outSliceNumb_5_value + 7'h01);
  assign _zz_when_ArraySlice_l307_5 = {1'd0, _zz_when_ArraySlice_l307_5_1};
  assign _zz_when_ArraySlice_l307_5_2 = (realValue1_0_41 / aReg);
  assign _zz_selectReadFifo_5_30 = (selectReadFifo_5 - _zz_selectReadFifo_5_31);
  assign _zz_selectReadFifo_5_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_344 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_344_1);
  assign _zz_when_ArraySlice_l158_344_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_344_1 = {4'd0, _zz_when_ArraySlice_l158_344_2};
  assign _zz_when_ArraySlice_l158_344_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_344 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_344_1 = (_zz_when_ArraySlice_l159_344_2 - _zz_when_ArraySlice_l159_344_3);
  assign _zz_when_ArraySlice_l159_344_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_344_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_344_4);
  assign _zz_when_ArraySlice_l159_344_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_344_4 = {4'd0, _zz_when_ArraySlice_l159_344_5};
  assign _zz__zz_realValue_0_344 = {1'd0, wReg};
  assign _zz__zz_realValue_0_344_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_344_1 = (_zz_realValue_0_344_2 + _zz_realValue_0_344_3);
  assign _zz_realValue_0_344_2 = {1'd0, wReg};
  assign _zz_realValue_0_344_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_344 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_344_1 = (_zz_when_ArraySlice_l166_344_2 + _zz_when_ArraySlice_l166_344_6);
  assign _zz_when_ArraySlice_l166_344_2 = (realValue_0_344 - _zz_when_ArraySlice_l166_344_3);
  assign _zz_when_ArraySlice_l166_344_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_344_4);
  assign _zz_when_ArraySlice_l166_344_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_344_4 = {4'd0, _zz_when_ArraySlice_l166_344_5};
  assign _zz_when_ArraySlice_l166_344_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_345 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_345_1);
  assign _zz_when_ArraySlice_l158_345_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_345_1 = {3'd0, _zz_when_ArraySlice_l158_345_2};
  assign _zz_when_ArraySlice_l158_345_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_345_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_345 = {1'd0, _zz_when_ArraySlice_l159_345_1};
  assign _zz_when_ArraySlice_l159_345_2 = (_zz_when_ArraySlice_l159_345_3 - _zz_when_ArraySlice_l159_345_4);
  assign _zz_when_ArraySlice_l159_345_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_345_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_345_5);
  assign _zz_when_ArraySlice_l159_345_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_345_5 = {3'd0, _zz_when_ArraySlice_l159_345_6};
  assign _zz__zz_realValue_0_345 = {1'd0, wReg};
  assign _zz__zz_realValue_0_345_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_345_1 = (_zz_realValue_0_345_2 + _zz_realValue_0_345_3);
  assign _zz_realValue_0_345_2 = {1'd0, wReg};
  assign _zz_realValue_0_345_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_345_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_345 = {1'd0, _zz_when_ArraySlice_l166_345_1};
  assign _zz_when_ArraySlice_l166_345_2 = (_zz_when_ArraySlice_l166_345_3 + _zz_when_ArraySlice_l166_345_7);
  assign _zz_when_ArraySlice_l166_345_3 = (realValue_0_345 - _zz_when_ArraySlice_l166_345_4);
  assign _zz_when_ArraySlice_l166_345_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_345_5);
  assign _zz_when_ArraySlice_l166_345_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_345_5 = {3'd0, _zz_when_ArraySlice_l166_345_6};
  assign _zz_when_ArraySlice_l166_345_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_346 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_346_1);
  assign _zz_when_ArraySlice_l158_346_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_346_1 = {2'd0, _zz_when_ArraySlice_l158_346_2};
  assign _zz_when_ArraySlice_l158_346_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_346_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_346 = {1'd0, _zz_when_ArraySlice_l159_346_1};
  assign _zz_when_ArraySlice_l159_346_2 = (_zz_when_ArraySlice_l159_346_3 - _zz_when_ArraySlice_l159_346_4);
  assign _zz_when_ArraySlice_l159_346_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_346_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_346_5);
  assign _zz_when_ArraySlice_l159_346_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_346_5 = {2'd0, _zz_when_ArraySlice_l159_346_6};
  assign _zz__zz_realValue_0_346 = {1'd0, wReg};
  assign _zz__zz_realValue_0_346_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_346_1 = (_zz_realValue_0_346_2 + _zz_realValue_0_346_3);
  assign _zz_realValue_0_346_2 = {1'd0, wReg};
  assign _zz_realValue_0_346_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_346_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_346 = {1'd0, _zz_when_ArraySlice_l166_346_1};
  assign _zz_when_ArraySlice_l166_346_2 = (_zz_when_ArraySlice_l166_346_3 + _zz_when_ArraySlice_l166_346_7);
  assign _zz_when_ArraySlice_l166_346_3 = (realValue_0_346 - _zz_when_ArraySlice_l166_346_4);
  assign _zz_when_ArraySlice_l166_346_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_346_5);
  assign _zz_when_ArraySlice_l166_346_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_346_5 = {2'd0, _zz_when_ArraySlice_l166_346_6};
  assign _zz_when_ArraySlice_l166_346_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_347 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_347_1);
  assign _zz_when_ArraySlice_l158_347_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_347_1 = {2'd0, _zz_when_ArraySlice_l158_347_2};
  assign _zz_when_ArraySlice_l158_347_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_347_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_347 = {1'd0, _zz_when_ArraySlice_l159_347_1};
  assign _zz_when_ArraySlice_l159_347_2 = (_zz_when_ArraySlice_l159_347_3 - _zz_when_ArraySlice_l159_347_4);
  assign _zz_when_ArraySlice_l159_347_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_347_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_347_5);
  assign _zz_when_ArraySlice_l159_347_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_347_5 = {2'd0, _zz_when_ArraySlice_l159_347_6};
  assign _zz__zz_realValue_0_347 = {1'd0, wReg};
  assign _zz__zz_realValue_0_347_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_347_1 = (_zz_realValue_0_347_2 + _zz_realValue_0_347_3);
  assign _zz_realValue_0_347_2 = {1'd0, wReg};
  assign _zz_realValue_0_347_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_347_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_347 = {1'd0, _zz_when_ArraySlice_l166_347_1};
  assign _zz_when_ArraySlice_l166_347_2 = (_zz_when_ArraySlice_l166_347_3 + _zz_when_ArraySlice_l166_347_7);
  assign _zz_when_ArraySlice_l166_347_3 = (realValue_0_347 - _zz_when_ArraySlice_l166_347_4);
  assign _zz_when_ArraySlice_l166_347_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_347_5);
  assign _zz_when_ArraySlice_l166_347_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_347_5 = {2'd0, _zz_when_ArraySlice_l166_347_6};
  assign _zz_when_ArraySlice_l166_347_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_348 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_348_1);
  assign _zz_when_ArraySlice_l158_348_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_348_1 = {1'd0, _zz_when_ArraySlice_l158_348_2};
  assign _zz_when_ArraySlice_l158_348_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_348_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_348 = {1'd0, _zz_when_ArraySlice_l159_348_1};
  assign _zz_when_ArraySlice_l159_348_2 = (_zz_when_ArraySlice_l159_348_3 - _zz_when_ArraySlice_l159_348_4);
  assign _zz_when_ArraySlice_l159_348_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_348_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_348_5);
  assign _zz_when_ArraySlice_l159_348_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_348_5 = {1'd0, _zz_when_ArraySlice_l159_348_6};
  assign _zz__zz_realValue_0_348 = {1'd0, wReg};
  assign _zz__zz_realValue_0_348_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_348_1 = (_zz_realValue_0_348_2 + _zz_realValue_0_348_3);
  assign _zz_realValue_0_348_2 = {1'd0, wReg};
  assign _zz_realValue_0_348_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_348_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_348 = {1'd0, _zz_when_ArraySlice_l166_348_1};
  assign _zz_when_ArraySlice_l166_348_2 = (_zz_when_ArraySlice_l166_348_3 + _zz_when_ArraySlice_l166_348_7);
  assign _zz_when_ArraySlice_l166_348_3 = (realValue_0_348 - _zz_when_ArraySlice_l166_348_4);
  assign _zz_when_ArraySlice_l166_348_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_348_5);
  assign _zz_when_ArraySlice_l166_348_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_348_5 = {1'd0, _zz_when_ArraySlice_l166_348_6};
  assign _zz_when_ArraySlice_l166_348_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_349 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_349_1);
  assign _zz_when_ArraySlice_l158_349_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_349_1 = {1'd0, _zz_when_ArraySlice_l158_349_2};
  assign _zz_when_ArraySlice_l158_349_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_349_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_349 = {2'd0, _zz_when_ArraySlice_l159_349_1};
  assign _zz_when_ArraySlice_l159_349_2 = (_zz_when_ArraySlice_l159_349_3 - _zz_when_ArraySlice_l159_349_4);
  assign _zz_when_ArraySlice_l159_349_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_349_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_349_5);
  assign _zz_when_ArraySlice_l159_349_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_349_5 = {1'd0, _zz_when_ArraySlice_l159_349_6};
  assign _zz__zz_realValue_0_349 = {1'd0, wReg};
  assign _zz__zz_realValue_0_349_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_349_1 = (_zz_realValue_0_349_2 + _zz_realValue_0_349_3);
  assign _zz_realValue_0_349_2 = {1'd0, wReg};
  assign _zz_realValue_0_349_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_349_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_349 = {2'd0, _zz_when_ArraySlice_l166_349_1};
  assign _zz_when_ArraySlice_l166_349_2 = (_zz_when_ArraySlice_l166_349_3 + _zz_when_ArraySlice_l166_349_7);
  assign _zz_when_ArraySlice_l166_349_3 = (realValue_0_349 - _zz_when_ArraySlice_l166_349_4);
  assign _zz_when_ArraySlice_l166_349_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_349_5);
  assign _zz_when_ArraySlice_l166_349_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_349_5 = {1'd0, _zz_when_ArraySlice_l166_349_6};
  assign _zz_when_ArraySlice_l166_349_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_350 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_350_1);
  assign _zz_when_ArraySlice_l158_350_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_350_1 = {1'd0, _zz_when_ArraySlice_l158_350_2};
  assign _zz_when_ArraySlice_l158_350_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_350_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_350 = {2'd0, _zz_when_ArraySlice_l159_350_1};
  assign _zz_when_ArraySlice_l159_350_2 = (_zz_when_ArraySlice_l159_350_3 - _zz_when_ArraySlice_l159_350_4);
  assign _zz_when_ArraySlice_l159_350_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_350_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_350_5);
  assign _zz_when_ArraySlice_l159_350_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_350_5 = {1'd0, _zz_when_ArraySlice_l159_350_6};
  assign _zz__zz_realValue_0_350 = {1'd0, wReg};
  assign _zz__zz_realValue_0_350_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_350_1 = (_zz_realValue_0_350_2 + _zz_realValue_0_350_3);
  assign _zz_realValue_0_350_2 = {1'd0, wReg};
  assign _zz_realValue_0_350_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_350_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_350 = {2'd0, _zz_when_ArraySlice_l166_350_1};
  assign _zz_when_ArraySlice_l166_350_2 = (_zz_when_ArraySlice_l166_350_3 + _zz_when_ArraySlice_l166_350_7);
  assign _zz_when_ArraySlice_l166_350_3 = (realValue_0_350 - _zz_when_ArraySlice_l166_350_4);
  assign _zz_when_ArraySlice_l166_350_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_350_5);
  assign _zz_when_ArraySlice_l166_350_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_350_5 = {1'd0, _zz_when_ArraySlice_l166_350_6};
  assign _zz_when_ArraySlice_l166_350_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_351 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_351_1);
  assign _zz_when_ArraySlice_l158_351_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_351_1 = {1'd0, _zz_when_ArraySlice_l158_351_2};
  assign _zz_when_ArraySlice_l158_351_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_351_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_351 = {3'd0, _zz_when_ArraySlice_l159_351_1};
  assign _zz_when_ArraySlice_l159_351_2 = (_zz_when_ArraySlice_l159_351_3 - _zz_when_ArraySlice_l159_351_4);
  assign _zz_when_ArraySlice_l159_351_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_351_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_351_5);
  assign _zz_when_ArraySlice_l159_351_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_351_5 = {1'd0, _zz_when_ArraySlice_l159_351_6};
  assign _zz__zz_realValue_0_351 = {1'd0, wReg};
  assign _zz__zz_realValue_0_351_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_351_1 = (_zz_realValue_0_351_2 + _zz_realValue_0_351_3);
  assign _zz_realValue_0_351_2 = {1'd0, wReg};
  assign _zz_realValue_0_351_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_351_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_351 = {3'd0, _zz_when_ArraySlice_l166_351_1};
  assign _zz_when_ArraySlice_l166_351_2 = (_zz_when_ArraySlice_l166_351_3 + _zz_when_ArraySlice_l166_351_7);
  assign _zz_when_ArraySlice_l166_351_3 = (realValue_0_351 - _zz_when_ArraySlice_l166_351_4);
  assign _zz_when_ArraySlice_l166_351_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_351_5);
  assign _zz_when_ArraySlice_l166_351_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_351_5 = {1'd0, _zz_when_ArraySlice_l166_351_6};
  assign _zz_when_ArraySlice_l166_351_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_5 = (_zz_when_ArraySlice_l318_5_1 % aReg);
  assign _zz_when_ArraySlice_l318_5_1 = (handshakeTimes_5_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_5 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_5_1 = (selectReadFifo_5 + _zz_when_ArraySlice_l304_5_2);
  assign _zz_when_ArraySlice_l304_5_3 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l304_5_2 = {1'd0, _zz_when_ArraySlice_l304_5_3};
  assign _zz_when_ArraySlice_l325_5_1 = (_zz_when_ArraySlice_l325_5_2 - 8'h01);
  assign _zz_when_ArraySlice_l325_5 = {5'd0, _zz_when_ArraySlice_l325_5_1};
  assign _zz_when_ArraySlice_l325_5_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_6 = (selectReadFifo_6 + _zz_when_ArraySlice_l233_6_1);
  assign _zz_when_ArraySlice_l233_6_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l233_6_1 = {1'd0, _zz_when_ArraySlice_l233_6_2};
  assign _zz_when_ArraySlice_l233_6_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l234_6_3);
  assign _zz_when_ArraySlice_l234_6_1 = _zz_when_ArraySlice_l234_6_2[6:0];
  assign _zz_when_ArraySlice_l234_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l234_6_3 = {1'd0, _zz_when_ArraySlice_l234_6_4};
  assign _zz__zz_outputStreamArrayData_6_valid_1_2 = (bReg * 3'b110);
  assign _zz__zz_outputStreamArrayData_6_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_6_valid_1_2};
  assign _zz__zz_17 = _zz_outputStreamArrayData_6_valid_1[6:0];
  assign _zz_outputStreamArrayData_6_valid_5 = _zz_outputStreamArrayData_6_valid_1[6:0];
  assign _zz_outputStreamArrayData_6_payload_3 = _zz_outputStreamArrayData_6_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l240_6_3);
  assign _zz_when_ArraySlice_l240_6_1 = _zz_when_ArraySlice_l240_6_2[6:0];
  assign _zz_when_ArraySlice_l240_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l240_6_3 = {1'd0, _zz_when_ArraySlice_l240_6_4};
  assign _zz_when_ArraySlice_l241_6_1 = (_zz_when_ArraySlice_l241_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l241_6 = {5'd0, _zz_when_ArraySlice_l241_6_1};
  assign _zz_when_ArraySlice_l241_6_2 = (bReg * aReg);
  assign _zz_selectReadFifo_6_16 = (selectReadFifo_6 - _zz_selectReadFifo_6_17);
  assign _zz_selectReadFifo_6_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_6 = (_zz_when_ArraySlice_l244_6_1 % aReg);
  assign _zz_when_ArraySlice_l244_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l249_6_3);
  assign _zz_when_ArraySlice_l249_6_1 = _zz_when_ArraySlice_l249_6_2[6:0];
  assign _zz_when_ArraySlice_l249_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l249_6_3 = {1'd0, _zz_when_ArraySlice_l249_6_4};
  assign _zz_when_ArraySlice_l250_6_1 = (_zz_when_ArraySlice_l250_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l250_6 = {5'd0, _zz_when_ArraySlice_l250_6_1};
  assign _zz_when_ArraySlice_l250_6_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_42 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_42_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_42_1 = (_zz_realValue1_0_42_2 + _zz_realValue1_0_42_3);
  assign _zz_realValue1_0_42_2 = {1'd0, hReg};
  assign _zz_realValue1_0_42_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l252_6 = {1'd0, _zz_when_ArraySlice_l252_6_1};
  assign _zz_when_ArraySlice_l252_6_2 = (realValue1_0_42 / aReg);
  assign _zz_selectReadFifo_6_18 = (selectReadFifo_6 - _zz_selectReadFifo_6_19);
  assign _zz_selectReadFifo_6_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_6_21 = 1'b1;
  assign _zz_selectReadFifo_6_20 = {7'd0, _zz_selectReadFifo_6_21};
  assign _zz_when_ArraySlice_l158_352 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_352_1);
  assign _zz_when_ArraySlice_l158_352_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_352_1 = {4'd0, _zz_when_ArraySlice_l158_352_2};
  assign _zz_when_ArraySlice_l158_352_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_352 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_352_1 = (_zz_when_ArraySlice_l159_352_2 - _zz_when_ArraySlice_l159_352_3);
  assign _zz_when_ArraySlice_l159_352_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_352_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_352_4);
  assign _zz_when_ArraySlice_l159_352_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_352_4 = {4'd0, _zz_when_ArraySlice_l159_352_5};
  assign _zz__zz_realValue_0_352 = {1'd0, wReg};
  assign _zz__zz_realValue_0_352_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_352_1 = (_zz_realValue_0_352_2 + _zz_realValue_0_352_3);
  assign _zz_realValue_0_352_2 = {1'd0, wReg};
  assign _zz_realValue_0_352_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_352 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_352_1 = (_zz_when_ArraySlice_l166_352_2 + _zz_when_ArraySlice_l166_352_6);
  assign _zz_when_ArraySlice_l166_352_2 = (realValue_0_352 - _zz_when_ArraySlice_l166_352_3);
  assign _zz_when_ArraySlice_l166_352_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_352_4);
  assign _zz_when_ArraySlice_l166_352_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_352_4 = {4'd0, _zz_when_ArraySlice_l166_352_5};
  assign _zz_when_ArraySlice_l166_352_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_353 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_353_1);
  assign _zz_when_ArraySlice_l158_353_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_353_1 = {3'd0, _zz_when_ArraySlice_l158_353_2};
  assign _zz_when_ArraySlice_l158_353_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_353_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_353 = {1'd0, _zz_when_ArraySlice_l159_353_1};
  assign _zz_when_ArraySlice_l159_353_2 = (_zz_when_ArraySlice_l159_353_3 - _zz_when_ArraySlice_l159_353_4);
  assign _zz_when_ArraySlice_l159_353_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_353_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_353_5);
  assign _zz_when_ArraySlice_l159_353_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_353_5 = {3'd0, _zz_when_ArraySlice_l159_353_6};
  assign _zz__zz_realValue_0_353 = {1'd0, wReg};
  assign _zz__zz_realValue_0_353_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_353_1 = (_zz_realValue_0_353_2 + _zz_realValue_0_353_3);
  assign _zz_realValue_0_353_2 = {1'd0, wReg};
  assign _zz_realValue_0_353_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_353_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_353 = {1'd0, _zz_when_ArraySlice_l166_353_1};
  assign _zz_when_ArraySlice_l166_353_2 = (_zz_when_ArraySlice_l166_353_3 + _zz_when_ArraySlice_l166_353_7);
  assign _zz_when_ArraySlice_l166_353_3 = (realValue_0_353 - _zz_when_ArraySlice_l166_353_4);
  assign _zz_when_ArraySlice_l166_353_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_353_5);
  assign _zz_when_ArraySlice_l166_353_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_353_5 = {3'd0, _zz_when_ArraySlice_l166_353_6};
  assign _zz_when_ArraySlice_l166_353_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_354 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_354_1);
  assign _zz_when_ArraySlice_l158_354_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_354_1 = {2'd0, _zz_when_ArraySlice_l158_354_2};
  assign _zz_when_ArraySlice_l158_354_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_354_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_354 = {1'd0, _zz_when_ArraySlice_l159_354_1};
  assign _zz_when_ArraySlice_l159_354_2 = (_zz_when_ArraySlice_l159_354_3 - _zz_when_ArraySlice_l159_354_4);
  assign _zz_when_ArraySlice_l159_354_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_354_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_354_5);
  assign _zz_when_ArraySlice_l159_354_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_354_5 = {2'd0, _zz_when_ArraySlice_l159_354_6};
  assign _zz__zz_realValue_0_354 = {1'd0, wReg};
  assign _zz__zz_realValue_0_354_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_354_1 = (_zz_realValue_0_354_2 + _zz_realValue_0_354_3);
  assign _zz_realValue_0_354_2 = {1'd0, wReg};
  assign _zz_realValue_0_354_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_354_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_354 = {1'd0, _zz_when_ArraySlice_l166_354_1};
  assign _zz_when_ArraySlice_l166_354_2 = (_zz_when_ArraySlice_l166_354_3 + _zz_when_ArraySlice_l166_354_7);
  assign _zz_when_ArraySlice_l166_354_3 = (realValue_0_354 - _zz_when_ArraySlice_l166_354_4);
  assign _zz_when_ArraySlice_l166_354_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_354_5);
  assign _zz_when_ArraySlice_l166_354_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_354_5 = {2'd0, _zz_when_ArraySlice_l166_354_6};
  assign _zz_when_ArraySlice_l166_354_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_355 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_355_1);
  assign _zz_when_ArraySlice_l158_355_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_355_1 = {2'd0, _zz_when_ArraySlice_l158_355_2};
  assign _zz_when_ArraySlice_l158_355_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_355_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_355 = {1'd0, _zz_when_ArraySlice_l159_355_1};
  assign _zz_when_ArraySlice_l159_355_2 = (_zz_when_ArraySlice_l159_355_3 - _zz_when_ArraySlice_l159_355_4);
  assign _zz_when_ArraySlice_l159_355_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_355_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_355_5);
  assign _zz_when_ArraySlice_l159_355_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_355_5 = {2'd0, _zz_when_ArraySlice_l159_355_6};
  assign _zz__zz_realValue_0_355 = {1'd0, wReg};
  assign _zz__zz_realValue_0_355_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_355_1 = (_zz_realValue_0_355_2 + _zz_realValue_0_355_3);
  assign _zz_realValue_0_355_2 = {1'd0, wReg};
  assign _zz_realValue_0_355_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_355_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_355 = {1'd0, _zz_when_ArraySlice_l166_355_1};
  assign _zz_when_ArraySlice_l166_355_2 = (_zz_when_ArraySlice_l166_355_3 + _zz_when_ArraySlice_l166_355_7);
  assign _zz_when_ArraySlice_l166_355_3 = (realValue_0_355 - _zz_when_ArraySlice_l166_355_4);
  assign _zz_when_ArraySlice_l166_355_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_355_5);
  assign _zz_when_ArraySlice_l166_355_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_355_5 = {2'd0, _zz_when_ArraySlice_l166_355_6};
  assign _zz_when_ArraySlice_l166_355_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_356 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_356_1);
  assign _zz_when_ArraySlice_l158_356_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_356_1 = {1'd0, _zz_when_ArraySlice_l158_356_2};
  assign _zz_when_ArraySlice_l158_356_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_356_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_356 = {1'd0, _zz_when_ArraySlice_l159_356_1};
  assign _zz_when_ArraySlice_l159_356_2 = (_zz_when_ArraySlice_l159_356_3 - _zz_when_ArraySlice_l159_356_4);
  assign _zz_when_ArraySlice_l159_356_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_356_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_356_5);
  assign _zz_when_ArraySlice_l159_356_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_356_5 = {1'd0, _zz_when_ArraySlice_l159_356_6};
  assign _zz__zz_realValue_0_356 = {1'd0, wReg};
  assign _zz__zz_realValue_0_356_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_356_1 = (_zz_realValue_0_356_2 + _zz_realValue_0_356_3);
  assign _zz_realValue_0_356_2 = {1'd0, wReg};
  assign _zz_realValue_0_356_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_356_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_356 = {1'd0, _zz_when_ArraySlice_l166_356_1};
  assign _zz_when_ArraySlice_l166_356_2 = (_zz_when_ArraySlice_l166_356_3 + _zz_when_ArraySlice_l166_356_7);
  assign _zz_when_ArraySlice_l166_356_3 = (realValue_0_356 - _zz_when_ArraySlice_l166_356_4);
  assign _zz_when_ArraySlice_l166_356_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_356_5);
  assign _zz_when_ArraySlice_l166_356_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_356_5 = {1'd0, _zz_when_ArraySlice_l166_356_6};
  assign _zz_when_ArraySlice_l166_356_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_357 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_357_1);
  assign _zz_when_ArraySlice_l158_357_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_357_1 = {1'd0, _zz_when_ArraySlice_l158_357_2};
  assign _zz_when_ArraySlice_l158_357_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_357_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_357 = {2'd0, _zz_when_ArraySlice_l159_357_1};
  assign _zz_when_ArraySlice_l159_357_2 = (_zz_when_ArraySlice_l159_357_3 - _zz_when_ArraySlice_l159_357_4);
  assign _zz_when_ArraySlice_l159_357_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_357_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_357_5);
  assign _zz_when_ArraySlice_l159_357_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_357_5 = {1'd0, _zz_when_ArraySlice_l159_357_6};
  assign _zz__zz_realValue_0_357 = {1'd0, wReg};
  assign _zz__zz_realValue_0_357_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_357_1 = (_zz_realValue_0_357_2 + _zz_realValue_0_357_3);
  assign _zz_realValue_0_357_2 = {1'd0, wReg};
  assign _zz_realValue_0_357_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_357_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_357 = {2'd0, _zz_when_ArraySlice_l166_357_1};
  assign _zz_when_ArraySlice_l166_357_2 = (_zz_when_ArraySlice_l166_357_3 + _zz_when_ArraySlice_l166_357_7);
  assign _zz_when_ArraySlice_l166_357_3 = (realValue_0_357 - _zz_when_ArraySlice_l166_357_4);
  assign _zz_when_ArraySlice_l166_357_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_357_5);
  assign _zz_when_ArraySlice_l166_357_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_357_5 = {1'd0, _zz_when_ArraySlice_l166_357_6};
  assign _zz_when_ArraySlice_l166_357_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_358 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_358_1);
  assign _zz_when_ArraySlice_l158_358_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_358_1 = {1'd0, _zz_when_ArraySlice_l158_358_2};
  assign _zz_when_ArraySlice_l158_358_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_358_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_358 = {2'd0, _zz_when_ArraySlice_l159_358_1};
  assign _zz_when_ArraySlice_l159_358_2 = (_zz_when_ArraySlice_l159_358_3 - _zz_when_ArraySlice_l159_358_4);
  assign _zz_when_ArraySlice_l159_358_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_358_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_358_5);
  assign _zz_when_ArraySlice_l159_358_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_358_5 = {1'd0, _zz_when_ArraySlice_l159_358_6};
  assign _zz__zz_realValue_0_358 = {1'd0, wReg};
  assign _zz__zz_realValue_0_358_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_358_1 = (_zz_realValue_0_358_2 + _zz_realValue_0_358_3);
  assign _zz_realValue_0_358_2 = {1'd0, wReg};
  assign _zz_realValue_0_358_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_358_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_358 = {2'd0, _zz_when_ArraySlice_l166_358_1};
  assign _zz_when_ArraySlice_l166_358_2 = (_zz_when_ArraySlice_l166_358_3 + _zz_when_ArraySlice_l166_358_7);
  assign _zz_when_ArraySlice_l166_358_3 = (realValue_0_358 - _zz_when_ArraySlice_l166_358_4);
  assign _zz_when_ArraySlice_l166_358_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_358_5);
  assign _zz_when_ArraySlice_l166_358_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_358_5 = {1'd0, _zz_when_ArraySlice_l166_358_6};
  assign _zz_when_ArraySlice_l166_358_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_359 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_359_1);
  assign _zz_when_ArraySlice_l158_359_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_359_1 = {1'd0, _zz_when_ArraySlice_l158_359_2};
  assign _zz_when_ArraySlice_l158_359_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_359_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_359 = {3'd0, _zz_when_ArraySlice_l159_359_1};
  assign _zz_when_ArraySlice_l159_359_2 = (_zz_when_ArraySlice_l159_359_3 - _zz_when_ArraySlice_l159_359_4);
  assign _zz_when_ArraySlice_l159_359_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_359_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_359_5);
  assign _zz_when_ArraySlice_l159_359_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_359_5 = {1'd0, _zz_when_ArraySlice_l159_359_6};
  assign _zz__zz_realValue_0_359 = {1'd0, wReg};
  assign _zz__zz_realValue_0_359_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_359_1 = (_zz_realValue_0_359_2 + _zz_realValue_0_359_3);
  assign _zz_realValue_0_359_2 = {1'd0, wReg};
  assign _zz_realValue_0_359_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_359_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_359 = {3'd0, _zz_when_ArraySlice_l166_359_1};
  assign _zz_when_ArraySlice_l166_359_2 = (_zz_when_ArraySlice_l166_359_3 + _zz_when_ArraySlice_l166_359_7);
  assign _zz_when_ArraySlice_l166_359_3 = (realValue_0_359 - _zz_when_ArraySlice_l166_359_4);
  assign _zz_when_ArraySlice_l166_359_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_359_5);
  assign _zz_when_ArraySlice_l166_359_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_359_5 = {1'd0, _zz_when_ArraySlice_l166_359_6};
  assign _zz_when_ArraySlice_l166_359_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_6_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_6_2 = (_zz_when_ArraySlice_l260_6_3 + _zz_when_ArraySlice_l260_6_7);
  assign _zz_when_ArraySlice_l260_6_3 = (_zz_when_ArraySlice_l260_6_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_6_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l260_6_5);
  assign _zz_when_ArraySlice_l260_6_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_6_5 = {1'd0, _zz_when_ArraySlice_l260_6_6};
  assign _zz_when_ArraySlice_l260_6_8 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l260_6_7 = {1'd0, _zz_when_ArraySlice_l260_6_8};
  assign _zz_when_ArraySlice_l263_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_6_1 = (_zz_when_ArraySlice_l263_6_2 + 8'h01);
  assign _zz_when_ArraySlice_l263_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l263_6_3);
  assign _zz_when_ArraySlice_l263_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_6_3 = {1'd0, _zz_when_ArraySlice_l263_6_4};
  assign _zz_selectReadFifo_6_22 = (selectReadFifo_6 + _zz_selectReadFifo_6_23);
  assign _zz_selectReadFifo_6_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_23 = {1'd0, _zz_selectReadFifo_6_24};
  assign _zz_when_ArraySlice_l270_6 = (_zz_when_ArraySlice_l270_6_1 % aReg);
  assign _zz_when_ArraySlice_l270_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l274_6_3);
  assign _zz_when_ArraySlice_l274_6_1 = _zz_when_ArraySlice_l274_6_2[6:0];
  assign _zz_when_ArraySlice_l274_6_4 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l274_6_3 = {1'd0, _zz_when_ArraySlice_l274_6_4};
  assign _zz_when_ArraySlice_l275_6_1 = (_zz_when_ArraySlice_l275_6_2 - _zz_when_ArraySlice_l275_6_3);
  assign _zz_when_ArraySlice_l275_6 = {5'd0, _zz_when_ArraySlice_l275_6_1};
  assign _zz_when_ArraySlice_l275_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_6_4 = 1'b1;
  assign _zz_when_ArraySlice_l275_6_3 = {7'd0, _zz_when_ArraySlice_l275_6_4};
  assign _zz__zz_realValue1_0_43 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_43_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_43_1 = (_zz_realValue1_0_43_2 + _zz_realValue1_0_43_3);
  assign _zz_realValue1_0_43_2 = {1'd0, hReg};
  assign _zz_realValue1_0_43_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l277_6 = {1'd0, _zz_when_ArraySlice_l277_6_1};
  assign _zz_when_ArraySlice_l277_6_2 = (realValue1_0_43 / aReg);
  assign _zz_selectReadFifo_6_25 = (selectReadFifo_6 - _zz_selectReadFifo_6_26);
  assign _zz_selectReadFifo_6_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_360 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_360_1);
  assign _zz_when_ArraySlice_l158_360_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_360_1 = {4'd0, _zz_when_ArraySlice_l158_360_2};
  assign _zz_when_ArraySlice_l158_360_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_360 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_360_1 = (_zz_when_ArraySlice_l159_360_2 - _zz_when_ArraySlice_l159_360_3);
  assign _zz_when_ArraySlice_l159_360_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_360_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_360_4);
  assign _zz_when_ArraySlice_l159_360_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_360_4 = {4'd0, _zz_when_ArraySlice_l159_360_5};
  assign _zz__zz_realValue_0_360 = {1'd0, wReg};
  assign _zz__zz_realValue_0_360_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_360_1 = (_zz_realValue_0_360_2 + _zz_realValue_0_360_3);
  assign _zz_realValue_0_360_2 = {1'd0, wReg};
  assign _zz_realValue_0_360_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_360 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_360_1 = (_zz_when_ArraySlice_l166_360_2 + _zz_when_ArraySlice_l166_360_6);
  assign _zz_when_ArraySlice_l166_360_2 = (realValue_0_360 - _zz_when_ArraySlice_l166_360_3);
  assign _zz_when_ArraySlice_l166_360_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_360_4);
  assign _zz_when_ArraySlice_l166_360_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_360_4 = {4'd0, _zz_when_ArraySlice_l166_360_5};
  assign _zz_when_ArraySlice_l166_360_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_361 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_361_1);
  assign _zz_when_ArraySlice_l158_361_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_361_1 = {3'd0, _zz_when_ArraySlice_l158_361_2};
  assign _zz_when_ArraySlice_l158_361_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_361_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_361 = {1'd0, _zz_when_ArraySlice_l159_361_1};
  assign _zz_when_ArraySlice_l159_361_2 = (_zz_when_ArraySlice_l159_361_3 - _zz_when_ArraySlice_l159_361_4);
  assign _zz_when_ArraySlice_l159_361_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_361_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_361_5);
  assign _zz_when_ArraySlice_l159_361_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_361_5 = {3'd0, _zz_when_ArraySlice_l159_361_6};
  assign _zz__zz_realValue_0_361 = {1'd0, wReg};
  assign _zz__zz_realValue_0_361_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_361_1 = (_zz_realValue_0_361_2 + _zz_realValue_0_361_3);
  assign _zz_realValue_0_361_2 = {1'd0, wReg};
  assign _zz_realValue_0_361_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_361_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_361 = {1'd0, _zz_when_ArraySlice_l166_361_1};
  assign _zz_when_ArraySlice_l166_361_2 = (_zz_when_ArraySlice_l166_361_3 + _zz_when_ArraySlice_l166_361_7);
  assign _zz_when_ArraySlice_l166_361_3 = (realValue_0_361 - _zz_when_ArraySlice_l166_361_4);
  assign _zz_when_ArraySlice_l166_361_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_361_5);
  assign _zz_when_ArraySlice_l166_361_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_361_5 = {3'd0, _zz_when_ArraySlice_l166_361_6};
  assign _zz_when_ArraySlice_l166_361_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_362 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_362_1);
  assign _zz_when_ArraySlice_l158_362_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_362_1 = {2'd0, _zz_when_ArraySlice_l158_362_2};
  assign _zz_when_ArraySlice_l158_362_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_362_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_362 = {1'd0, _zz_when_ArraySlice_l159_362_1};
  assign _zz_when_ArraySlice_l159_362_2 = (_zz_when_ArraySlice_l159_362_3 - _zz_when_ArraySlice_l159_362_4);
  assign _zz_when_ArraySlice_l159_362_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_362_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_362_5);
  assign _zz_when_ArraySlice_l159_362_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_362_5 = {2'd0, _zz_when_ArraySlice_l159_362_6};
  assign _zz__zz_realValue_0_362 = {1'd0, wReg};
  assign _zz__zz_realValue_0_362_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_362_1 = (_zz_realValue_0_362_2 + _zz_realValue_0_362_3);
  assign _zz_realValue_0_362_2 = {1'd0, wReg};
  assign _zz_realValue_0_362_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_362_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_362 = {1'd0, _zz_when_ArraySlice_l166_362_1};
  assign _zz_when_ArraySlice_l166_362_2 = (_zz_when_ArraySlice_l166_362_3 + _zz_when_ArraySlice_l166_362_7);
  assign _zz_when_ArraySlice_l166_362_3 = (realValue_0_362 - _zz_when_ArraySlice_l166_362_4);
  assign _zz_when_ArraySlice_l166_362_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_362_5);
  assign _zz_when_ArraySlice_l166_362_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_362_5 = {2'd0, _zz_when_ArraySlice_l166_362_6};
  assign _zz_when_ArraySlice_l166_362_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_363 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_363_1);
  assign _zz_when_ArraySlice_l158_363_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_363_1 = {2'd0, _zz_when_ArraySlice_l158_363_2};
  assign _zz_when_ArraySlice_l158_363_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_363_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_363 = {1'd0, _zz_when_ArraySlice_l159_363_1};
  assign _zz_when_ArraySlice_l159_363_2 = (_zz_when_ArraySlice_l159_363_3 - _zz_when_ArraySlice_l159_363_4);
  assign _zz_when_ArraySlice_l159_363_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_363_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_363_5);
  assign _zz_when_ArraySlice_l159_363_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_363_5 = {2'd0, _zz_when_ArraySlice_l159_363_6};
  assign _zz__zz_realValue_0_363 = {1'd0, wReg};
  assign _zz__zz_realValue_0_363_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_363_1 = (_zz_realValue_0_363_2 + _zz_realValue_0_363_3);
  assign _zz_realValue_0_363_2 = {1'd0, wReg};
  assign _zz_realValue_0_363_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_363_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_363 = {1'd0, _zz_when_ArraySlice_l166_363_1};
  assign _zz_when_ArraySlice_l166_363_2 = (_zz_when_ArraySlice_l166_363_3 + _zz_when_ArraySlice_l166_363_7);
  assign _zz_when_ArraySlice_l166_363_3 = (realValue_0_363 - _zz_when_ArraySlice_l166_363_4);
  assign _zz_when_ArraySlice_l166_363_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_363_5);
  assign _zz_when_ArraySlice_l166_363_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_363_5 = {2'd0, _zz_when_ArraySlice_l166_363_6};
  assign _zz_when_ArraySlice_l166_363_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_364 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_364_1);
  assign _zz_when_ArraySlice_l158_364_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_364_1 = {1'd0, _zz_when_ArraySlice_l158_364_2};
  assign _zz_when_ArraySlice_l158_364_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_364_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_364 = {1'd0, _zz_when_ArraySlice_l159_364_1};
  assign _zz_when_ArraySlice_l159_364_2 = (_zz_when_ArraySlice_l159_364_3 - _zz_when_ArraySlice_l159_364_4);
  assign _zz_when_ArraySlice_l159_364_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_364_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_364_5);
  assign _zz_when_ArraySlice_l159_364_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_364_5 = {1'd0, _zz_when_ArraySlice_l159_364_6};
  assign _zz__zz_realValue_0_364 = {1'd0, wReg};
  assign _zz__zz_realValue_0_364_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_364_1 = (_zz_realValue_0_364_2 + _zz_realValue_0_364_3);
  assign _zz_realValue_0_364_2 = {1'd0, wReg};
  assign _zz_realValue_0_364_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_364_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_364 = {1'd0, _zz_when_ArraySlice_l166_364_1};
  assign _zz_when_ArraySlice_l166_364_2 = (_zz_when_ArraySlice_l166_364_3 + _zz_when_ArraySlice_l166_364_7);
  assign _zz_when_ArraySlice_l166_364_3 = (realValue_0_364 - _zz_when_ArraySlice_l166_364_4);
  assign _zz_when_ArraySlice_l166_364_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_364_5);
  assign _zz_when_ArraySlice_l166_364_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_364_5 = {1'd0, _zz_when_ArraySlice_l166_364_6};
  assign _zz_when_ArraySlice_l166_364_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_365 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_365_1);
  assign _zz_when_ArraySlice_l158_365_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_365_1 = {1'd0, _zz_when_ArraySlice_l158_365_2};
  assign _zz_when_ArraySlice_l158_365_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_365_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_365 = {2'd0, _zz_when_ArraySlice_l159_365_1};
  assign _zz_when_ArraySlice_l159_365_2 = (_zz_when_ArraySlice_l159_365_3 - _zz_when_ArraySlice_l159_365_4);
  assign _zz_when_ArraySlice_l159_365_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_365_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_365_5);
  assign _zz_when_ArraySlice_l159_365_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_365_5 = {1'd0, _zz_when_ArraySlice_l159_365_6};
  assign _zz__zz_realValue_0_365 = {1'd0, wReg};
  assign _zz__zz_realValue_0_365_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_365_1 = (_zz_realValue_0_365_2 + _zz_realValue_0_365_3);
  assign _zz_realValue_0_365_2 = {1'd0, wReg};
  assign _zz_realValue_0_365_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_365_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_365 = {2'd0, _zz_when_ArraySlice_l166_365_1};
  assign _zz_when_ArraySlice_l166_365_2 = (_zz_when_ArraySlice_l166_365_3 + _zz_when_ArraySlice_l166_365_7);
  assign _zz_when_ArraySlice_l166_365_3 = (realValue_0_365 - _zz_when_ArraySlice_l166_365_4);
  assign _zz_when_ArraySlice_l166_365_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_365_5);
  assign _zz_when_ArraySlice_l166_365_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_365_5 = {1'd0, _zz_when_ArraySlice_l166_365_6};
  assign _zz_when_ArraySlice_l166_365_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_366 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_366_1);
  assign _zz_when_ArraySlice_l158_366_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_366_1 = {1'd0, _zz_when_ArraySlice_l158_366_2};
  assign _zz_when_ArraySlice_l158_366_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_366_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_366 = {2'd0, _zz_when_ArraySlice_l159_366_1};
  assign _zz_when_ArraySlice_l159_366_2 = (_zz_when_ArraySlice_l159_366_3 - _zz_when_ArraySlice_l159_366_4);
  assign _zz_when_ArraySlice_l159_366_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_366_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_366_5);
  assign _zz_when_ArraySlice_l159_366_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_366_5 = {1'd0, _zz_when_ArraySlice_l159_366_6};
  assign _zz__zz_realValue_0_366 = {1'd0, wReg};
  assign _zz__zz_realValue_0_366_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_366_1 = (_zz_realValue_0_366_2 + _zz_realValue_0_366_3);
  assign _zz_realValue_0_366_2 = {1'd0, wReg};
  assign _zz_realValue_0_366_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_366_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_366 = {2'd0, _zz_when_ArraySlice_l166_366_1};
  assign _zz_when_ArraySlice_l166_366_2 = (_zz_when_ArraySlice_l166_366_3 + _zz_when_ArraySlice_l166_366_7);
  assign _zz_when_ArraySlice_l166_366_3 = (realValue_0_366 - _zz_when_ArraySlice_l166_366_4);
  assign _zz_when_ArraySlice_l166_366_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_366_5);
  assign _zz_when_ArraySlice_l166_366_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_366_5 = {1'd0, _zz_when_ArraySlice_l166_366_6};
  assign _zz_when_ArraySlice_l166_366_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_367 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_367_1);
  assign _zz_when_ArraySlice_l158_367_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_367_1 = {1'd0, _zz_when_ArraySlice_l158_367_2};
  assign _zz_when_ArraySlice_l158_367_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_367_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_367 = {3'd0, _zz_when_ArraySlice_l159_367_1};
  assign _zz_when_ArraySlice_l159_367_2 = (_zz_when_ArraySlice_l159_367_3 - _zz_when_ArraySlice_l159_367_4);
  assign _zz_when_ArraySlice_l159_367_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_367_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_367_5);
  assign _zz_when_ArraySlice_l159_367_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_367_5 = {1'd0, _zz_when_ArraySlice_l159_367_6};
  assign _zz__zz_realValue_0_367 = {1'd0, wReg};
  assign _zz__zz_realValue_0_367_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_367_1 = (_zz_realValue_0_367_2 + _zz_realValue_0_367_3);
  assign _zz_realValue_0_367_2 = {1'd0, wReg};
  assign _zz_realValue_0_367_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_367_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_367 = {3'd0, _zz_when_ArraySlice_l166_367_1};
  assign _zz_when_ArraySlice_l166_367_2 = (_zz_when_ArraySlice_l166_367_3 + _zz_when_ArraySlice_l166_367_7);
  assign _zz_when_ArraySlice_l166_367_3 = (realValue_0_367 - _zz_when_ArraySlice_l166_367_4);
  assign _zz_when_ArraySlice_l166_367_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_367_5);
  assign _zz_when_ArraySlice_l166_367_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_367_5 = {1'd0, _zz_when_ArraySlice_l166_367_6};
  assign _zz_when_ArraySlice_l166_367_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_6_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_6_2 = (_zz_when_ArraySlice_l285_6_3 + _zz_when_ArraySlice_l285_6_7);
  assign _zz_when_ArraySlice_l285_6_3 = (_zz_when_ArraySlice_l285_6_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_6_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l285_6_5);
  assign _zz_when_ArraySlice_l285_6_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_6_5 = {1'd0, _zz_when_ArraySlice_l285_6_6};
  assign _zz_when_ArraySlice_l285_6_8 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l285_6_7 = {1'd0, _zz_when_ArraySlice_l285_6_8};
  assign _zz_when_ArraySlice_l288_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_6_1 = (_zz_when_ArraySlice_l288_6_2 + 8'h01);
  assign _zz_when_ArraySlice_l288_6_2 = (selectReadFifo_6 + _zz_when_ArraySlice_l288_6_3);
  assign _zz_when_ArraySlice_l288_6_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_6_3 = {1'd0, _zz_when_ArraySlice_l288_6_4};
  assign _zz_selectReadFifo_6_27 = (selectReadFifo_6 + _zz_selectReadFifo_6_28);
  assign _zz_selectReadFifo_6_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_6_28 = {1'd0, _zz_selectReadFifo_6_29};
  assign _zz_when_ArraySlice_l295_6 = (_zz_when_ArraySlice_l295_6_1 % aReg);
  assign _zz_when_ArraySlice_l295_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_6_1 = (_zz_when_ArraySlice_l306_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l306_6 = {5'd0, _zz_when_ArraySlice_l306_6_1};
  assign _zz_when_ArraySlice_l306_6_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_44 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_44_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_44_1 = (_zz_realValue1_0_44_2 + _zz_realValue1_0_44_3);
  assign _zz_realValue1_0_44_2 = {1'd0, hReg};
  assign _zz_realValue1_0_44_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_6_1 = (outSliceNumb_6_value + 7'h01);
  assign _zz_when_ArraySlice_l307_6 = {1'd0, _zz_when_ArraySlice_l307_6_1};
  assign _zz_when_ArraySlice_l307_6_2 = (realValue1_0_44 / aReg);
  assign _zz_selectReadFifo_6_30 = (selectReadFifo_6 - _zz_selectReadFifo_6_31);
  assign _zz_selectReadFifo_6_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_368 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_368_1);
  assign _zz_when_ArraySlice_l158_368_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_368_1 = {4'd0, _zz_when_ArraySlice_l158_368_2};
  assign _zz_when_ArraySlice_l158_368_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_368 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_368_1 = (_zz_when_ArraySlice_l159_368_2 - _zz_when_ArraySlice_l159_368_3);
  assign _zz_when_ArraySlice_l159_368_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_368_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_368_4);
  assign _zz_when_ArraySlice_l159_368_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_368_4 = {4'd0, _zz_when_ArraySlice_l159_368_5};
  assign _zz__zz_realValue_0_368 = {1'd0, wReg};
  assign _zz__zz_realValue_0_368_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_368_1 = (_zz_realValue_0_368_2 + _zz_realValue_0_368_3);
  assign _zz_realValue_0_368_2 = {1'd0, wReg};
  assign _zz_realValue_0_368_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_368 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_368_1 = (_zz_when_ArraySlice_l166_368_2 + _zz_when_ArraySlice_l166_368_6);
  assign _zz_when_ArraySlice_l166_368_2 = (realValue_0_368 - _zz_when_ArraySlice_l166_368_3);
  assign _zz_when_ArraySlice_l166_368_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_368_4);
  assign _zz_when_ArraySlice_l166_368_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_368_4 = {4'd0, _zz_when_ArraySlice_l166_368_5};
  assign _zz_when_ArraySlice_l166_368_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_369 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_369_1);
  assign _zz_when_ArraySlice_l158_369_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_369_1 = {3'd0, _zz_when_ArraySlice_l158_369_2};
  assign _zz_when_ArraySlice_l158_369_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_369_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_369 = {1'd0, _zz_when_ArraySlice_l159_369_1};
  assign _zz_when_ArraySlice_l159_369_2 = (_zz_when_ArraySlice_l159_369_3 - _zz_when_ArraySlice_l159_369_4);
  assign _zz_when_ArraySlice_l159_369_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_369_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_369_5);
  assign _zz_when_ArraySlice_l159_369_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_369_5 = {3'd0, _zz_when_ArraySlice_l159_369_6};
  assign _zz__zz_realValue_0_369 = {1'd0, wReg};
  assign _zz__zz_realValue_0_369_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_369_1 = (_zz_realValue_0_369_2 + _zz_realValue_0_369_3);
  assign _zz_realValue_0_369_2 = {1'd0, wReg};
  assign _zz_realValue_0_369_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_369_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_369 = {1'd0, _zz_when_ArraySlice_l166_369_1};
  assign _zz_when_ArraySlice_l166_369_2 = (_zz_when_ArraySlice_l166_369_3 + _zz_when_ArraySlice_l166_369_7);
  assign _zz_when_ArraySlice_l166_369_3 = (realValue_0_369 - _zz_when_ArraySlice_l166_369_4);
  assign _zz_when_ArraySlice_l166_369_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_369_5);
  assign _zz_when_ArraySlice_l166_369_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_369_5 = {3'd0, _zz_when_ArraySlice_l166_369_6};
  assign _zz_when_ArraySlice_l166_369_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_370 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_370_1);
  assign _zz_when_ArraySlice_l158_370_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_370_1 = {2'd0, _zz_when_ArraySlice_l158_370_2};
  assign _zz_when_ArraySlice_l158_370_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_370_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_370 = {1'd0, _zz_when_ArraySlice_l159_370_1};
  assign _zz_when_ArraySlice_l159_370_2 = (_zz_when_ArraySlice_l159_370_3 - _zz_when_ArraySlice_l159_370_4);
  assign _zz_when_ArraySlice_l159_370_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_370_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_370_5);
  assign _zz_when_ArraySlice_l159_370_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_370_5 = {2'd0, _zz_when_ArraySlice_l159_370_6};
  assign _zz__zz_realValue_0_370 = {1'd0, wReg};
  assign _zz__zz_realValue_0_370_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_370_1 = (_zz_realValue_0_370_2 + _zz_realValue_0_370_3);
  assign _zz_realValue_0_370_2 = {1'd0, wReg};
  assign _zz_realValue_0_370_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_370_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_370 = {1'd0, _zz_when_ArraySlice_l166_370_1};
  assign _zz_when_ArraySlice_l166_370_2 = (_zz_when_ArraySlice_l166_370_3 + _zz_when_ArraySlice_l166_370_7);
  assign _zz_when_ArraySlice_l166_370_3 = (realValue_0_370 - _zz_when_ArraySlice_l166_370_4);
  assign _zz_when_ArraySlice_l166_370_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_370_5);
  assign _zz_when_ArraySlice_l166_370_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_370_5 = {2'd0, _zz_when_ArraySlice_l166_370_6};
  assign _zz_when_ArraySlice_l166_370_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_371 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_371_1);
  assign _zz_when_ArraySlice_l158_371_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_371_1 = {2'd0, _zz_when_ArraySlice_l158_371_2};
  assign _zz_when_ArraySlice_l158_371_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_371_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_371 = {1'd0, _zz_when_ArraySlice_l159_371_1};
  assign _zz_when_ArraySlice_l159_371_2 = (_zz_when_ArraySlice_l159_371_3 - _zz_when_ArraySlice_l159_371_4);
  assign _zz_when_ArraySlice_l159_371_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_371_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_371_5);
  assign _zz_when_ArraySlice_l159_371_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_371_5 = {2'd0, _zz_when_ArraySlice_l159_371_6};
  assign _zz__zz_realValue_0_371 = {1'd0, wReg};
  assign _zz__zz_realValue_0_371_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_371_1 = (_zz_realValue_0_371_2 + _zz_realValue_0_371_3);
  assign _zz_realValue_0_371_2 = {1'd0, wReg};
  assign _zz_realValue_0_371_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_371_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_371 = {1'd0, _zz_when_ArraySlice_l166_371_1};
  assign _zz_when_ArraySlice_l166_371_2 = (_zz_when_ArraySlice_l166_371_3 + _zz_when_ArraySlice_l166_371_7);
  assign _zz_when_ArraySlice_l166_371_3 = (realValue_0_371 - _zz_when_ArraySlice_l166_371_4);
  assign _zz_when_ArraySlice_l166_371_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_371_5);
  assign _zz_when_ArraySlice_l166_371_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_371_5 = {2'd0, _zz_when_ArraySlice_l166_371_6};
  assign _zz_when_ArraySlice_l166_371_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_372 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_372_1);
  assign _zz_when_ArraySlice_l158_372_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_372_1 = {1'd0, _zz_when_ArraySlice_l158_372_2};
  assign _zz_when_ArraySlice_l158_372_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_372_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_372 = {1'd0, _zz_when_ArraySlice_l159_372_1};
  assign _zz_when_ArraySlice_l159_372_2 = (_zz_when_ArraySlice_l159_372_3 - _zz_when_ArraySlice_l159_372_4);
  assign _zz_when_ArraySlice_l159_372_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_372_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_372_5);
  assign _zz_when_ArraySlice_l159_372_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_372_5 = {1'd0, _zz_when_ArraySlice_l159_372_6};
  assign _zz__zz_realValue_0_372 = {1'd0, wReg};
  assign _zz__zz_realValue_0_372_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_372_1 = (_zz_realValue_0_372_2 + _zz_realValue_0_372_3);
  assign _zz_realValue_0_372_2 = {1'd0, wReg};
  assign _zz_realValue_0_372_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_372_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_372 = {1'd0, _zz_when_ArraySlice_l166_372_1};
  assign _zz_when_ArraySlice_l166_372_2 = (_zz_when_ArraySlice_l166_372_3 + _zz_when_ArraySlice_l166_372_7);
  assign _zz_when_ArraySlice_l166_372_3 = (realValue_0_372 - _zz_when_ArraySlice_l166_372_4);
  assign _zz_when_ArraySlice_l166_372_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_372_5);
  assign _zz_when_ArraySlice_l166_372_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_372_5 = {1'd0, _zz_when_ArraySlice_l166_372_6};
  assign _zz_when_ArraySlice_l166_372_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_373 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_373_1);
  assign _zz_when_ArraySlice_l158_373_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_373_1 = {1'd0, _zz_when_ArraySlice_l158_373_2};
  assign _zz_when_ArraySlice_l158_373_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_373_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_373 = {2'd0, _zz_when_ArraySlice_l159_373_1};
  assign _zz_when_ArraySlice_l159_373_2 = (_zz_when_ArraySlice_l159_373_3 - _zz_when_ArraySlice_l159_373_4);
  assign _zz_when_ArraySlice_l159_373_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_373_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_373_5);
  assign _zz_when_ArraySlice_l159_373_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_373_5 = {1'd0, _zz_when_ArraySlice_l159_373_6};
  assign _zz__zz_realValue_0_373 = {1'd0, wReg};
  assign _zz__zz_realValue_0_373_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_373_1 = (_zz_realValue_0_373_2 + _zz_realValue_0_373_3);
  assign _zz_realValue_0_373_2 = {1'd0, wReg};
  assign _zz_realValue_0_373_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_373_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_373 = {2'd0, _zz_when_ArraySlice_l166_373_1};
  assign _zz_when_ArraySlice_l166_373_2 = (_zz_when_ArraySlice_l166_373_3 + _zz_when_ArraySlice_l166_373_7);
  assign _zz_when_ArraySlice_l166_373_3 = (realValue_0_373 - _zz_when_ArraySlice_l166_373_4);
  assign _zz_when_ArraySlice_l166_373_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_373_5);
  assign _zz_when_ArraySlice_l166_373_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_373_5 = {1'd0, _zz_when_ArraySlice_l166_373_6};
  assign _zz_when_ArraySlice_l166_373_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_374 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_374_1);
  assign _zz_when_ArraySlice_l158_374_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_374_1 = {1'd0, _zz_when_ArraySlice_l158_374_2};
  assign _zz_when_ArraySlice_l158_374_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_374_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_374 = {2'd0, _zz_when_ArraySlice_l159_374_1};
  assign _zz_when_ArraySlice_l159_374_2 = (_zz_when_ArraySlice_l159_374_3 - _zz_when_ArraySlice_l159_374_4);
  assign _zz_when_ArraySlice_l159_374_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_374_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_374_5);
  assign _zz_when_ArraySlice_l159_374_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_374_5 = {1'd0, _zz_when_ArraySlice_l159_374_6};
  assign _zz__zz_realValue_0_374 = {1'd0, wReg};
  assign _zz__zz_realValue_0_374_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_374_1 = (_zz_realValue_0_374_2 + _zz_realValue_0_374_3);
  assign _zz_realValue_0_374_2 = {1'd0, wReg};
  assign _zz_realValue_0_374_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_374_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_374 = {2'd0, _zz_when_ArraySlice_l166_374_1};
  assign _zz_when_ArraySlice_l166_374_2 = (_zz_when_ArraySlice_l166_374_3 + _zz_when_ArraySlice_l166_374_7);
  assign _zz_when_ArraySlice_l166_374_3 = (realValue_0_374 - _zz_when_ArraySlice_l166_374_4);
  assign _zz_when_ArraySlice_l166_374_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_374_5);
  assign _zz_when_ArraySlice_l166_374_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_374_5 = {1'd0, _zz_when_ArraySlice_l166_374_6};
  assign _zz_when_ArraySlice_l166_374_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_375 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_375_1);
  assign _zz_when_ArraySlice_l158_375_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_375_1 = {1'd0, _zz_when_ArraySlice_l158_375_2};
  assign _zz_when_ArraySlice_l158_375_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_375_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_375 = {3'd0, _zz_when_ArraySlice_l159_375_1};
  assign _zz_when_ArraySlice_l159_375_2 = (_zz_when_ArraySlice_l159_375_3 - _zz_when_ArraySlice_l159_375_4);
  assign _zz_when_ArraySlice_l159_375_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_375_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_375_5);
  assign _zz_when_ArraySlice_l159_375_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_375_5 = {1'd0, _zz_when_ArraySlice_l159_375_6};
  assign _zz__zz_realValue_0_375 = {1'd0, wReg};
  assign _zz__zz_realValue_0_375_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_375_1 = (_zz_realValue_0_375_2 + _zz_realValue_0_375_3);
  assign _zz_realValue_0_375_2 = {1'd0, wReg};
  assign _zz_realValue_0_375_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_375_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_375 = {3'd0, _zz_when_ArraySlice_l166_375_1};
  assign _zz_when_ArraySlice_l166_375_2 = (_zz_when_ArraySlice_l166_375_3 + _zz_when_ArraySlice_l166_375_7);
  assign _zz_when_ArraySlice_l166_375_3 = (realValue_0_375 - _zz_when_ArraySlice_l166_375_4);
  assign _zz_when_ArraySlice_l166_375_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_375_5);
  assign _zz_when_ArraySlice_l166_375_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_375_5 = {1'd0, _zz_when_ArraySlice_l166_375_6};
  assign _zz_when_ArraySlice_l166_375_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_6 = (_zz_when_ArraySlice_l318_6_1 % aReg);
  assign _zz_when_ArraySlice_l318_6_1 = (handshakeTimes_6_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_6 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_6_1 = (selectReadFifo_6 + _zz_when_ArraySlice_l304_6_2);
  assign _zz_when_ArraySlice_l304_6_3 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l304_6_2 = {1'd0, _zz_when_ArraySlice_l304_6_3};
  assign _zz_when_ArraySlice_l325_6_1 = (_zz_when_ArraySlice_l325_6_2 - 8'h01);
  assign _zz_when_ArraySlice_l325_6 = {5'd0, _zz_when_ArraySlice_l325_6_1};
  assign _zz_when_ArraySlice_l325_6_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l233_7 = (selectReadFifo_7 + _zz_when_ArraySlice_l233_7_1);
  assign _zz_when_ArraySlice_l233_7_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l233_7_1 = {1'd0, _zz_when_ArraySlice_l233_7_2};
  assign _zz_when_ArraySlice_l233_7_3 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l234_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l234_7_3);
  assign _zz_when_ArraySlice_l234_7_1 = _zz_when_ArraySlice_l234_7_2[6:0];
  assign _zz_when_ArraySlice_l234_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l234_7_3 = {1'd0, _zz_when_ArraySlice_l234_7_4};
  assign _zz__zz_outputStreamArrayData_7_valid_1_2 = (bReg * 3'b111);
  assign _zz__zz_outputStreamArrayData_7_valid_1_1 = {1'd0, _zz__zz_outputStreamArrayData_7_valid_1_2};
  assign _zz__zz_18 = _zz_outputStreamArrayData_7_valid_1[6:0];
  assign _zz_outputStreamArrayData_7_valid_5 = _zz_outputStreamArrayData_7_valid_1[6:0];
  assign _zz_outputStreamArrayData_7_payload_3 = _zz_outputStreamArrayData_7_valid_1[6:0];
  assign _zz_when_ArraySlice_l240_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l240_7_3);
  assign _zz_when_ArraySlice_l240_7_1 = _zz_when_ArraySlice_l240_7_2[6:0];
  assign _zz_when_ArraySlice_l240_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l240_7_3 = {1'd0, _zz_when_ArraySlice_l240_7_4};
  assign _zz_when_ArraySlice_l241_7_1 = (_zz_when_ArraySlice_l241_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l241_7 = {5'd0, _zz_when_ArraySlice_l241_7_1};
  assign _zz_when_ArraySlice_l241_7_2 = (bReg * aReg);
  assign _zz_selectReadFifo_7_16 = (selectReadFifo_7 - _zz_selectReadFifo_7_17);
  assign _zz_selectReadFifo_7_17 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l244_7 = (_zz_when_ArraySlice_l244_7_1 % aReg);
  assign _zz_when_ArraySlice_l244_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l249_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l249_7_3);
  assign _zz_when_ArraySlice_l249_7_1 = _zz_when_ArraySlice_l249_7_2[6:0];
  assign _zz_when_ArraySlice_l249_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l249_7_3 = {1'd0, _zz_when_ArraySlice_l249_7_4};
  assign _zz_when_ArraySlice_l250_7_1 = (_zz_when_ArraySlice_l250_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l250_7 = {5'd0, _zz_when_ArraySlice_l250_7_1};
  assign _zz_when_ArraySlice_l250_7_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_45 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_45_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_45_1 = (_zz_realValue1_0_45_2 + _zz_realValue1_0_45_3);
  assign _zz_realValue1_0_45_2 = {1'd0, hReg};
  assign _zz_realValue1_0_45_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l252_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l252_7 = {1'd0, _zz_when_ArraySlice_l252_7_1};
  assign _zz_when_ArraySlice_l252_7_2 = (realValue1_0_45 / aReg);
  assign _zz_selectReadFifo_7_18 = (selectReadFifo_7 - _zz_selectReadFifo_7_19);
  assign _zz_selectReadFifo_7_19 = {4'd0, bReg};
  assign _zz_selectReadFifo_7_21 = 1'b1;
  assign _zz_selectReadFifo_7_20 = {7'd0, _zz_selectReadFifo_7_21};
  assign _zz_when_ArraySlice_l158_376 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_376_1);
  assign _zz_when_ArraySlice_l158_376_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_376_1 = {4'd0, _zz_when_ArraySlice_l158_376_2};
  assign _zz_when_ArraySlice_l158_376_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_376 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_376_1 = (_zz_when_ArraySlice_l159_376_2 - _zz_when_ArraySlice_l159_376_3);
  assign _zz_when_ArraySlice_l159_376_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_376_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_376_4);
  assign _zz_when_ArraySlice_l159_376_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_376_4 = {4'd0, _zz_when_ArraySlice_l159_376_5};
  assign _zz__zz_realValue_0_376 = {1'd0, wReg};
  assign _zz__zz_realValue_0_376_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_376_1 = (_zz_realValue_0_376_2 + _zz_realValue_0_376_3);
  assign _zz_realValue_0_376_2 = {1'd0, wReg};
  assign _zz_realValue_0_376_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_376 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_376_1 = (_zz_when_ArraySlice_l166_376_2 + _zz_when_ArraySlice_l166_376_6);
  assign _zz_when_ArraySlice_l166_376_2 = (realValue_0_376 - _zz_when_ArraySlice_l166_376_3);
  assign _zz_when_ArraySlice_l166_376_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_376_4);
  assign _zz_when_ArraySlice_l166_376_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_376_4 = {4'd0, _zz_when_ArraySlice_l166_376_5};
  assign _zz_when_ArraySlice_l166_376_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_377 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_377_1);
  assign _zz_when_ArraySlice_l158_377_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_377_1 = {3'd0, _zz_when_ArraySlice_l158_377_2};
  assign _zz_when_ArraySlice_l158_377_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_377_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_377 = {1'd0, _zz_when_ArraySlice_l159_377_1};
  assign _zz_when_ArraySlice_l159_377_2 = (_zz_when_ArraySlice_l159_377_3 - _zz_when_ArraySlice_l159_377_4);
  assign _zz_when_ArraySlice_l159_377_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_377_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_377_5);
  assign _zz_when_ArraySlice_l159_377_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_377_5 = {3'd0, _zz_when_ArraySlice_l159_377_6};
  assign _zz__zz_realValue_0_377 = {1'd0, wReg};
  assign _zz__zz_realValue_0_377_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_377_1 = (_zz_realValue_0_377_2 + _zz_realValue_0_377_3);
  assign _zz_realValue_0_377_2 = {1'd0, wReg};
  assign _zz_realValue_0_377_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_377_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_377 = {1'd0, _zz_when_ArraySlice_l166_377_1};
  assign _zz_when_ArraySlice_l166_377_2 = (_zz_when_ArraySlice_l166_377_3 + _zz_when_ArraySlice_l166_377_7);
  assign _zz_when_ArraySlice_l166_377_3 = (realValue_0_377 - _zz_when_ArraySlice_l166_377_4);
  assign _zz_when_ArraySlice_l166_377_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_377_5);
  assign _zz_when_ArraySlice_l166_377_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_377_5 = {3'd0, _zz_when_ArraySlice_l166_377_6};
  assign _zz_when_ArraySlice_l166_377_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_378 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_378_1);
  assign _zz_when_ArraySlice_l158_378_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_378_1 = {2'd0, _zz_when_ArraySlice_l158_378_2};
  assign _zz_when_ArraySlice_l158_378_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_378_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_378 = {1'd0, _zz_when_ArraySlice_l159_378_1};
  assign _zz_when_ArraySlice_l159_378_2 = (_zz_when_ArraySlice_l159_378_3 - _zz_when_ArraySlice_l159_378_4);
  assign _zz_when_ArraySlice_l159_378_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_378_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_378_5);
  assign _zz_when_ArraySlice_l159_378_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_378_5 = {2'd0, _zz_when_ArraySlice_l159_378_6};
  assign _zz__zz_realValue_0_378 = {1'd0, wReg};
  assign _zz__zz_realValue_0_378_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_378_1 = (_zz_realValue_0_378_2 + _zz_realValue_0_378_3);
  assign _zz_realValue_0_378_2 = {1'd0, wReg};
  assign _zz_realValue_0_378_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_378_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_378 = {1'd0, _zz_when_ArraySlice_l166_378_1};
  assign _zz_when_ArraySlice_l166_378_2 = (_zz_when_ArraySlice_l166_378_3 + _zz_when_ArraySlice_l166_378_7);
  assign _zz_when_ArraySlice_l166_378_3 = (realValue_0_378 - _zz_when_ArraySlice_l166_378_4);
  assign _zz_when_ArraySlice_l166_378_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_378_5);
  assign _zz_when_ArraySlice_l166_378_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_378_5 = {2'd0, _zz_when_ArraySlice_l166_378_6};
  assign _zz_when_ArraySlice_l166_378_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_379 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_379_1);
  assign _zz_when_ArraySlice_l158_379_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_379_1 = {2'd0, _zz_when_ArraySlice_l158_379_2};
  assign _zz_when_ArraySlice_l158_379_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_379_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_379 = {1'd0, _zz_when_ArraySlice_l159_379_1};
  assign _zz_when_ArraySlice_l159_379_2 = (_zz_when_ArraySlice_l159_379_3 - _zz_when_ArraySlice_l159_379_4);
  assign _zz_when_ArraySlice_l159_379_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_379_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_379_5);
  assign _zz_when_ArraySlice_l159_379_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_379_5 = {2'd0, _zz_when_ArraySlice_l159_379_6};
  assign _zz__zz_realValue_0_379 = {1'd0, wReg};
  assign _zz__zz_realValue_0_379_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_379_1 = (_zz_realValue_0_379_2 + _zz_realValue_0_379_3);
  assign _zz_realValue_0_379_2 = {1'd0, wReg};
  assign _zz_realValue_0_379_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_379_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_379 = {1'd0, _zz_when_ArraySlice_l166_379_1};
  assign _zz_when_ArraySlice_l166_379_2 = (_zz_when_ArraySlice_l166_379_3 + _zz_when_ArraySlice_l166_379_7);
  assign _zz_when_ArraySlice_l166_379_3 = (realValue_0_379 - _zz_when_ArraySlice_l166_379_4);
  assign _zz_when_ArraySlice_l166_379_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_379_5);
  assign _zz_when_ArraySlice_l166_379_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_379_5 = {2'd0, _zz_when_ArraySlice_l166_379_6};
  assign _zz_when_ArraySlice_l166_379_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_380 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_380_1);
  assign _zz_when_ArraySlice_l158_380_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_380_1 = {1'd0, _zz_when_ArraySlice_l158_380_2};
  assign _zz_when_ArraySlice_l158_380_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_380_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_380 = {1'd0, _zz_when_ArraySlice_l159_380_1};
  assign _zz_when_ArraySlice_l159_380_2 = (_zz_when_ArraySlice_l159_380_3 - _zz_when_ArraySlice_l159_380_4);
  assign _zz_when_ArraySlice_l159_380_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_380_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_380_5);
  assign _zz_when_ArraySlice_l159_380_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_380_5 = {1'd0, _zz_when_ArraySlice_l159_380_6};
  assign _zz__zz_realValue_0_380 = {1'd0, wReg};
  assign _zz__zz_realValue_0_380_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_380_1 = (_zz_realValue_0_380_2 + _zz_realValue_0_380_3);
  assign _zz_realValue_0_380_2 = {1'd0, wReg};
  assign _zz_realValue_0_380_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_380_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_380 = {1'd0, _zz_when_ArraySlice_l166_380_1};
  assign _zz_when_ArraySlice_l166_380_2 = (_zz_when_ArraySlice_l166_380_3 + _zz_when_ArraySlice_l166_380_7);
  assign _zz_when_ArraySlice_l166_380_3 = (realValue_0_380 - _zz_when_ArraySlice_l166_380_4);
  assign _zz_when_ArraySlice_l166_380_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_380_5);
  assign _zz_when_ArraySlice_l166_380_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_380_5 = {1'd0, _zz_when_ArraySlice_l166_380_6};
  assign _zz_when_ArraySlice_l166_380_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_381 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_381_1);
  assign _zz_when_ArraySlice_l158_381_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_381_1 = {1'd0, _zz_when_ArraySlice_l158_381_2};
  assign _zz_when_ArraySlice_l158_381_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_381_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_381 = {2'd0, _zz_when_ArraySlice_l159_381_1};
  assign _zz_when_ArraySlice_l159_381_2 = (_zz_when_ArraySlice_l159_381_3 - _zz_when_ArraySlice_l159_381_4);
  assign _zz_when_ArraySlice_l159_381_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_381_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_381_5);
  assign _zz_when_ArraySlice_l159_381_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_381_5 = {1'd0, _zz_when_ArraySlice_l159_381_6};
  assign _zz__zz_realValue_0_381 = {1'd0, wReg};
  assign _zz__zz_realValue_0_381_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_381_1 = (_zz_realValue_0_381_2 + _zz_realValue_0_381_3);
  assign _zz_realValue_0_381_2 = {1'd0, wReg};
  assign _zz_realValue_0_381_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_381_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_381 = {2'd0, _zz_when_ArraySlice_l166_381_1};
  assign _zz_when_ArraySlice_l166_381_2 = (_zz_when_ArraySlice_l166_381_3 + _zz_when_ArraySlice_l166_381_7);
  assign _zz_when_ArraySlice_l166_381_3 = (realValue_0_381 - _zz_when_ArraySlice_l166_381_4);
  assign _zz_when_ArraySlice_l166_381_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_381_5);
  assign _zz_when_ArraySlice_l166_381_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_381_5 = {1'd0, _zz_when_ArraySlice_l166_381_6};
  assign _zz_when_ArraySlice_l166_381_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_382 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_382_1);
  assign _zz_when_ArraySlice_l158_382_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_382_1 = {1'd0, _zz_when_ArraySlice_l158_382_2};
  assign _zz_when_ArraySlice_l158_382_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_382_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_382 = {2'd0, _zz_when_ArraySlice_l159_382_1};
  assign _zz_when_ArraySlice_l159_382_2 = (_zz_when_ArraySlice_l159_382_3 - _zz_when_ArraySlice_l159_382_4);
  assign _zz_when_ArraySlice_l159_382_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_382_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_382_5);
  assign _zz_when_ArraySlice_l159_382_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_382_5 = {1'd0, _zz_when_ArraySlice_l159_382_6};
  assign _zz__zz_realValue_0_382 = {1'd0, wReg};
  assign _zz__zz_realValue_0_382_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_382_1 = (_zz_realValue_0_382_2 + _zz_realValue_0_382_3);
  assign _zz_realValue_0_382_2 = {1'd0, wReg};
  assign _zz_realValue_0_382_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_382_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_382 = {2'd0, _zz_when_ArraySlice_l166_382_1};
  assign _zz_when_ArraySlice_l166_382_2 = (_zz_when_ArraySlice_l166_382_3 + _zz_when_ArraySlice_l166_382_7);
  assign _zz_when_ArraySlice_l166_382_3 = (realValue_0_382 - _zz_when_ArraySlice_l166_382_4);
  assign _zz_when_ArraySlice_l166_382_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_382_5);
  assign _zz_when_ArraySlice_l166_382_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_382_5 = {1'd0, _zz_when_ArraySlice_l166_382_6};
  assign _zz_when_ArraySlice_l166_382_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_383 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_383_1);
  assign _zz_when_ArraySlice_l158_383_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_383_1 = {1'd0, _zz_when_ArraySlice_l158_383_2};
  assign _zz_when_ArraySlice_l158_383_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_383_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_383 = {3'd0, _zz_when_ArraySlice_l159_383_1};
  assign _zz_when_ArraySlice_l159_383_2 = (_zz_when_ArraySlice_l159_383_3 - _zz_when_ArraySlice_l159_383_4);
  assign _zz_when_ArraySlice_l159_383_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_383_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_383_5);
  assign _zz_when_ArraySlice_l159_383_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_383_5 = {1'd0, _zz_when_ArraySlice_l159_383_6};
  assign _zz__zz_realValue_0_383 = {1'd0, wReg};
  assign _zz__zz_realValue_0_383_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_383_1 = (_zz_realValue_0_383_2 + _zz_realValue_0_383_3);
  assign _zz_realValue_0_383_2 = {1'd0, wReg};
  assign _zz_realValue_0_383_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_383_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_383 = {3'd0, _zz_when_ArraySlice_l166_383_1};
  assign _zz_when_ArraySlice_l166_383_2 = (_zz_when_ArraySlice_l166_383_3 + _zz_when_ArraySlice_l166_383_7);
  assign _zz_when_ArraySlice_l166_383_3 = (realValue_0_383 - _zz_when_ArraySlice_l166_383_4);
  assign _zz_when_ArraySlice_l166_383_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_383_5);
  assign _zz_when_ArraySlice_l166_383_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_383_5 = {1'd0, _zz_when_ArraySlice_l166_383_6};
  assign _zz_when_ArraySlice_l166_383_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l260_7_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l260_7_2 = (_zz_when_ArraySlice_l260_7_3 + _zz_when_ArraySlice_l260_7_7);
  assign _zz_when_ArraySlice_l260_7_3 = (_zz_when_ArraySlice_l260_7_4 + 8'h01);
  assign _zz_when_ArraySlice_l260_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l260_7_5);
  assign _zz_when_ArraySlice_l260_7_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l260_7_5 = {1'd0, _zz_when_ArraySlice_l260_7_6};
  assign _zz_when_ArraySlice_l260_7_8 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l260_7_7 = {1'd0, _zz_when_ArraySlice_l260_7_8};
  assign _zz_when_ArraySlice_l263_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l263_7_1 = (_zz_when_ArraySlice_l263_7_2 + 8'h01);
  assign _zz_when_ArraySlice_l263_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l263_7_3);
  assign _zz_when_ArraySlice_l263_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l263_7_3 = {1'd0, _zz_when_ArraySlice_l263_7_4};
  assign _zz_selectReadFifo_7_22 = (selectReadFifo_7 + _zz_selectReadFifo_7_23);
  assign _zz_selectReadFifo_7_24 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_23 = {1'd0, _zz_selectReadFifo_7_24};
  assign _zz_when_ArraySlice_l270_7 = (_zz_when_ArraySlice_l270_7_1 % aReg);
  assign _zz_when_ArraySlice_l270_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l274_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l274_7_3);
  assign _zz_when_ArraySlice_l274_7_1 = _zz_when_ArraySlice_l274_7_2[6:0];
  assign _zz_when_ArraySlice_l274_7_4 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l274_7_3 = {1'd0, _zz_when_ArraySlice_l274_7_4};
  assign _zz_when_ArraySlice_l275_7_1 = (_zz_when_ArraySlice_l275_7_2 - _zz_when_ArraySlice_l275_7_3);
  assign _zz_when_ArraySlice_l275_7 = {5'd0, _zz_when_ArraySlice_l275_7_1};
  assign _zz_when_ArraySlice_l275_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l275_7_4 = 1'b1;
  assign _zz_when_ArraySlice_l275_7_3 = {7'd0, _zz_when_ArraySlice_l275_7_4};
  assign _zz__zz_realValue1_0_46 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_46_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_46_1 = (_zz_realValue1_0_46_2 + _zz_realValue1_0_46_3);
  assign _zz_realValue1_0_46_2 = {1'd0, hReg};
  assign _zz_realValue1_0_46_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l277_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l277_7 = {1'd0, _zz_when_ArraySlice_l277_7_1};
  assign _zz_when_ArraySlice_l277_7_2 = (realValue1_0_46 / aReg);
  assign _zz_selectReadFifo_7_25 = (selectReadFifo_7 - _zz_selectReadFifo_7_26);
  assign _zz_selectReadFifo_7_26 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_384 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_384_1);
  assign _zz_when_ArraySlice_l158_384_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_384_1 = {4'd0, _zz_when_ArraySlice_l158_384_2};
  assign _zz_when_ArraySlice_l158_384_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_384 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_384_1 = (_zz_when_ArraySlice_l159_384_2 - _zz_when_ArraySlice_l159_384_3);
  assign _zz_when_ArraySlice_l159_384_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_384_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_384_4);
  assign _zz_when_ArraySlice_l159_384_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_384_4 = {4'd0, _zz_when_ArraySlice_l159_384_5};
  assign _zz__zz_realValue_0_384 = {1'd0, wReg};
  assign _zz__zz_realValue_0_384_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_384_1 = (_zz_realValue_0_384_2 + _zz_realValue_0_384_3);
  assign _zz_realValue_0_384_2 = {1'd0, wReg};
  assign _zz_realValue_0_384_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_384 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_384_1 = (_zz_when_ArraySlice_l166_384_2 + _zz_when_ArraySlice_l166_384_6);
  assign _zz_when_ArraySlice_l166_384_2 = (realValue_0_384 - _zz_when_ArraySlice_l166_384_3);
  assign _zz_when_ArraySlice_l166_384_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_384_4);
  assign _zz_when_ArraySlice_l166_384_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_384_4 = {4'd0, _zz_when_ArraySlice_l166_384_5};
  assign _zz_when_ArraySlice_l166_384_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_385 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_385_1);
  assign _zz_when_ArraySlice_l158_385_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_385_1 = {3'd0, _zz_when_ArraySlice_l158_385_2};
  assign _zz_when_ArraySlice_l158_385_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_385_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_385 = {1'd0, _zz_when_ArraySlice_l159_385_1};
  assign _zz_when_ArraySlice_l159_385_2 = (_zz_when_ArraySlice_l159_385_3 - _zz_when_ArraySlice_l159_385_4);
  assign _zz_when_ArraySlice_l159_385_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_385_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_385_5);
  assign _zz_when_ArraySlice_l159_385_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_385_5 = {3'd0, _zz_when_ArraySlice_l159_385_6};
  assign _zz__zz_realValue_0_385 = {1'd0, wReg};
  assign _zz__zz_realValue_0_385_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_385_1 = (_zz_realValue_0_385_2 + _zz_realValue_0_385_3);
  assign _zz_realValue_0_385_2 = {1'd0, wReg};
  assign _zz_realValue_0_385_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_385_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_385 = {1'd0, _zz_when_ArraySlice_l166_385_1};
  assign _zz_when_ArraySlice_l166_385_2 = (_zz_when_ArraySlice_l166_385_3 + _zz_when_ArraySlice_l166_385_7);
  assign _zz_when_ArraySlice_l166_385_3 = (realValue_0_385 - _zz_when_ArraySlice_l166_385_4);
  assign _zz_when_ArraySlice_l166_385_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_385_5);
  assign _zz_when_ArraySlice_l166_385_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_385_5 = {3'd0, _zz_when_ArraySlice_l166_385_6};
  assign _zz_when_ArraySlice_l166_385_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_386 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_386_1);
  assign _zz_when_ArraySlice_l158_386_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_386_1 = {2'd0, _zz_when_ArraySlice_l158_386_2};
  assign _zz_when_ArraySlice_l158_386_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_386_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_386 = {1'd0, _zz_when_ArraySlice_l159_386_1};
  assign _zz_when_ArraySlice_l159_386_2 = (_zz_when_ArraySlice_l159_386_3 - _zz_when_ArraySlice_l159_386_4);
  assign _zz_when_ArraySlice_l159_386_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_386_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_386_5);
  assign _zz_when_ArraySlice_l159_386_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_386_5 = {2'd0, _zz_when_ArraySlice_l159_386_6};
  assign _zz__zz_realValue_0_386 = {1'd0, wReg};
  assign _zz__zz_realValue_0_386_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_386_1 = (_zz_realValue_0_386_2 + _zz_realValue_0_386_3);
  assign _zz_realValue_0_386_2 = {1'd0, wReg};
  assign _zz_realValue_0_386_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_386_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_386 = {1'd0, _zz_when_ArraySlice_l166_386_1};
  assign _zz_when_ArraySlice_l166_386_2 = (_zz_when_ArraySlice_l166_386_3 + _zz_when_ArraySlice_l166_386_7);
  assign _zz_when_ArraySlice_l166_386_3 = (realValue_0_386 - _zz_when_ArraySlice_l166_386_4);
  assign _zz_when_ArraySlice_l166_386_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_386_5);
  assign _zz_when_ArraySlice_l166_386_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_386_5 = {2'd0, _zz_when_ArraySlice_l166_386_6};
  assign _zz_when_ArraySlice_l166_386_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_387 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_387_1);
  assign _zz_when_ArraySlice_l158_387_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_387_1 = {2'd0, _zz_when_ArraySlice_l158_387_2};
  assign _zz_when_ArraySlice_l158_387_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_387_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_387 = {1'd0, _zz_when_ArraySlice_l159_387_1};
  assign _zz_when_ArraySlice_l159_387_2 = (_zz_when_ArraySlice_l159_387_3 - _zz_when_ArraySlice_l159_387_4);
  assign _zz_when_ArraySlice_l159_387_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_387_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_387_5);
  assign _zz_when_ArraySlice_l159_387_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_387_5 = {2'd0, _zz_when_ArraySlice_l159_387_6};
  assign _zz__zz_realValue_0_387 = {1'd0, wReg};
  assign _zz__zz_realValue_0_387_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_387_1 = (_zz_realValue_0_387_2 + _zz_realValue_0_387_3);
  assign _zz_realValue_0_387_2 = {1'd0, wReg};
  assign _zz_realValue_0_387_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_387_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_387 = {1'd0, _zz_when_ArraySlice_l166_387_1};
  assign _zz_when_ArraySlice_l166_387_2 = (_zz_when_ArraySlice_l166_387_3 + _zz_when_ArraySlice_l166_387_7);
  assign _zz_when_ArraySlice_l166_387_3 = (realValue_0_387 - _zz_when_ArraySlice_l166_387_4);
  assign _zz_when_ArraySlice_l166_387_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_387_5);
  assign _zz_when_ArraySlice_l166_387_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_387_5 = {2'd0, _zz_when_ArraySlice_l166_387_6};
  assign _zz_when_ArraySlice_l166_387_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_388 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_388_1);
  assign _zz_when_ArraySlice_l158_388_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_388_1 = {1'd0, _zz_when_ArraySlice_l158_388_2};
  assign _zz_when_ArraySlice_l158_388_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_388_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_388 = {1'd0, _zz_when_ArraySlice_l159_388_1};
  assign _zz_when_ArraySlice_l159_388_2 = (_zz_when_ArraySlice_l159_388_3 - _zz_when_ArraySlice_l159_388_4);
  assign _zz_when_ArraySlice_l159_388_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_388_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_388_5);
  assign _zz_when_ArraySlice_l159_388_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_388_5 = {1'd0, _zz_when_ArraySlice_l159_388_6};
  assign _zz__zz_realValue_0_388 = {1'd0, wReg};
  assign _zz__zz_realValue_0_388_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_388_1 = (_zz_realValue_0_388_2 + _zz_realValue_0_388_3);
  assign _zz_realValue_0_388_2 = {1'd0, wReg};
  assign _zz_realValue_0_388_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_388_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_388 = {1'd0, _zz_when_ArraySlice_l166_388_1};
  assign _zz_when_ArraySlice_l166_388_2 = (_zz_when_ArraySlice_l166_388_3 + _zz_when_ArraySlice_l166_388_7);
  assign _zz_when_ArraySlice_l166_388_3 = (realValue_0_388 - _zz_when_ArraySlice_l166_388_4);
  assign _zz_when_ArraySlice_l166_388_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_388_5);
  assign _zz_when_ArraySlice_l166_388_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_388_5 = {1'd0, _zz_when_ArraySlice_l166_388_6};
  assign _zz_when_ArraySlice_l166_388_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_389 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_389_1);
  assign _zz_when_ArraySlice_l158_389_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_389_1 = {1'd0, _zz_when_ArraySlice_l158_389_2};
  assign _zz_when_ArraySlice_l158_389_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_389_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_389 = {2'd0, _zz_when_ArraySlice_l159_389_1};
  assign _zz_when_ArraySlice_l159_389_2 = (_zz_when_ArraySlice_l159_389_3 - _zz_when_ArraySlice_l159_389_4);
  assign _zz_when_ArraySlice_l159_389_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_389_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_389_5);
  assign _zz_when_ArraySlice_l159_389_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_389_5 = {1'd0, _zz_when_ArraySlice_l159_389_6};
  assign _zz__zz_realValue_0_389 = {1'd0, wReg};
  assign _zz__zz_realValue_0_389_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_389_1 = (_zz_realValue_0_389_2 + _zz_realValue_0_389_3);
  assign _zz_realValue_0_389_2 = {1'd0, wReg};
  assign _zz_realValue_0_389_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_389_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_389 = {2'd0, _zz_when_ArraySlice_l166_389_1};
  assign _zz_when_ArraySlice_l166_389_2 = (_zz_when_ArraySlice_l166_389_3 + _zz_when_ArraySlice_l166_389_7);
  assign _zz_when_ArraySlice_l166_389_3 = (realValue_0_389 - _zz_when_ArraySlice_l166_389_4);
  assign _zz_when_ArraySlice_l166_389_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_389_5);
  assign _zz_when_ArraySlice_l166_389_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_389_5 = {1'd0, _zz_when_ArraySlice_l166_389_6};
  assign _zz_when_ArraySlice_l166_389_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_390 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_390_1);
  assign _zz_when_ArraySlice_l158_390_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_390_1 = {1'd0, _zz_when_ArraySlice_l158_390_2};
  assign _zz_when_ArraySlice_l158_390_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_390_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_390 = {2'd0, _zz_when_ArraySlice_l159_390_1};
  assign _zz_when_ArraySlice_l159_390_2 = (_zz_when_ArraySlice_l159_390_3 - _zz_when_ArraySlice_l159_390_4);
  assign _zz_when_ArraySlice_l159_390_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_390_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_390_5);
  assign _zz_when_ArraySlice_l159_390_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_390_5 = {1'd0, _zz_when_ArraySlice_l159_390_6};
  assign _zz__zz_realValue_0_390 = {1'd0, wReg};
  assign _zz__zz_realValue_0_390_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_390_1 = (_zz_realValue_0_390_2 + _zz_realValue_0_390_3);
  assign _zz_realValue_0_390_2 = {1'd0, wReg};
  assign _zz_realValue_0_390_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_390_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_390 = {2'd0, _zz_when_ArraySlice_l166_390_1};
  assign _zz_when_ArraySlice_l166_390_2 = (_zz_when_ArraySlice_l166_390_3 + _zz_when_ArraySlice_l166_390_7);
  assign _zz_when_ArraySlice_l166_390_3 = (realValue_0_390 - _zz_when_ArraySlice_l166_390_4);
  assign _zz_when_ArraySlice_l166_390_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_390_5);
  assign _zz_when_ArraySlice_l166_390_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_390_5 = {1'd0, _zz_when_ArraySlice_l166_390_6};
  assign _zz_when_ArraySlice_l166_390_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_391 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_391_1);
  assign _zz_when_ArraySlice_l158_391_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_391_1 = {1'd0, _zz_when_ArraySlice_l158_391_2};
  assign _zz_when_ArraySlice_l158_391_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_391_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_391 = {3'd0, _zz_when_ArraySlice_l159_391_1};
  assign _zz_when_ArraySlice_l159_391_2 = (_zz_when_ArraySlice_l159_391_3 - _zz_when_ArraySlice_l159_391_4);
  assign _zz_when_ArraySlice_l159_391_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_391_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_391_5);
  assign _zz_when_ArraySlice_l159_391_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_391_5 = {1'd0, _zz_when_ArraySlice_l159_391_6};
  assign _zz__zz_realValue_0_391 = {1'd0, wReg};
  assign _zz__zz_realValue_0_391_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_391_1 = (_zz_realValue_0_391_2 + _zz_realValue_0_391_3);
  assign _zz_realValue_0_391_2 = {1'd0, wReg};
  assign _zz_realValue_0_391_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_391_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_391 = {3'd0, _zz_when_ArraySlice_l166_391_1};
  assign _zz_when_ArraySlice_l166_391_2 = (_zz_when_ArraySlice_l166_391_3 + _zz_when_ArraySlice_l166_391_7);
  assign _zz_when_ArraySlice_l166_391_3 = (realValue_0_391 - _zz_when_ArraySlice_l166_391_4);
  assign _zz_when_ArraySlice_l166_391_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_391_5);
  assign _zz_when_ArraySlice_l166_391_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_391_5 = {1'd0, _zz_when_ArraySlice_l166_391_6};
  assign _zz_when_ArraySlice_l166_391_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l285_7_1 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l285_7_2 = (_zz_when_ArraySlice_l285_7_3 + _zz_when_ArraySlice_l285_7_7);
  assign _zz_when_ArraySlice_l285_7_3 = (_zz_when_ArraySlice_l285_7_4 + 8'h01);
  assign _zz_when_ArraySlice_l285_7_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l285_7_5);
  assign _zz_when_ArraySlice_l285_7_6 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l285_7_5 = {1'd0, _zz_when_ArraySlice_l285_7_6};
  assign _zz_when_ArraySlice_l285_7_8 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l285_7_7 = {1'd0, _zz_when_ArraySlice_l285_7_8};
  assign _zz_when_ArraySlice_l288_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l288_7_1 = (_zz_when_ArraySlice_l288_7_2 + 8'h01);
  assign _zz_when_ArraySlice_l288_7_2 = (selectReadFifo_7 + _zz_when_ArraySlice_l288_7_3);
  assign _zz_when_ArraySlice_l288_7_4 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l288_7_3 = {1'd0, _zz_when_ArraySlice_l288_7_4};
  assign _zz_selectReadFifo_7_27 = (selectReadFifo_7 + _zz_selectReadFifo_7_28);
  assign _zz_selectReadFifo_7_29 = (3'b111 * bReg);
  assign _zz_selectReadFifo_7_28 = {1'd0, _zz_selectReadFifo_7_29};
  assign _zz_when_ArraySlice_l295_7 = (_zz_when_ArraySlice_l295_7_1 % aReg);
  assign _zz_when_ArraySlice_l295_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l306_7_1 = (_zz_when_ArraySlice_l306_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l306_7 = {5'd0, _zz_when_ArraySlice_l306_7_1};
  assign _zz_when_ArraySlice_l306_7_2 = (bReg * aReg);
  assign _zz__zz_realValue1_0_47 = {1'd0, hReg};
  assign _zz__zz_realValue1_0_47_1 = (aReg * 4'b1000);
  assign _zz_realValue1_0_47_1 = (_zz_realValue1_0_47_2 + _zz_realValue1_0_47_3);
  assign _zz_realValue1_0_47_2 = {1'd0, hReg};
  assign _zz_realValue1_0_47_3 = (aReg * 4'b1000);
  assign _zz_when_ArraySlice_l307_7_1 = (outSliceNumb_7_value + 7'h01);
  assign _zz_when_ArraySlice_l307_7 = {1'd0, _zz_when_ArraySlice_l307_7_1};
  assign _zz_when_ArraySlice_l307_7_2 = (realValue1_0_47 / aReg);
  assign _zz_selectReadFifo_7_30 = (selectReadFifo_7 - _zz_selectReadFifo_7_31);
  assign _zz_selectReadFifo_7_31 = {4'd0, bReg};
  assign _zz_when_ArraySlice_l158_392 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_392_1);
  assign _zz_when_ArraySlice_l158_392_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_392_1 = {4'd0, _zz_when_ArraySlice_l158_392_2};
  assign _zz_when_ArraySlice_l158_392_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_392 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_392_1 = (_zz_when_ArraySlice_l159_392_2 - _zz_when_ArraySlice_l159_392_3);
  assign _zz_when_ArraySlice_l159_392_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_392_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_392_4);
  assign _zz_when_ArraySlice_l159_392_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_392_4 = {4'd0, _zz_when_ArraySlice_l159_392_5};
  assign _zz__zz_realValue_0_392 = {1'd0, wReg};
  assign _zz__zz_realValue_0_392_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_392_1 = (_zz_realValue_0_392_2 + _zz_realValue_0_392_3);
  assign _zz_realValue_0_392_2 = {1'd0, wReg};
  assign _zz_realValue_0_392_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_392 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_392_1 = (_zz_when_ArraySlice_l166_392_2 + _zz_when_ArraySlice_l166_392_6);
  assign _zz_when_ArraySlice_l166_392_2 = (realValue_0_392 - _zz_when_ArraySlice_l166_392_3);
  assign _zz_when_ArraySlice_l166_392_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_392_4);
  assign _zz_when_ArraySlice_l166_392_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_392_4 = {4'd0, _zz_when_ArraySlice_l166_392_5};
  assign _zz_when_ArraySlice_l166_392_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_393 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_393_1);
  assign _zz_when_ArraySlice_l158_393_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_393_1 = {3'd0, _zz_when_ArraySlice_l158_393_2};
  assign _zz_when_ArraySlice_l158_393_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_393_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_393 = {1'd0, _zz_when_ArraySlice_l159_393_1};
  assign _zz_when_ArraySlice_l159_393_2 = (_zz_when_ArraySlice_l159_393_3 - _zz_when_ArraySlice_l159_393_4);
  assign _zz_when_ArraySlice_l159_393_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_393_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_393_5);
  assign _zz_when_ArraySlice_l159_393_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_393_5 = {3'd0, _zz_when_ArraySlice_l159_393_6};
  assign _zz__zz_realValue_0_393 = {1'd0, wReg};
  assign _zz__zz_realValue_0_393_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_393_1 = (_zz_realValue_0_393_2 + _zz_realValue_0_393_3);
  assign _zz_realValue_0_393_2 = {1'd0, wReg};
  assign _zz_realValue_0_393_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_393_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_393 = {1'd0, _zz_when_ArraySlice_l166_393_1};
  assign _zz_when_ArraySlice_l166_393_2 = (_zz_when_ArraySlice_l166_393_3 + _zz_when_ArraySlice_l166_393_7);
  assign _zz_when_ArraySlice_l166_393_3 = (realValue_0_393 - _zz_when_ArraySlice_l166_393_4);
  assign _zz_when_ArraySlice_l166_393_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_393_5);
  assign _zz_when_ArraySlice_l166_393_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_393_5 = {3'd0, _zz_when_ArraySlice_l166_393_6};
  assign _zz_when_ArraySlice_l166_393_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_394 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_394_1);
  assign _zz_when_ArraySlice_l158_394_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_394_1 = {2'd0, _zz_when_ArraySlice_l158_394_2};
  assign _zz_when_ArraySlice_l158_394_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_394_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_394 = {1'd0, _zz_when_ArraySlice_l159_394_1};
  assign _zz_when_ArraySlice_l159_394_2 = (_zz_when_ArraySlice_l159_394_3 - _zz_when_ArraySlice_l159_394_4);
  assign _zz_when_ArraySlice_l159_394_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_394_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_394_5);
  assign _zz_when_ArraySlice_l159_394_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_394_5 = {2'd0, _zz_when_ArraySlice_l159_394_6};
  assign _zz__zz_realValue_0_394 = {1'd0, wReg};
  assign _zz__zz_realValue_0_394_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_394_1 = (_zz_realValue_0_394_2 + _zz_realValue_0_394_3);
  assign _zz_realValue_0_394_2 = {1'd0, wReg};
  assign _zz_realValue_0_394_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_394_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_394 = {1'd0, _zz_when_ArraySlice_l166_394_1};
  assign _zz_when_ArraySlice_l166_394_2 = (_zz_when_ArraySlice_l166_394_3 + _zz_when_ArraySlice_l166_394_7);
  assign _zz_when_ArraySlice_l166_394_3 = (realValue_0_394 - _zz_when_ArraySlice_l166_394_4);
  assign _zz_when_ArraySlice_l166_394_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_394_5);
  assign _zz_when_ArraySlice_l166_394_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_394_5 = {2'd0, _zz_when_ArraySlice_l166_394_6};
  assign _zz_when_ArraySlice_l166_394_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_395 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_395_1);
  assign _zz_when_ArraySlice_l158_395_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_395_1 = {2'd0, _zz_when_ArraySlice_l158_395_2};
  assign _zz_when_ArraySlice_l158_395_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_395_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_395 = {1'd0, _zz_when_ArraySlice_l159_395_1};
  assign _zz_when_ArraySlice_l159_395_2 = (_zz_when_ArraySlice_l159_395_3 - _zz_when_ArraySlice_l159_395_4);
  assign _zz_when_ArraySlice_l159_395_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_395_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_395_5);
  assign _zz_when_ArraySlice_l159_395_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_395_5 = {2'd0, _zz_when_ArraySlice_l159_395_6};
  assign _zz__zz_realValue_0_395 = {1'd0, wReg};
  assign _zz__zz_realValue_0_395_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_395_1 = (_zz_realValue_0_395_2 + _zz_realValue_0_395_3);
  assign _zz_realValue_0_395_2 = {1'd0, wReg};
  assign _zz_realValue_0_395_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_395_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_395 = {1'd0, _zz_when_ArraySlice_l166_395_1};
  assign _zz_when_ArraySlice_l166_395_2 = (_zz_when_ArraySlice_l166_395_3 + _zz_when_ArraySlice_l166_395_7);
  assign _zz_when_ArraySlice_l166_395_3 = (realValue_0_395 - _zz_when_ArraySlice_l166_395_4);
  assign _zz_when_ArraySlice_l166_395_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_395_5);
  assign _zz_when_ArraySlice_l166_395_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_395_5 = {2'd0, _zz_when_ArraySlice_l166_395_6};
  assign _zz_when_ArraySlice_l166_395_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_396 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_396_1);
  assign _zz_when_ArraySlice_l158_396_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_396_1 = {1'd0, _zz_when_ArraySlice_l158_396_2};
  assign _zz_when_ArraySlice_l158_396_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_396_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_396 = {1'd0, _zz_when_ArraySlice_l159_396_1};
  assign _zz_when_ArraySlice_l159_396_2 = (_zz_when_ArraySlice_l159_396_3 - _zz_when_ArraySlice_l159_396_4);
  assign _zz_when_ArraySlice_l159_396_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_396_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_396_5);
  assign _zz_when_ArraySlice_l159_396_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_396_5 = {1'd0, _zz_when_ArraySlice_l159_396_6};
  assign _zz__zz_realValue_0_396 = {1'd0, wReg};
  assign _zz__zz_realValue_0_396_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_396_1 = (_zz_realValue_0_396_2 + _zz_realValue_0_396_3);
  assign _zz_realValue_0_396_2 = {1'd0, wReg};
  assign _zz_realValue_0_396_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_396_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_396 = {1'd0, _zz_when_ArraySlice_l166_396_1};
  assign _zz_when_ArraySlice_l166_396_2 = (_zz_when_ArraySlice_l166_396_3 + _zz_when_ArraySlice_l166_396_7);
  assign _zz_when_ArraySlice_l166_396_3 = (realValue_0_396 - _zz_when_ArraySlice_l166_396_4);
  assign _zz_when_ArraySlice_l166_396_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_396_5);
  assign _zz_when_ArraySlice_l166_396_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_396_5 = {1'd0, _zz_when_ArraySlice_l166_396_6};
  assign _zz_when_ArraySlice_l166_396_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_397 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_397_1);
  assign _zz_when_ArraySlice_l158_397_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_397_1 = {1'd0, _zz_when_ArraySlice_l158_397_2};
  assign _zz_when_ArraySlice_l158_397_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_397_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_397 = {2'd0, _zz_when_ArraySlice_l159_397_1};
  assign _zz_when_ArraySlice_l159_397_2 = (_zz_when_ArraySlice_l159_397_3 - _zz_when_ArraySlice_l159_397_4);
  assign _zz_when_ArraySlice_l159_397_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_397_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_397_5);
  assign _zz_when_ArraySlice_l159_397_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_397_5 = {1'd0, _zz_when_ArraySlice_l159_397_6};
  assign _zz__zz_realValue_0_397 = {1'd0, wReg};
  assign _zz__zz_realValue_0_397_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_397_1 = (_zz_realValue_0_397_2 + _zz_realValue_0_397_3);
  assign _zz_realValue_0_397_2 = {1'd0, wReg};
  assign _zz_realValue_0_397_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_397_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_397 = {2'd0, _zz_when_ArraySlice_l166_397_1};
  assign _zz_when_ArraySlice_l166_397_2 = (_zz_when_ArraySlice_l166_397_3 + _zz_when_ArraySlice_l166_397_7);
  assign _zz_when_ArraySlice_l166_397_3 = (realValue_0_397 - _zz_when_ArraySlice_l166_397_4);
  assign _zz_when_ArraySlice_l166_397_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_397_5);
  assign _zz_when_ArraySlice_l166_397_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_397_5 = {1'd0, _zz_when_ArraySlice_l166_397_6};
  assign _zz_when_ArraySlice_l166_397_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_398 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_398_1);
  assign _zz_when_ArraySlice_l158_398_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_398_1 = {1'd0, _zz_when_ArraySlice_l158_398_2};
  assign _zz_when_ArraySlice_l158_398_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_398_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_398 = {2'd0, _zz_when_ArraySlice_l159_398_1};
  assign _zz_when_ArraySlice_l159_398_2 = (_zz_when_ArraySlice_l159_398_3 - _zz_when_ArraySlice_l159_398_4);
  assign _zz_when_ArraySlice_l159_398_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_398_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_398_5);
  assign _zz_when_ArraySlice_l159_398_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_398_5 = {1'd0, _zz_when_ArraySlice_l159_398_6};
  assign _zz__zz_realValue_0_398 = {1'd0, wReg};
  assign _zz__zz_realValue_0_398_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_398_1 = (_zz_realValue_0_398_2 + _zz_realValue_0_398_3);
  assign _zz_realValue_0_398_2 = {1'd0, wReg};
  assign _zz_realValue_0_398_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_398_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_398 = {2'd0, _zz_when_ArraySlice_l166_398_1};
  assign _zz_when_ArraySlice_l166_398_2 = (_zz_when_ArraySlice_l166_398_3 + _zz_when_ArraySlice_l166_398_7);
  assign _zz_when_ArraySlice_l166_398_3 = (realValue_0_398 - _zz_when_ArraySlice_l166_398_4);
  assign _zz_when_ArraySlice_l166_398_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_398_5);
  assign _zz_when_ArraySlice_l166_398_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_398_5 = {1'd0, _zz_when_ArraySlice_l166_398_6};
  assign _zz_when_ArraySlice_l166_398_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_399 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_399_1);
  assign _zz_when_ArraySlice_l158_399_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_399_1 = {1'd0, _zz_when_ArraySlice_l158_399_2};
  assign _zz_when_ArraySlice_l158_399_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_399_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_399 = {3'd0, _zz_when_ArraySlice_l159_399_1};
  assign _zz_when_ArraySlice_l159_399_2 = (_zz_when_ArraySlice_l159_399_3 - _zz_when_ArraySlice_l159_399_4);
  assign _zz_when_ArraySlice_l159_399_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_399_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_399_5);
  assign _zz_when_ArraySlice_l159_399_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_399_5 = {1'd0, _zz_when_ArraySlice_l159_399_6};
  assign _zz__zz_realValue_0_399 = {1'd0, wReg};
  assign _zz__zz_realValue_0_399_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_399_1 = (_zz_realValue_0_399_2 + _zz_realValue_0_399_3);
  assign _zz_realValue_0_399_2 = {1'd0, wReg};
  assign _zz_realValue_0_399_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_399_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_399 = {3'd0, _zz_when_ArraySlice_l166_399_1};
  assign _zz_when_ArraySlice_l166_399_2 = (_zz_when_ArraySlice_l166_399_3 + _zz_when_ArraySlice_l166_399_7);
  assign _zz_when_ArraySlice_l166_399_3 = (realValue_0_399 - _zz_when_ArraySlice_l166_399_4);
  assign _zz_when_ArraySlice_l166_399_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_399_5);
  assign _zz_when_ArraySlice_l166_399_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_399_5 = {1'd0, _zz_when_ArraySlice_l166_399_6};
  assign _zz_when_ArraySlice_l166_399_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l318_7 = (_zz_when_ArraySlice_l318_7_1 % aReg);
  assign _zz_when_ArraySlice_l318_7_1 = (handshakeTimes_7_value + 13'h0001);
  assign _zz_when_ArraySlice_l304_7 = {1'd0, wReg};
  assign _zz_when_ArraySlice_l304_7_1 = (selectReadFifo_7 + _zz_when_ArraySlice_l304_7_2);
  assign _zz_when_ArraySlice_l304_7_3 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l304_7_2 = {1'd0, _zz_when_ArraySlice_l304_7_3};
  assign _zz_when_ArraySlice_l325_7_1 = (_zz_when_ArraySlice_l325_7_2 - 8'h01);
  assign _zz_when_ArraySlice_l325_7 = {5'd0, _zz_when_ArraySlice_l325_7_1};
  assign _zz_when_ArraySlice_l325_7_2 = (bReg * aReg);
  assign _zz_when_ArraySlice_l182 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_1 = (selectReadFifo_0 - _zz_when_ArraySlice_l182_2);
  assign _zz_when_ArraySlice_l182_2 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l182_1_1 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_1_2 = (selectReadFifo_1 - _zz_when_ArraySlice_l182_1_3);
  assign _zz_when_ArraySlice_l182_1_3 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l182_2_1 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_2_2 = (selectReadFifo_2 - _zz_when_ArraySlice_l182_2_3);
  assign _zz_when_ArraySlice_l182_2_3 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l182_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_3_1 = (selectReadFifo_3 - _zz_when_ArraySlice_l182_3_2);
  assign _zz_when_ArraySlice_l182_3_2 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l182_4 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_4_1 = (selectReadFifo_4 - _zz_when_ArraySlice_l182_4_2);
  assign _zz_when_ArraySlice_l182_4_2 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l182_5 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_5_1 = (selectReadFifo_5 - _zz_when_ArraySlice_l182_5_2);
  assign _zz_when_ArraySlice_l182_5_2 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l182_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_6_1 = (selectReadFifo_6 - _zz_when_ArraySlice_l182_6_2);
  assign _zz_when_ArraySlice_l182_6_2 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l182_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_7_1 = (selectReadFifo_7 - _zz_when_ArraySlice_l182_7_2);
  assign _zz_when_ArraySlice_l182_7_2 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l341_1 = (hReg - 7'h01);
  assign _zz_when_ArraySlice_l342 = (wReg - 7'h01);
  assign _zz_when_ArraySlice_l158_400 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_400_1);
  assign _zz_when_ArraySlice_l158_400_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_400_1 = {4'd0, _zz_when_ArraySlice_l158_400_2};
  assign _zz_when_ArraySlice_l158_400_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_400 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_400_1 = (_zz_when_ArraySlice_l159_400_2 - _zz_when_ArraySlice_l159_400_3);
  assign _zz_when_ArraySlice_l159_400_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_400_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_400_4);
  assign _zz_when_ArraySlice_l159_400_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_400_4 = {4'd0, _zz_when_ArraySlice_l159_400_5};
  assign _zz__zz_realValue_0_400 = {1'd0, wReg};
  assign _zz__zz_realValue_0_400_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_400_1 = (_zz_realValue_0_400_2 + _zz_realValue_0_400_3);
  assign _zz_realValue_0_400_2 = {1'd0, wReg};
  assign _zz_realValue_0_400_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_400 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_400_1 = (_zz_when_ArraySlice_l166_400_2 + _zz_when_ArraySlice_l166_400_6);
  assign _zz_when_ArraySlice_l166_400_2 = (realValue_0_400 - _zz_when_ArraySlice_l166_400_3);
  assign _zz_when_ArraySlice_l166_400_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_400_4);
  assign _zz_when_ArraySlice_l166_400_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_400_4 = {4'd0, _zz_when_ArraySlice_l166_400_5};
  assign _zz_when_ArraySlice_l166_400_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_401 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_401_1);
  assign _zz_when_ArraySlice_l158_401_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_401_1 = {3'd0, _zz_when_ArraySlice_l158_401_2};
  assign _zz_when_ArraySlice_l158_401_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_401_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_401 = {1'd0, _zz_when_ArraySlice_l159_401_1};
  assign _zz_when_ArraySlice_l159_401_2 = (_zz_when_ArraySlice_l159_401_3 - _zz_when_ArraySlice_l159_401_4);
  assign _zz_when_ArraySlice_l159_401_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_401_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_401_5);
  assign _zz_when_ArraySlice_l159_401_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_401_5 = {3'd0, _zz_when_ArraySlice_l159_401_6};
  assign _zz__zz_realValue_0_401 = {1'd0, wReg};
  assign _zz__zz_realValue_0_401_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_401_1 = (_zz_realValue_0_401_2 + _zz_realValue_0_401_3);
  assign _zz_realValue_0_401_2 = {1'd0, wReg};
  assign _zz_realValue_0_401_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_401_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_401 = {1'd0, _zz_when_ArraySlice_l166_401_1};
  assign _zz_when_ArraySlice_l166_401_2 = (_zz_when_ArraySlice_l166_401_3 + _zz_when_ArraySlice_l166_401_7);
  assign _zz_when_ArraySlice_l166_401_3 = (realValue_0_401 - _zz_when_ArraySlice_l166_401_4);
  assign _zz_when_ArraySlice_l166_401_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_401_5);
  assign _zz_when_ArraySlice_l166_401_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_401_5 = {3'd0, _zz_when_ArraySlice_l166_401_6};
  assign _zz_when_ArraySlice_l166_401_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_402 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_402_1);
  assign _zz_when_ArraySlice_l158_402_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_402_1 = {2'd0, _zz_when_ArraySlice_l158_402_2};
  assign _zz_when_ArraySlice_l158_402_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_402_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_402 = {1'd0, _zz_when_ArraySlice_l159_402_1};
  assign _zz_when_ArraySlice_l159_402_2 = (_zz_when_ArraySlice_l159_402_3 - _zz_when_ArraySlice_l159_402_4);
  assign _zz_when_ArraySlice_l159_402_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_402_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_402_5);
  assign _zz_when_ArraySlice_l159_402_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_402_5 = {2'd0, _zz_when_ArraySlice_l159_402_6};
  assign _zz__zz_realValue_0_402 = {1'd0, wReg};
  assign _zz__zz_realValue_0_402_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_402_1 = (_zz_realValue_0_402_2 + _zz_realValue_0_402_3);
  assign _zz_realValue_0_402_2 = {1'd0, wReg};
  assign _zz_realValue_0_402_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_402_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_402 = {1'd0, _zz_when_ArraySlice_l166_402_1};
  assign _zz_when_ArraySlice_l166_402_2 = (_zz_when_ArraySlice_l166_402_3 + _zz_when_ArraySlice_l166_402_7);
  assign _zz_when_ArraySlice_l166_402_3 = (realValue_0_402 - _zz_when_ArraySlice_l166_402_4);
  assign _zz_when_ArraySlice_l166_402_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_402_5);
  assign _zz_when_ArraySlice_l166_402_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_402_5 = {2'd0, _zz_when_ArraySlice_l166_402_6};
  assign _zz_when_ArraySlice_l166_402_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_403 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_403_1);
  assign _zz_when_ArraySlice_l158_403_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_403_1 = {2'd0, _zz_when_ArraySlice_l158_403_2};
  assign _zz_when_ArraySlice_l158_403_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_403_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_403 = {1'd0, _zz_when_ArraySlice_l159_403_1};
  assign _zz_when_ArraySlice_l159_403_2 = (_zz_when_ArraySlice_l159_403_3 - _zz_when_ArraySlice_l159_403_4);
  assign _zz_when_ArraySlice_l159_403_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_403_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_403_5);
  assign _zz_when_ArraySlice_l159_403_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_403_5 = {2'd0, _zz_when_ArraySlice_l159_403_6};
  assign _zz__zz_realValue_0_403 = {1'd0, wReg};
  assign _zz__zz_realValue_0_403_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_403_1 = (_zz_realValue_0_403_2 + _zz_realValue_0_403_3);
  assign _zz_realValue_0_403_2 = {1'd0, wReg};
  assign _zz_realValue_0_403_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_403_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_403 = {1'd0, _zz_when_ArraySlice_l166_403_1};
  assign _zz_when_ArraySlice_l166_403_2 = (_zz_when_ArraySlice_l166_403_3 + _zz_when_ArraySlice_l166_403_7);
  assign _zz_when_ArraySlice_l166_403_3 = (realValue_0_403 - _zz_when_ArraySlice_l166_403_4);
  assign _zz_when_ArraySlice_l166_403_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_403_5);
  assign _zz_when_ArraySlice_l166_403_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_403_5 = {2'd0, _zz_when_ArraySlice_l166_403_6};
  assign _zz_when_ArraySlice_l166_403_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_404 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_404_1);
  assign _zz_when_ArraySlice_l158_404_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_404_1 = {1'd0, _zz_when_ArraySlice_l158_404_2};
  assign _zz_when_ArraySlice_l158_404_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_404_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_404 = {1'd0, _zz_when_ArraySlice_l159_404_1};
  assign _zz_when_ArraySlice_l159_404_2 = (_zz_when_ArraySlice_l159_404_3 - _zz_when_ArraySlice_l159_404_4);
  assign _zz_when_ArraySlice_l159_404_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_404_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_404_5);
  assign _zz_when_ArraySlice_l159_404_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_404_5 = {1'd0, _zz_when_ArraySlice_l159_404_6};
  assign _zz__zz_realValue_0_404 = {1'd0, wReg};
  assign _zz__zz_realValue_0_404_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_404_1 = (_zz_realValue_0_404_2 + _zz_realValue_0_404_3);
  assign _zz_realValue_0_404_2 = {1'd0, wReg};
  assign _zz_realValue_0_404_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_404_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_404 = {1'd0, _zz_when_ArraySlice_l166_404_1};
  assign _zz_when_ArraySlice_l166_404_2 = (_zz_when_ArraySlice_l166_404_3 + _zz_when_ArraySlice_l166_404_7);
  assign _zz_when_ArraySlice_l166_404_3 = (realValue_0_404 - _zz_when_ArraySlice_l166_404_4);
  assign _zz_when_ArraySlice_l166_404_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_404_5);
  assign _zz_when_ArraySlice_l166_404_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_404_5 = {1'd0, _zz_when_ArraySlice_l166_404_6};
  assign _zz_when_ArraySlice_l166_404_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_405 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_405_1);
  assign _zz_when_ArraySlice_l158_405_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_405_1 = {1'd0, _zz_when_ArraySlice_l158_405_2};
  assign _zz_when_ArraySlice_l158_405_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_405_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_405 = {2'd0, _zz_when_ArraySlice_l159_405_1};
  assign _zz_when_ArraySlice_l159_405_2 = (_zz_when_ArraySlice_l159_405_3 - _zz_when_ArraySlice_l159_405_4);
  assign _zz_when_ArraySlice_l159_405_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_405_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_405_5);
  assign _zz_when_ArraySlice_l159_405_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_405_5 = {1'd0, _zz_when_ArraySlice_l159_405_6};
  assign _zz__zz_realValue_0_405 = {1'd0, wReg};
  assign _zz__zz_realValue_0_405_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_405_1 = (_zz_realValue_0_405_2 + _zz_realValue_0_405_3);
  assign _zz_realValue_0_405_2 = {1'd0, wReg};
  assign _zz_realValue_0_405_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_405_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_405 = {2'd0, _zz_when_ArraySlice_l166_405_1};
  assign _zz_when_ArraySlice_l166_405_2 = (_zz_when_ArraySlice_l166_405_3 + _zz_when_ArraySlice_l166_405_7);
  assign _zz_when_ArraySlice_l166_405_3 = (realValue_0_405 - _zz_when_ArraySlice_l166_405_4);
  assign _zz_when_ArraySlice_l166_405_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_405_5);
  assign _zz_when_ArraySlice_l166_405_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_405_5 = {1'd0, _zz_when_ArraySlice_l166_405_6};
  assign _zz_when_ArraySlice_l166_405_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_406 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_406_1);
  assign _zz_when_ArraySlice_l158_406_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_406_1 = {1'd0, _zz_when_ArraySlice_l158_406_2};
  assign _zz_when_ArraySlice_l158_406_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_406_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_406 = {2'd0, _zz_when_ArraySlice_l159_406_1};
  assign _zz_when_ArraySlice_l159_406_2 = (_zz_when_ArraySlice_l159_406_3 - _zz_when_ArraySlice_l159_406_4);
  assign _zz_when_ArraySlice_l159_406_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_406_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_406_5);
  assign _zz_when_ArraySlice_l159_406_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_406_5 = {1'd0, _zz_when_ArraySlice_l159_406_6};
  assign _zz__zz_realValue_0_406 = {1'd0, wReg};
  assign _zz__zz_realValue_0_406_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_406_1 = (_zz_realValue_0_406_2 + _zz_realValue_0_406_3);
  assign _zz_realValue_0_406_2 = {1'd0, wReg};
  assign _zz_realValue_0_406_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_406_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_406 = {2'd0, _zz_when_ArraySlice_l166_406_1};
  assign _zz_when_ArraySlice_l166_406_2 = (_zz_when_ArraySlice_l166_406_3 + _zz_when_ArraySlice_l166_406_7);
  assign _zz_when_ArraySlice_l166_406_3 = (realValue_0_406 - _zz_when_ArraySlice_l166_406_4);
  assign _zz_when_ArraySlice_l166_406_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_406_5);
  assign _zz_when_ArraySlice_l166_406_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_406_5 = {1'd0, _zz_when_ArraySlice_l166_406_6};
  assign _zz_when_ArraySlice_l166_406_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_407 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_407_1);
  assign _zz_when_ArraySlice_l158_407_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_407_1 = {1'd0, _zz_when_ArraySlice_l158_407_2};
  assign _zz_when_ArraySlice_l158_407_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_407_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_407 = {3'd0, _zz_when_ArraySlice_l159_407_1};
  assign _zz_when_ArraySlice_l159_407_2 = (_zz_when_ArraySlice_l159_407_3 - _zz_when_ArraySlice_l159_407_4);
  assign _zz_when_ArraySlice_l159_407_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_407_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_407_5);
  assign _zz_when_ArraySlice_l159_407_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_407_5 = {1'd0, _zz_when_ArraySlice_l159_407_6};
  assign _zz__zz_realValue_0_407 = {1'd0, wReg};
  assign _zz__zz_realValue_0_407_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_407_1 = (_zz_realValue_0_407_2 + _zz_realValue_0_407_3);
  assign _zz_realValue_0_407_2 = {1'd0, wReg};
  assign _zz_realValue_0_407_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_407_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_407 = {3'd0, _zz_when_ArraySlice_l166_407_1};
  assign _zz_when_ArraySlice_l166_407_2 = (_zz_when_ArraySlice_l166_407_3 + _zz_when_ArraySlice_l166_407_7);
  assign _zz_when_ArraySlice_l166_407_3 = (realValue_0_407 - _zz_when_ArraySlice_l166_407_4);
  assign _zz_when_ArraySlice_l166_407_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_407_5);
  assign _zz_when_ArraySlice_l166_407_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_407_5 = {1'd0, _zz_when_ArraySlice_l166_407_6};
  assign _zz_when_ArraySlice_l166_407_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_408 = (selectReadFifo_0 + _zz_when_ArraySlice_l158_408_1);
  assign _zz_when_ArraySlice_l158_408_2 = 4'b0000;
  assign _zz_when_ArraySlice_l158_408_1 = {4'd0, _zz_when_ArraySlice_l158_408_2};
  assign _zz_when_ArraySlice_l158_408_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_408 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l159_408_1 = (_zz_when_ArraySlice_l159_408_2 - _zz_when_ArraySlice_l159_408_3);
  assign _zz_when_ArraySlice_l159_408_2 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_408_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l159_408_4);
  assign _zz_when_ArraySlice_l159_408_5 = 4'b0000;
  assign _zz_when_ArraySlice_l159_408_4 = {4'd0, _zz_when_ArraySlice_l159_408_5};
  assign _zz__zz_realValue_0_408 = {1'd0, wReg};
  assign _zz__zz_realValue_0_408_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_408_1 = (_zz_realValue_0_408_2 + _zz_realValue_0_408_3);
  assign _zz_realValue_0_408_2 = {1'd0, wReg};
  assign _zz_realValue_0_408_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_408 = (4'b1000 * bReg);
  assign _zz_when_ArraySlice_l166_408_1 = (_zz_when_ArraySlice_l166_408_2 + _zz_when_ArraySlice_l166_408_6);
  assign _zz_when_ArraySlice_l166_408_2 = (realValue_0_408 - _zz_when_ArraySlice_l166_408_3);
  assign _zz_when_ArraySlice_l166_408_3 = (selectReadFifo_0 + _zz_when_ArraySlice_l166_408_4);
  assign _zz_when_ArraySlice_l166_408_5 = 4'b0000;
  assign _zz_when_ArraySlice_l166_408_4 = {4'd0, _zz_when_ArraySlice_l166_408_5};
  assign _zz_when_ArraySlice_l166_408_6 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_409 = (selectReadFifo_1 + _zz_when_ArraySlice_l158_409_1);
  assign _zz_when_ArraySlice_l158_409_2 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l158_409_1 = {3'd0, _zz_when_ArraySlice_l158_409_2};
  assign _zz_when_ArraySlice_l158_409_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_409_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l159_409 = {1'd0, _zz_when_ArraySlice_l159_409_1};
  assign _zz_when_ArraySlice_l159_409_2 = (_zz_when_ArraySlice_l159_409_3 - _zz_when_ArraySlice_l159_409_4);
  assign _zz_when_ArraySlice_l159_409_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_409_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l159_409_5);
  assign _zz_when_ArraySlice_l159_409_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l159_409_5 = {3'd0, _zz_when_ArraySlice_l159_409_6};
  assign _zz__zz_realValue_0_409 = {1'd0, wReg};
  assign _zz__zz_realValue_0_409_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_409_1 = (_zz_realValue_0_409_2 + _zz_realValue_0_409_3);
  assign _zz_realValue_0_409_2 = {1'd0, wReg};
  assign _zz_realValue_0_409_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_409_1 = (3'b111 * bReg);
  assign _zz_when_ArraySlice_l166_409 = {1'd0, _zz_when_ArraySlice_l166_409_1};
  assign _zz_when_ArraySlice_l166_409_2 = (_zz_when_ArraySlice_l166_409_3 + _zz_when_ArraySlice_l166_409_7);
  assign _zz_when_ArraySlice_l166_409_3 = (realValue_0_409 - _zz_when_ArraySlice_l166_409_4);
  assign _zz_when_ArraySlice_l166_409_4 = (selectReadFifo_1 + _zz_when_ArraySlice_l166_409_5);
  assign _zz_when_ArraySlice_l166_409_6 = (bReg * 1'b1);
  assign _zz_when_ArraySlice_l166_409_5 = {3'd0, _zz_when_ArraySlice_l166_409_6};
  assign _zz_when_ArraySlice_l166_409_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_410 = (selectReadFifo_2 + _zz_when_ArraySlice_l158_410_1);
  assign _zz_when_ArraySlice_l158_410_2 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l158_410_1 = {2'd0, _zz_when_ArraySlice_l158_410_2};
  assign _zz_when_ArraySlice_l158_410_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_410_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l159_410 = {1'd0, _zz_when_ArraySlice_l159_410_1};
  assign _zz_when_ArraySlice_l159_410_2 = (_zz_when_ArraySlice_l159_410_3 - _zz_when_ArraySlice_l159_410_4);
  assign _zz_when_ArraySlice_l159_410_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_410_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l159_410_5);
  assign _zz_when_ArraySlice_l159_410_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l159_410_5 = {2'd0, _zz_when_ArraySlice_l159_410_6};
  assign _zz__zz_realValue_0_410 = {1'd0, wReg};
  assign _zz__zz_realValue_0_410_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_410_1 = (_zz_realValue_0_410_2 + _zz_realValue_0_410_3);
  assign _zz_realValue_0_410_2 = {1'd0, wReg};
  assign _zz_realValue_0_410_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_410_1 = (3'b110 * bReg);
  assign _zz_when_ArraySlice_l166_410 = {1'd0, _zz_when_ArraySlice_l166_410_1};
  assign _zz_when_ArraySlice_l166_410_2 = (_zz_when_ArraySlice_l166_410_3 + _zz_when_ArraySlice_l166_410_7);
  assign _zz_when_ArraySlice_l166_410_3 = (realValue_0_410 - _zz_when_ArraySlice_l166_410_4);
  assign _zz_when_ArraySlice_l166_410_4 = (selectReadFifo_2 + _zz_when_ArraySlice_l166_410_5);
  assign _zz_when_ArraySlice_l166_410_6 = (bReg * 2'b10);
  assign _zz_when_ArraySlice_l166_410_5 = {2'd0, _zz_when_ArraySlice_l166_410_6};
  assign _zz_when_ArraySlice_l166_410_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_411 = (selectReadFifo_3 + _zz_when_ArraySlice_l158_411_1);
  assign _zz_when_ArraySlice_l158_411_2 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l158_411_1 = {2'd0, _zz_when_ArraySlice_l158_411_2};
  assign _zz_when_ArraySlice_l158_411_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_411_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l159_411 = {1'd0, _zz_when_ArraySlice_l159_411_1};
  assign _zz_when_ArraySlice_l159_411_2 = (_zz_when_ArraySlice_l159_411_3 - _zz_when_ArraySlice_l159_411_4);
  assign _zz_when_ArraySlice_l159_411_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_411_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l159_411_5);
  assign _zz_when_ArraySlice_l159_411_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l159_411_5 = {2'd0, _zz_when_ArraySlice_l159_411_6};
  assign _zz__zz_realValue_0_411 = {1'd0, wReg};
  assign _zz__zz_realValue_0_411_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_411_1 = (_zz_realValue_0_411_2 + _zz_realValue_0_411_3);
  assign _zz_realValue_0_411_2 = {1'd0, wReg};
  assign _zz_realValue_0_411_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_411_1 = (3'b101 * bReg);
  assign _zz_when_ArraySlice_l166_411 = {1'd0, _zz_when_ArraySlice_l166_411_1};
  assign _zz_when_ArraySlice_l166_411_2 = (_zz_when_ArraySlice_l166_411_3 + _zz_when_ArraySlice_l166_411_7);
  assign _zz_when_ArraySlice_l166_411_3 = (realValue_0_411 - _zz_when_ArraySlice_l166_411_4);
  assign _zz_when_ArraySlice_l166_411_4 = (selectReadFifo_3 + _zz_when_ArraySlice_l166_411_5);
  assign _zz_when_ArraySlice_l166_411_6 = (bReg * 2'b11);
  assign _zz_when_ArraySlice_l166_411_5 = {2'd0, _zz_when_ArraySlice_l166_411_6};
  assign _zz_when_ArraySlice_l166_411_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_412 = (selectReadFifo_4 + _zz_when_ArraySlice_l158_412_1);
  assign _zz_when_ArraySlice_l158_412_2 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l158_412_1 = {1'd0, _zz_when_ArraySlice_l158_412_2};
  assign _zz_when_ArraySlice_l158_412_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_412_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l159_412 = {1'd0, _zz_when_ArraySlice_l159_412_1};
  assign _zz_when_ArraySlice_l159_412_2 = (_zz_when_ArraySlice_l159_412_3 - _zz_when_ArraySlice_l159_412_4);
  assign _zz_when_ArraySlice_l159_412_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_412_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l159_412_5);
  assign _zz_when_ArraySlice_l159_412_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l159_412_5 = {1'd0, _zz_when_ArraySlice_l159_412_6};
  assign _zz__zz_realValue_0_412 = {1'd0, wReg};
  assign _zz__zz_realValue_0_412_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_412_1 = (_zz_realValue_0_412_2 + _zz_realValue_0_412_3);
  assign _zz_realValue_0_412_2 = {1'd0, wReg};
  assign _zz_realValue_0_412_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_412_1 = (3'b100 * bReg);
  assign _zz_when_ArraySlice_l166_412 = {1'd0, _zz_when_ArraySlice_l166_412_1};
  assign _zz_when_ArraySlice_l166_412_2 = (_zz_when_ArraySlice_l166_412_3 + _zz_when_ArraySlice_l166_412_7);
  assign _zz_when_ArraySlice_l166_412_3 = (realValue_0_412 - _zz_when_ArraySlice_l166_412_4);
  assign _zz_when_ArraySlice_l166_412_4 = (selectReadFifo_4 + _zz_when_ArraySlice_l166_412_5);
  assign _zz_when_ArraySlice_l166_412_6 = (bReg * 3'b100);
  assign _zz_when_ArraySlice_l166_412_5 = {1'd0, _zz_when_ArraySlice_l166_412_6};
  assign _zz_when_ArraySlice_l166_412_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_413 = (selectReadFifo_5 + _zz_when_ArraySlice_l158_413_1);
  assign _zz_when_ArraySlice_l158_413_2 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l158_413_1 = {1'd0, _zz_when_ArraySlice_l158_413_2};
  assign _zz_when_ArraySlice_l158_413_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_413_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l159_413 = {2'd0, _zz_when_ArraySlice_l159_413_1};
  assign _zz_when_ArraySlice_l159_413_2 = (_zz_when_ArraySlice_l159_413_3 - _zz_when_ArraySlice_l159_413_4);
  assign _zz_when_ArraySlice_l159_413_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_413_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l159_413_5);
  assign _zz_when_ArraySlice_l159_413_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l159_413_5 = {1'd0, _zz_when_ArraySlice_l159_413_6};
  assign _zz__zz_realValue_0_413 = {1'd0, wReg};
  assign _zz__zz_realValue_0_413_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_413_1 = (_zz_realValue_0_413_2 + _zz_realValue_0_413_3);
  assign _zz_realValue_0_413_2 = {1'd0, wReg};
  assign _zz_realValue_0_413_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_413_1 = (2'b11 * bReg);
  assign _zz_when_ArraySlice_l166_413 = {2'd0, _zz_when_ArraySlice_l166_413_1};
  assign _zz_when_ArraySlice_l166_413_2 = (_zz_when_ArraySlice_l166_413_3 + _zz_when_ArraySlice_l166_413_7);
  assign _zz_when_ArraySlice_l166_413_3 = (realValue_0_413 - _zz_when_ArraySlice_l166_413_4);
  assign _zz_when_ArraySlice_l166_413_4 = (selectReadFifo_5 + _zz_when_ArraySlice_l166_413_5);
  assign _zz_when_ArraySlice_l166_413_6 = (bReg * 3'b101);
  assign _zz_when_ArraySlice_l166_413_5 = {1'd0, _zz_when_ArraySlice_l166_413_6};
  assign _zz_when_ArraySlice_l166_413_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_414 = (selectReadFifo_6 + _zz_when_ArraySlice_l158_414_1);
  assign _zz_when_ArraySlice_l158_414_2 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l158_414_1 = {1'd0, _zz_when_ArraySlice_l158_414_2};
  assign _zz_when_ArraySlice_l158_414_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_414_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l159_414 = {2'd0, _zz_when_ArraySlice_l159_414_1};
  assign _zz_when_ArraySlice_l159_414_2 = (_zz_when_ArraySlice_l159_414_3 - _zz_when_ArraySlice_l159_414_4);
  assign _zz_when_ArraySlice_l159_414_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_414_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l159_414_5);
  assign _zz_when_ArraySlice_l159_414_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l159_414_5 = {1'd0, _zz_when_ArraySlice_l159_414_6};
  assign _zz__zz_realValue_0_414 = {1'd0, wReg};
  assign _zz__zz_realValue_0_414_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_414_1 = (_zz_realValue_0_414_2 + _zz_realValue_0_414_3);
  assign _zz_realValue_0_414_2 = {1'd0, wReg};
  assign _zz_realValue_0_414_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_414_1 = (2'b10 * bReg);
  assign _zz_when_ArraySlice_l166_414 = {2'd0, _zz_when_ArraySlice_l166_414_1};
  assign _zz_when_ArraySlice_l166_414_2 = (_zz_when_ArraySlice_l166_414_3 + _zz_when_ArraySlice_l166_414_7);
  assign _zz_when_ArraySlice_l166_414_3 = (realValue_0_414 - _zz_when_ArraySlice_l166_414_4);
  assign _zz_when_ArraySlice_l166_414_4 = (selectReadFifo_6 + _zz_when_ArraySlice_l166_414_5);
  assign _zz_when_ArraySlice_l166_414_6 = (bReg * 3'b110);
  assign _zz_when_ArraySlice_l166_414_5 = {1'd0, _zz_when_ArraySlice_l166_414_6};
  assign _zz_when_ArraySlice_l166_414_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l158_415 = (selectReadFifo_7 + _zz_when_ArraySlice_l158_415_1);
  assign _zz_when_ArraySlice_l158_415_2 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l158_415_1 = {1'd0, _zz_when_ArraySlice_l158_415_2};
  assign _zz_when_ArraySlice_l158_415_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_415_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l159_415 = {3'd0, _zz_when_ArraySlice_l159_415_1};
  assign _zz_when_ArraySlice_l159_415_2 = (_zz_when_ArraySlice_l159_415_3 - _zz_when_ArraySlice_l159_415_4);
  assign _zz_when_ArraySlice_l159_415_3 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l159_415_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l159_415_5);
  assign _zz_when_ArraySlice_l159_415_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l159_415_5 = {1'd0, _zz_when_ArraySlice_l159_415_6};
  assign _zz__zz_realValue_0_415 = {1'd0, wReg};
  assign _zz__zz_realValue_0_415_1 = (bReg * 4'b1000);
  assign _zz_realValue_0_415_1 = (_zz_realValue_0_415_2 + _zz_realValue_0_415_3);
  assign _zz_realValue_0_415_2 = {1'd0, wReg};
  assign _zz_realValue_0_415_3 = (bReg * 4'b1000);
  assign _zz_when_ArraySlice_l166_415_1 = (1'b1 * bReg);
  assign _zz_when_ArraySlice_l166_415 = {3'd0, _zz_when_ArraySlice_l166_415_1};
  assign _zz_when_ArraySlice_l166_415_2 = (_zz_when_ArraySlice_l166_415_3 + _zz_when_ArraySlice_l166_415_7);
  assign _zz_when_ArraySlice_l166_415_3 = (realValue_0_415 - _zz_when_ArraySlice_l166_415_4);
  assign _zz_when_ArraySlice_l166_415_4 = (selectReadFifo_7 + _zz_when_ArraySlice_l166_415_5);
  assign _zz_when_ArraySlice_l166_415_6 = (bReg * 3'b111);
  assign _zz_when_ArraySlice_l166_415_5 = {1'd0, _zz_when_ArraySlice_l166_415_6};
  assign _zz_when_ArraySlice_l166_415_7 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_8 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_8_1 = (selectReadFifo_0 - _zz_when_ArraySlice_l182_8_2);
  assign _zz_when_ArraySlice_l182_8_2 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l182_9 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_9_1 = (selectReadFifo_1 - _zz_when_ArraySlice_l182_9_2);
  assign _zz_when_ArraySlice_l182_9_2 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l182_10 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_10_1 = (selectReadFifo_2 - _zz_when_ArraySlice_l182_10_2);
  assign _zz_when_ArraySlice_l182_10_2 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l182_11 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_11_1 = (selectReadFifo_3 - _zz_when_ArraySlice_l182_11_2);
  assign _zz_when_ArraySlice_l182_11_2 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l182_12 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_12_1 = (selectReadFifo_4 - _zz_when_ArraySlice_l182_12_2);
  assign _zz_when_ArraySlice_l182_12_2 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l182_13 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_13_1 = (selectReadFifo_5 - _zz_when_ArraySlice_l182_13_2);
  assign _zz_when_ArraySlice_l182_13_2 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l182_14 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_14_1 = (selectReadFifo_6 - _zz_when_ArraySlice_l182_14_2);
  assign _zz_when_ArraySlice_l182_14_2 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l182_15 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_15_1 = (selectReadFifo_7 - _zz_when_ArraySlice_l182_15_2);
  assign _zz_when_ArraySlice_l182_15_2 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l182_16 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_16_1 = (selectReadFifo_0 - _zz_when_ArraySlice_l182_16_2);
  assign _zz_when_ArraySlice_l182_16_2 = (selectReadFifo_0 % bReg);
  assign _zz_when_ArraySlice_l182_17 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_17_1 = (selectReadFifo_1 - _zz_when_ArraySlice_l182_17_2);
  assign _zz_when_ArraySlice_l182_17_2 = (selectReadFifo_1 % bReg);
  assign _zz_when_ArraySlice_l182_18 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_18_1 = (selectReadFifo_2 - _zz_when_ArraySlice_l182_18_2);
  assign _zz_when_ArraySlice_l182_18_2 = (selectReadFifo_2 % bReg);
  assign _zz_when_ArraySlice_l182_19 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_19_1 = (selectReadFifo_3 - _zz_when_ArraySlice_l182_19_2);
  assign _zz_when_ArraySlice_l182_19_2 = (selectReadFifo_3 % bReg);
  assign _zz_when_ArraySlice_l182_20 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_20_1 = (selectReadFifo_4 - _zz_when_ArraySlice_l182_20_2);
  assign _zz_when_ArraySlice_l182_20_2 = (selectReadFifo_4 % bReg);
  assign _zz_when_ArraySlice_l182_21 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_21_1 = (selectReadFifo_5 - _zz_when_ArraySlice_l182_21_2);
  assign _zz_when_ArraySlice_l182_21_2 = (selectReadFifo_5 % bReg);
  assign _zz_when_ArraySlice_l182_22 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_22_1 = (selectReadFifo_6 - _zz_when_ArraySlice_l182_22_2);
  assign _zz_when_ArraySlice_l182_22_2 = (selectReadFifo_6 % bReg);
  assign _zz_when_ArraySlice_l182_23 = {1'd0, selectWriteFifo};
  assign _zz_when_ArraySlice_l182_23_1 = (selectReadFifo_7 - _zz_when_ArraySlice_l182_23_2);
  assign _zz_when_ArraySlice_l182_23_2 = (selectReadFifo_7 % bReg);
  assign _zz_when_ArraySlice_l400 = ((((holdReadOp_0 == _zz_when_ArraySlice_l400_1) && (holdReadOp_1 == _zz_when_ArraySlice_l400_2)) && (holdReadOp_2 == 1'b1)) && (holdReadOp_3 == 1'b1));
  assign _zz_when_ArraySlice_l400_3 = (holdReadOp_4 == 1'b1);
  assign _zz_when_ArraySlice_l400_4 = 1'b1;
  assign _zz_when_ArraySlice_l400_5 = ((((debug_0_1 == _zz_when_ArraySlice_l400_6) && (debug_1_1 == _zz_when_ArraySlice_l400_7)) && (debug_2_1 == 1'b1)) && (debug_3_1 == 1'b1));
  assign _zz_when_ArraySlice_l400_8 = (debug_4_1 == 1'b1);
  assign _zz_when_ArraySlice_l400_9 = 1'b1;
  assign _zz_when_ArraySlice_l400_1 = 1'b1;
  assign _zz_when_ArraySlice_l400_2 = 1'b1;
  assign _zz_when_ArraySlice_l400_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_7 = 1'b1;
  assign _zz_when_ArraySlice_l425 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_2 = 1'b1;
  assign _zz_when_ArraySlice_l425_3 = (((debug_0_2 == 1'b1) && (debug_1_2 == 1'b1)) && (debug_2_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_4 = (debug_3_2 == 1'b1);
  assign _zz_when_ArraySlice_l425_5 = 1'b1;
  assign _zz_when_ArraySlice_l457 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_2 = 1'b1;
  assign _zz_when_ArraySlice_l457_3 = (((debug_0_3 == 1'b1) && (debug_1_3 == 1'b1)) && (debug_2_3 == 1'b1));
  assign _zz_when_ArraySlice_l457_4 = (debug_3_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_5 = 1'b1;
  assign _zz_when_ArraySlice_l400_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_1_4 = (((debug_0_4 == 1'b1) && (debug_1_4 == 1'b1)) && (debug_2_4 == 1'b1));
  assign _zz_when_ArraySlice_l400_1_5 = (debug_3_4 == 1'b1);
  assign _zz_when_ArraySlice_l400_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_1_4 = (((debug_0_5 == 1'b1) && (debug_1_5 == 1'b1)) && (debug_2_5 == 1'b1));
  assign _zz_when_ArraySlice_l425_1_5 = (debug_3_5 == 1'b1);
  assign _zz_when_ArraySlice_l425_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l457_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l457_1_4 = (((debug_0_6 == 1'b1) && (debug_1_6 == 1'b1)) && (debug_2_6 == 1'b1));
  assign _zz_when_ArraySlice_l457_1_5 = (debug_3_6 == 1'b1);
  assign _zz_when_ArraySlice_l457_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_2_4 = (((debug_0_7 == 1'b1) && (debug_1_7 == 1'b1)) && (debug_2_7 == 1'b1));
  assign _zz_when_ArraySlice_l400_2_5 = (debug_3_7 == 1'b1);
  assign _zz_when_ArraySlice_l400_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_2_4 = (((debug_0_8 == 1'b1) && (debug_1_8 == 1'b1)) && (debug_2_8 == 1'b1));
  assign _zz_when_ArraySlice_l425_2_5 = (debug_3_8 == 1'b1);
  assign _zz_when_ArraySlice_l425_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l457_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l457_2_4 = (((debug_0_9 == 1'b1) && (debug_1_9 == 1'b1)) && (debug_2_9 == 1'b1));
  assign _zz_when_ArraySlice_l457_2_5 = (debug_3_9 == 1'b1);
  assign _zz_when_ArraySlice_l457_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_3_4 = (((debug_0_10 == 1'b1) && (debug_1_10 == 1'b1)) && (debug_2_10 == 1'b1));
  assign _zz_when_ArraySlice_l400_3_5 = (debug_3_10 == 1'b1);
  assign _zz_when_ArraySlice_l400_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_3_4 = (((debug_0_11 == 1'b1) && (debug_1_11 == 1'b1)) && (debug_2_11 == 1'b1));
  assign _zz_when_ArraySlice_l425_3_5 = (debug_3_11 == 1'b1);
  assign _zz_when_ArraySlice_l425_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l457_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l457_3_4 = (((debug_0_12 == 1'b1) && (debug_1_12 == 1'b1)) && (debug_2_12 == 1'b1));
  assign _zz_when_ArraySlice_l457_3_5 = (debug_3_12 == 1'b1);
  assign _zz_when_ArraySlice_l457_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_4_4 = (((debug_0_13 == 1'b1) && (debug_1_13 == 1'b1)) && (debug_2_13 == 1'b1));
  assign _zz_when_ArraySlice_l400_4_5 = (debug_3_13 == 1'b1);
  assign _zz_when_ArraySlice_l400_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_4_4 = (((debug_0_14 == 1'b1) && (debug_1_14 == 1'b1)) && (debug_2_14 == 1'b1));
  assign _zz_when_ArraySlice_l425_4_5 = (debug_3_14 == 1'b1);
  assign _zz_when_ArraySlice_l425_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l457_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l457_4_4 = (((debug_0_15 == 1'b1) && (debug_1_15 == 1'b1)) && (debug_2_15 == 1'b1));
  assign _zz_when_ArraySlice_l457_4_5 = (debug_3_15 == 1'b1);
  assign _zz_when_ArraySlice_l457_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_5_4 = (((debug_0_16 == 1'b1) && (debug_1_16 == 1'b1)) && (debug_2_16 == 1'b1));
  assign _zz_when_ArraySlice_l400_5_5 = (debug_3_16 == 1'b1);
  assign _zz_when_ArraySlice_l400_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l425_5_4 = (((debug_0_17 == 1'b1) && (debug_1_17 == 1'b1)) && (debug_2_17 == 1'b1));
  assign _zz_when_ArraySlice_l425_5_5 = (debug_3_17 == 1'b1);
  assign _zz_when_ArraySlice_l425_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l457_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l457_5_4 = (((debug_0_18 == 1'b1) && (debug_1_18 == 1'b1)) && (debug_2_18 == 1'b1));
  assign _zz_when_ArraySlice_l457_5_5 = (debug_3_18 == 1'b1);
  assign _zz_when_ArraySlice_l457_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l400_6_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_6_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_6_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_6_4 = (((debug_0_19 == 1'b1) && (debug_1_19 == 1'b1)) && (debug_2_19 == 1'b1));
  assign _zz_when_ArraySlice_l400_6_5 = (debug_3_19 == 1'b1);
  assign _zz_when_ArraySlice_l400_6_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l425_6_3 = (((debug_0_20 == 1'b1) && (debug_1_20 == 1'b1)) && (debug_2_20 == 1'b1));
  assign _zz_when_ArraySlice_l425_6_4 = (debug_3_20 == 1'b1);
  assign _zz_when_ArraySlice_l425_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l457_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l457_6_3 = (((debug_0_21 == 1'b1) && (debug_1_21 == 1'b1)) && (debug_2_21 == 1'b1));
  assign _zz_when_ArraySlice_l457_6_4 = (debug_3_21 == 1'b1);
  assign _zz_when_ArraySlice_l457_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l400_7_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l400_7_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l400_7_3 = 1'b1;
  assign _zz_when_ArraySlice_l400_7_4 = (((debug_0_22 == 1'b1) && (debug_1_22 == 1'b1)) && (debug_2_22 == 1'b1));
  assign _zz_when_ArraySlice_l400_7_5 = (debug_3_22 == 1'b1);
  assign _zz_when_ArraySlice_l400_7_6 = 1'b1;
  assign _zz_when_ArraySlice_l425_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l425_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l425_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l425_7_3 = (((debug_0_23 == 1'b1) && (debug_1_23 == 1'b1)) && (debug_2_23 == 1'b1));
  assign _zz_when_ArraySlice_l425_7_4 = (debug_3_23 == 1'b1);
  assign _zz_when_ArraySlice_l425_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l457_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l457_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l457_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l457_7_3 = (((debug_0_24 == 1'b1) && (debug_1_24 == 1'b1)) && (debug_2_24 == 1'b1));
  assign _zz_when_ArraySlice_l457_7_4 = (debug_3_24 == 1'b1);
  assign _zz_when_ArraySlice_l457_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l478 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l478_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l478_2 = 1'b1;
  assign _zz_when_ArraySlice_l478_3 = (((debug_0_25 == 1'b1) && (debug_1_25 == 1'b1)) && (debug_2_25 == 1'b1));
  assign _zz_when_ArraySlice_l478_4 = (debug_3_25 == 1'b1);
  assign _zz_when_ArraySlice_l478_5 = 1'b1;
  assign _zz_when_ArraySlice_l257 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_2 = 1'b1;
  assign _zz_when_ArraySlice_l257_3 = (((debug_0_26 == 1'b1) && (debug_1_26 == 1'b1)) && (debug_2_26 == 1'b1));
  assign _zz_when_ArraySlice_l257_4 = (debug_3_26 == 1'b1);
  assign _zz_when_ArraySlice_l257_5 = 1'b1;
  assign _zz_when_ArraySlice_l282 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_2 = 1'b1;
  assign _zz_when_ArraySlice_l282_3 = (((debug_0_27 == 1'b1) && (debug_1_27 == 1'b1)) && (debug_2_27 == 1'b1));
  assign _zz_when_ArraySlice_l282_4 = (debug_3_27 == 1'b1);
  assign _zz_when_ArraySlice_l282_5 = 1'b1;
  assign _zz_when_ArraySlice_l314 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_2 = 1'b1;
  assign _zz_when_ArraySlice_l314_3 = (((debug_0_28 == 1'b1) && (debug_1_28 == 1'b1)) && (debug_2_28 == 1'b1));
  assign _zz_when_ArraySlice_l314_4 = (debug_3_28 == 1'b1);
  assign _zz_when_ArraySlice_l314_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l257_1_4 = (((debug_0_29 == 1'b1) && (debug_1_29 == 1'b1)) && (debug_2_29 == 1'b1));
  assign _zz_when_ArraySlice_l257_1_5 = (debug_3_29 == 1'b1);
  assign _zz_when_ArraySlice_l257_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l282_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l282_1_4 = (((debug_0_30 == 1'b1) && (debug_1_30 == 1'b1)) && (debug_2_30 == 1'b1));
  assign _zz_when_ArraySlice_l282_1_5 = (debug_3_30 == 1'b1);
  assign _zz_when_ArraySlice_l282_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l314_1_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_1_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_1_3 = 1'b1;
  assign _zz_when_ArraySlice_l314_1_4 = (((debug_0_31 == 1'b1) && (debug_1_31 == 1'b1)) && (debug_2_31 == 1'b1));
  assign _zz_when_ArraySlice_l314_1_5 = (debug_3_31 == 1'b1);
  assign _zz_when_ArraySlice_l314_1_6 = 1'b1;
  assign _zz_when_ArraySlice_l257_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l257_2_4 = (((debug_0_32 == 1'b1) && (debug_1_32 == 1'b1)) && (debug_2_32 == 1'b1));
  assign _zz_when_ArraySlice_l257_2_5 = (debug_3_32 == 1'b1);
  assign _zz_when_ArraySlice_l257_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l282_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l282_2_4 = (((debug_0_33 == 1'b1) && (debug_1_33 == 1'b1)) && (debug_2_33 == 1'b1));
  assign _zz_when_ArraySlice_l282_2_5 = (debug_3_33 == 1'b1);
  assign _zz_when_ArraySlice_l282_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l314_2_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_2_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_2_3 = 1'b1;
  assign _zz_when_ArraySlice_l314_2_4 = (((debug_0_34 == 1'b1) && (debug_1_34 == 1'b1)) && (debug_2_34 == 1'b1));
  assign _zz_when_ArraySlice_l314_2_5 = (debug_3_34 == 1'b1);
  assign _zz_when_ArraySlice_l314_2_6 = 1'b1;
  assign _zz_when_ArraySlice_l257_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l257_3_4 = (((debug_0_35 == 1'b1) && (debug_1_35 == 1'b1)) && (debug_2_35 == 1'b1));
  assign _zz_when_ArraySlice_l257_3_5 = (debug_3_35 == 1'b1);
  assign _zz_when_ArraySlice_l257_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l282_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l282_3_4 = (((debug_0_36 == 1'b1) && (debug_1_36 == 1'b1)) && (debug_2_36 == 1'b1));
  assign _zz_when_ArraySlice_l282_3_5 = (debug_3_36 == 1'b1);
  assign _zz_when_ArraySlice_l282_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l314_3_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_3_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_3_3 = 1'b1;
  assign _zz_when_ArraySlice_l314_3_4 = (((debug_0_37 == 1'b1) && (debug_1_37 == 1'b1)) && (debug_2_37 == 1'b1));
  assign _zz_when_ArraySlice_l314_3_5 = (debug_3_37 == 1'b1);
  assign _zz_when_ArraySlice_l314_3_6 = 1'b1;
  assign _zz_when_ArraySlice_l257_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l257_4_4 = (((debug_0_38 == 1'b1) && (debug_1_38 == 1'b1)) && (debug_2_38 == 1'b1));
  assign _zz_when_ArraySlice_l257_4_5 = (debug_3_38 == 1'b1);
  assign _zz_when_ArraySlice_l257_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l282_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l282_4_4 = (((debug_0_39 == 1'b1) && (debug_1_39 == 1'b1)) && (debug_2_39 == 1'b1));
  assign _zz_when_ArraySlice_l282_4_5 = (debug_3_39 == 1'b1);
  assign _zz_when_ArraySlice_l282_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l314_4_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_4_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_4_3 = 1'b1;
  assign _zz_when_ArraySlice_l314_4_4 = (((debug_0_40 == 1'b1) && (debug_1_40 == 1'b1)) && (debug_2_40 == 1'b1));
  assign _zz_when_ArraySlice_l314_4_5 = (debug_3_40 == 1'b1);
  assign _zz_when_ArraySlice_l314_4_6 = 1'b1;
  assign _zz_when_ArraySlice_l257_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l257_5_4 = (((debug_0_41 == 1'b1) && (debug_1_41 == 1'b1)) && (debug_2_41 == 1'b1));
  assign _zz_when_ArraySlice_l257_5_5 = (debug_3_41 == 1'b1);
  assign _zz_when_ArraySlice_l257_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l282_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l282_5_4 = (((debug_0_42 == 1'b1) && (debug_1_42 == 1'b1)) && (debug_2_42 == 1'b1));
  assign _zz_when_ArraySlice_l282_5_5 = (debug_3_42 == 1'b1);
  assign _zz_when_ArraySlice_l282_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l314_5_1 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_5_2 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_5_3 = 1'b1;
  assign _zz_when_ArraySlice_l314_5_4 = (((debug_0_43 == 1'b1) && (debug_1_43 == 1'b1)) && (debug_2_43 == 1'b1));
  assign _zz_when_ArraySlice_l314_5_5 = (debug_3_43 == 1'b1);
  assign _zz_when_ArraySlice_l314_5_6 = 1'b1;
  assign _zz_when_ArraySlice_l257_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l257_6_3 = (((debug_0_44 == 1'b1) && (debug_1_44 == 1'b1)) && (debug_2_44 == 1'b1));
  assign _zz_when_ArraySlice_l257_6_4 = (debug_3_44 == 1'b1);
  assign _zz_when_ArraySlice_l257_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l282_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l282_6_3 = (((debug_0_45 == 1'b1) && (debug_1_45 == 1'b1)) && (debug_2_45 == 1'b1));
  assign _zz_when_ArraySlice_l282_6_4 = (debug_3_45 == 1'b1);
  assign _zz_when_ArraySlice_l282_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l314_6 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_6_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_6_2 = 1'b1;
  assign _zz_when_ArraySlice_l314_6_3 = (((debug_0_46 == 1'b1) && (debug_1_46 == 1'b1)) && (debug_2_46 == 1'b1));
  assign _zz_when_ArraySlice_l314_6_4 = (debug_3_46 == 1'b1);
  assign _zz_when_ArraySlice_l314_6_5 = 1'b1;
  assign _zz_when_ArraySlice_l257_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l257_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l257_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l257_7_3 = (((debug_0_47 == 1'b1) && (debug_1_47 == 1'b1)) && (debug_2_47 == 1'b1));
  assign _zz_when_ArraySlice_l257_7_4 = (debug_3_47 == 1'b1);
  assign _zz_when_ArraySlice_l257_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l282_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l282_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l282_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l282_7_3 = (((debug_0_48 == 1'b1) && (debug_1_48 == 1'b1)) && (debug_2_48 == 1'b1));
  assign _zz_when_ArraySlice_l282_7_4 = (debug_3_48 == 1'b1);
  assign _zz_when_ArraySlice_l282_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l314_7 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l314_7_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l314_7_2 = 1'b1;
  assign _zz_when_ArraySlice_l314_7_3 = (((debug_0_49 == 1'b1) && (debug_1_49 == 1'b1)) && (debug_2_49 == 1'b1));
  assign _zz_when_ArraySlice_l314_7_4 = (debug_3_49 == 1'b1);
  assign _zz_when_ArraySlice_l314_7_5 = 1'b1;
  assign _zz_when_ArraySlice_l336_8 = 1'b0;
  assign _zz_when_ArraySlice_l336_9 = 1'b0;
  assign _zz_when_ArraySlice_l353 = (((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1)) && (holdReadOp_2 == 1'b1));
  assign _zz_when_ArraySlice_l353_1 = (holdReadOp_3 == 1'b1);
  assign _zz_when_ArraySlice_l353_2 = 1'b1;
  assign _zz_when_ArraySlice_l353_3 = (((debug_0_50 == 1'b1) && (debug_1_50 == 1'b1)) && (debug_2_50 == 1'b1));
  assign _zz_when_ArraySlice_l353_4 = (debug_3_50 == 1'b1);
  assign _zz_when_ArraySlice_l353_5 = 1'b1;
  assign _zz_when_ArraySlice_l357_8 = (((_zz_when_ArraySlice_l357_9 && _zz_when_ArraySlice_l357_10) && (holdReadOp_3 == _zz_when_ArraySlice_l357_11)) && (holdReadOp_4 == 1'b1));
  assign _zz_when_ArraySlice_l357_12 = (holdReadOp_5 == 1'b1);
  assign _zz_when_ArraySlice_l357_13 = 1'b1;
  assign _zz_when_ArraySlice_l357_14 = (((_zz_when_ArraySlice_l357_15 && _zz_when_ArraySlice_l357_16) && (debug_4_51 == _zz_when_ArraySlice_l357_17)) && (debug_5_51 == 1'b1));
  assign _zz_when_ArraySlice_l357_18 = (debug_6_51 == 1'b1);
  assign _zz_when_ArraySlice_l357_19 = 1'b1;
  assign _zz_when_ArraySlice_l357_20 = (((_zz_when_ArraySlice_l357_21 || _zz_when_ArraySlice_l357_22) || (_zz_when_ArraySlice_l357_3 != _zz_when_ArraySlice_l357_23)) || (_zz_when_ArraySlice_l357_4 != 1'b0));
  assign _zz_when_ArraySlice_l357_24 = (_zz_when_ArraySlice_l357_5 != 1'b0);
  assign _zz_when_ArraySlice_l357_25 = 1'b0;
  assign _zz_when_ArraySlice_l357_9 = ((holdReadOp_0 == 1'b1) && (holdReadOp_1 == 1'b1));
  assign _zz_when_ArraySlice_l357_10 = (holdReadOp_2 == 1'b1);
  assign _zz_when_ArraySlice_l357_11 = 1'b1;
  assign _zz_when_ArraySlice_l357_15 = (((debug_0_51 == 1'b1) && (debug_1_51 == 1'b1)) && (debug_2_51 == 1'b1));
  assign _zz_when_ArraySlice_l357_16 = (debug_3_51 == 1'b1);
  assign _zz_when_ArraySlice_l357_17 = 1'b1;
  assign _zz_when_ArraySlice_l357_21 = ((_zz_when_ArraySlice_l357 != 1'b0) || (_zz_when_ArraySlice_l357_1 != 1'b0));
  assign _zz_when_ArraySlice_l357_22 = (_zz_when_ArraySlice_l357_2 != 1'b0);
  assign _zz_when_ArraySlice_l357_23 = 1'b0;
  StreamFifo fifoGroup_0 (
    .io_push_valid   (fifoGroup_0_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_0_io_push_ready        ), //o
    .io_push_payload (fifoGroup_0_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_0_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_0_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_0_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_0_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_0_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_1 (
    .io_push_valid   (fifoGroup_1_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_1_io_push_ready        ), //o
    .io_push_payload (fifoGroup_1_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_1_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_1_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_1_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_1_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_1_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_2 (
    .io_push_valid   (fifoGroup_2_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_2_io_push_ready        ), //o
    .io_push_payload (fifoGroup_2_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_2_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_2_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_2_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_2_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_2_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_3 (
    .io_push_valid   (fifoGroup_3_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_3_io_push_ready        ), //o
    .io_push_payload (fifoGroup_3_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_3_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_3_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_3_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_3_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_3_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_4 (
    .io_push_valid   (fifoGroup_4_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_4_io_push_ready        ), //o
    .io_push_payload (fifoGroup_4_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_4_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_4_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_4_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_4_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_4_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_5 (
    .io_push_valid   (fifoGroup_5_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_5_io_push_ready        ), //o
    .io_push_payload (fifoGroup_5_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_5_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_5_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_5_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_5_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_5_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_6 (
    .io_push_valid   (fifoGroup_6_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_6_io_push_ready        ), //o
    .io_push_payload (fifoGroup_6_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_6_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_6_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_6_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_6_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_6_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_7 (
    .io_push_valid   (fifoGroup_7_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_7_io_push_ready        ), //o
    .io_push_payload (fifoGroup_7_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_7_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_7_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_7_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_7_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_7_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_8 (
    .io_push_valid   (fifoGroup_8_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_8_io_push_ready        ), //o
    .io_push_payload (fifoGroup_8_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_8_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_8_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_8_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_8_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_8_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_9 (
    .io_push_valid   (fifoGroup_9_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_9_io_push_ready        ), //o
    .io_push_payload (fifoGroup_9_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_9_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_9_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_9_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                             ), //i
    .io_occupancy    (fifoGroup_9_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_9_io_availability[6:0] ), //o
    .clk             (clk                              ), //i
    .resetn          (resetn                           )  //i
  );
  StreamFifo fifoGroup_10 (
    .io_push_valid   (fifoGroup_10_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_10_io_push_ready        ), //o
    .io_push_payload (fifoGroup_10_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_10_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_10_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_10_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_10_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_10_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_11 (
    .io_push_valid   (fifoGroup_11_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_11_io_push_ready        ), //o
    .io_push_payload (fifoGroup_11_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_11_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_11_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_11_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_11_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_11_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_12 (
    .io_push_valid   (fifoGroup_12_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_12_io_push_ready        ), //o
    .io_push_payload (fifoGroup_12_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_12_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_12_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_12_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_12_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_12_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_13 (
    .io_push_valid   (fifoGroup_13_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_13_io_push_ready        ), //o
    .io_push_payload (fifoGroup_13_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_13_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_13_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_13_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_13_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_13_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_14 (
    .io_push_valid   (fifoGroup_14_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_14_io_push_ready        ), //o
    .io_push_payload (fifoGroup_14_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_14_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_14_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_14_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_14_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_14_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_15 (
    .io_push_valid   (fifoGroup_15_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_15_io_push_ready        ), //o
    .io_push_payload (fifoGroup_15_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_15_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_15_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_15_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_15_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_15_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_16 (
    .io_push_valid   (fifoGroup_16_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_16_io_push_ready        ), //o
    .io_push_payload (fifoGroup_16_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_16_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_16_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_16_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_16_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_16_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_17 (
    .io_push_valid   (fifoGroup_17_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_17_io_push_ready        ), //o
    .io_push_payload (fifoGroup_17_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_17_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_17_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_17_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_17_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_17_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_18 (
    .io_push_valid   (fifoGroup_18_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_18_io_push_ready        ), //o
    .io_push_payload (fifoGroup_18_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_18_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_18_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_18_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_18_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_18_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_19 (
    .io_push_valid   (fifoGroup_19_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_19_io_push_ready        ), //o
    .io_push_payload (fifoGroup_19_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_19_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_19_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_19_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_19_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_19_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_20 (
    .io_push_valid   (fifoGroup_20_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_20_io_push_ready        ), //o
    .io_push_payload (fifoGroup_20_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_20_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_20_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_20_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_20_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_20_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_21 (
    .io_push_valid   (fifoGroup_21_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_21_io_push_ready        ), //o
    .io_push_payload (fifoGroup_21_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_21_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_21_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_21_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_21_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_21_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_22 (
    .io_push_valid   (fifoGroup_22_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_22_io_push_ready        ), //o
    .io_push_payload (fifoGroup_22_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_22_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_22_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_22_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_22_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_22_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_23 (
    .io_push_valid   (fifoGroup_23_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_23_io_push_ready        ), //o
    .io_push_payload (fifoGroup_23_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_23_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_23_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_23_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_23_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_23_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_24 (
    .io_push_valid   (fifoGroup_24_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_24_io_push_ready        ), //o
    .io_push_payload (fifoGroup_24_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_24_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_24_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_24_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_24_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_24_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_25 (
    .io_push_valid   (fifoGroup_25_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_25_io_push_ready        ), //o
    .io_push_payload (fifoGroup_25_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_25_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_25_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_25_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_25_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_25_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_26 (
    .io_push_valid   (fifoGroup_26_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_26_io_push_ready        ), //o
    .io_push_payload (fifoGroup_26_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_26_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_26_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_26_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_26_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_26_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_27 (
    .io_push_valid   (fifoGroup_27_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_27_io_push_ready        ), //o
    .io_push_payload (fifoGroup_27_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_27_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_27_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_27_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_27_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_27_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_28 (
    .io_push_valid   (fifoGroup_28_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_28_io_push_ready        ), //o
    .io_push_payload (fifoGroup_28_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_28_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_28_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_28_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_28_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_28_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_29 (
    .io_push_valid   (fifoGroup_29_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_29_io_push_ready        ), //o
    .io_push_payload (fifoGroup_29_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_29_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_29_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_29_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_29_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_29_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_30 (
    .io_push_valid   (fifoGroup_30_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_30_io_push_ready        ), //o
    .io_push_payload (fifoGroup_30_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_30_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_30_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_30_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_30_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_30_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_31 (
    .io_push_valid   (fifoGroup_31_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_31_io_push_ready        ), //o
    .io_push_payload (fifoGroup_31_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_31_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_31_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_31_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_31_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_31_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_32 (
    .io_push_valid   (fifoGroup_32_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_32_io_push_ready        ), //o
    .io_push_payload (fifoGroup_32_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_32_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_32_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_32_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_32_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_32_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_33 (
    .io_push_valid   (fifoGroup_33_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_33_io_push_ready        ), //o
    .io_push_payload (fifoGroup_33_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_33_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_33_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_33_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_33_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_33_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_34 (
    .io_push_valid   (fifoGroup_34_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_34_io_push_ready        ), //o
    .io_push_payload (fifoGroup_34_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_34_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_34_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_34_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_34_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_34_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_35 (
    .io_push_valid   (fifoGroup_35_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_35_io_push_ready        ), //o
    .io_push_payload (fifoGroup_35_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_35_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_35_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_35_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_35_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_35_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_36 (
    .io_push_valid   (fifoGroup_36_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_36_io_push_ready        ), //o
    .io_push_payload (fifoGroup_36_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_36_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_36_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_36_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_36_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_36_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_37 (
    .io_push_valid   (fifoGroup_37_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_37_io_push_ready        ), //o
    .io_push_payload (fifoGroup_37_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_37_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_37_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_37_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_37_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_37_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_38 (
    .io_push_valid   (fifoGroup_38_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_38_io_push_ready        ), //o
    .io_push_payload (fifoGroup_38_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_38_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_38_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_38_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_38_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_38_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_39 (
    .io_push_valid   (fifoGroup_39_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_39_io_push_ready        ), //o
    .io_push_payload (fifoGroup_39_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_39_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_39_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_39_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_39_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_39_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_40 (
    .io_push_valid   (fifoGroup_40_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_40_io_push_ready        ), //o
    .io_push_payload (fifoGroup_40_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_40_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_40_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_40_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_40_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_40_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_41 (
    .io_push_valid   (fifoGroup_41_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_41_io_push_ready        ), //o
    .io_push_payload (fifoGroup_41_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_41_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_41_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_41_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_41_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_41_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_42 (
    .io_push_valid   (fifoGroup_42_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_42_io_push_ready        ), //o
    .io_push_payload (fifoGroup_42_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_42_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_42_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_42_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_42_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_42_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_43 (
    .io_push_valid   (fifoGroup_43_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_43_io_push_ready        ), //o
    .io_push_payload (fifoGroup_43_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_43_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_43_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_43_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_43_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_43_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_44 (
    .io_push_valid   (fifoGroup_44_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_44_io_push_ready        ), //o
    .io_push_payload (fifoGroup_44_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_44_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_44_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_44_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_44_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_44_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_45 (
    .io_push_valid   (fifoGroup_45_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_45_io_push_ready        ), //o
    .io_push_payload (fifoGroup_45_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_45_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_45_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_45_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_45_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_45_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_46 (
    .io_push_valid   (fifoGroup_46_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_46_io_push_ready        ), //o
    .io_push_payload (fifoGroup_46_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_46_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_46_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_46_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_46_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_46_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_47 (
    .io_push_valid   (fifoGroup_47_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_47_io_push_ready        ), //o
    .io_push_payload (fifoGroup_47_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_47_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_47_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_47_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_47_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_47_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_48 (
    .io_push_valid   (fifoGroup_48_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_48_io_push_ready        ), //o
    .io_push_payload (fifoGroup_48_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_48_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_48_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_48_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_48_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_48_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_49 (
    .io_push_valid   (fifoGroup_49_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_49_io_push_ready        ), //o
    .io_push_payload (fifoGroup_49_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_49_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_49_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_49_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_49_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_49_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_50 (
    .io_push_valid   (fifoGroup_50_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_50_io_push_ready        ), //o
    .io_push_payload (fifoGroup_50_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_50_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_50_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_50_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_50_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_50_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_51 (
    .io_push_valid   (fifoGroup_51_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_51_io_push_ready        ), //o
    .io_push_payload (fifoGroup_51_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_51_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_51_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_51_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_51_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_51_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_52 (
    .io_push_valid   (fifoGroup_52_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_52_io_push_ready        ), //o
    .io_push_payload (fifoGroup_52_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_52_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_52_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_52_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_52_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_52_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_53 (
    .io_push_valid   (fifoGroup_53_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_53_io_push_ready        ), //o
    .io_push_payload (fifoGroup_53_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_53_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_53_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_53_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_53_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_53_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_54 (
    .io_push_valid   (fifoGroup_54_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_54_io_push_ready        ), //o
    .io_push_payload (fifoGroup_54_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_54_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_54_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_54_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_54_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_54_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_55 (
    .io_push_valid   (fifoGroup_55_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_55_io_push_ready        ), //o
    .io_push_payload (fifoGroup_55_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_55_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_55_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_55_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_55_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_55_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_56 (
    .io_push_valid   (fifoGroup_56_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_56_io_push_ready        ), //o
    .io_push_payload (fifoGroup_56_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_56_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_56_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_56_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_56_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_56_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_57 (
    .io_push_valid   (fifoGroup_57_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_57_io_push_ready        ), //o
    .io_push_payload (fifoGroup_57_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_57_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_57_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_57_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_57_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_57_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_58 (
    .io_push_valid   (fifoGroup_58_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_58_io_push_ready        ), //o
    .io_push_payload (fifoGroup_58_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_58_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_58_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_58_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_58_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_58_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_59 (
    .io_push_valid   (fifoGroup_59_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_59_io_push_ready        ), //o
    .io_push_payload (fifoGroup_59_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_59_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_59_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_59_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_59_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_59_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_60 (
    .io_push_valid   (fifoGroup_60_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_60_io_push_ready        ), //o
    .io_push_payload (fifoGroup_60_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_60_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_60_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_60_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_60_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_60_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_61 (
    .io_push_valid   (fifoGroup_61_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_61_io_push_ready        ), //o
    .io_push_payload (fifoGroup_61_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_61_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_61_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_61_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_61_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_61_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_62 (
    .io_push_valid   (fifoGroup_62_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_62_io_push_ready        ), //o
    .io_push_payload (fifoGroup_62_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_62_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_62_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_62_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_62_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_62_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_63 (
    .io_push_valid   (fifoGroup_63_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_63_io_push_ready        ), //o
    .io_push_payload (fifoGroup_63_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_63_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_63_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_63_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_63_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_63_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_64 (
    .io_push_valid   (fifoGroup_64_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_64_io_push_ready        ), //o
    .io_push_payload (fifoGroup_64_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_64_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_64_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_64_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_64_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_64_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_65 (
    .io_push_valid   (fifoGroup_65_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_65_io_push_ready        ), //o
    .io_push_payload (fifoGroup_65_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_65_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_65_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_65_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_65_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_65_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_66 (
    .io_push_valid   (fifoGroup_66_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_66_io_push_ready        ), //o
    .io_push_payload (fifoGroup_66_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_66_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_66_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_66_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_66_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_66_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_67 (
    .io_push_valid   (fifoGroup_67_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_67_io_push_ready        ), //o
    .io_push_payload (fifoGroup_67_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_67_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_67_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_67_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_67_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_67_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_68 (
    .io_push_valid   (fifoGroup_68_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_68_io_push_ready        ), //o
    .io_push_payload (fifoGroup_68_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_68_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_68_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_68_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_68_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_68_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_69 (
    .io_push_valid   (fifoGroup_69_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_69_io_push_ready        ), //o
    .io_push_payload (fifoGroup_69_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_69_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_69_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_69_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_69_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_69_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_70 (
    .io_push_valid   (fifoGroup_70_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_70_io_push_ready        ), //o
    .io_push_payload (fifoGroup_70_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_70_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_70_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_70_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_70_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_70_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_71 (
    .io_push_valid   (fifoGroup_71_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_71_io_push_ready        ), //o
    .io_push_payload (fifoGroup_71_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_71_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_71_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_71_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_71_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_71_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_72 (
    .io_push_valid   (fifoGroup_72_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_72_io_push_ready        ), //o
    .io_push_payload (fifoGroup_72_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_72_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_72_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_72_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_72_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_72_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_73 (
    .io_push_valid   (fifoGroup_73_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_73_io_push_ready        ), //o
    .io_push_payload (fifoGroup_73_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_73_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_73_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_73_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_73_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_73_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_74 (
    .io_push_valid   (fifoGroup_74_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_74_io_push_ready        ), //o
    .io_push_payload (fifoGroup_74_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_74_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_74_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_74_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_74_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_74_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_75 (
    .io_push_valid   (fifoGroup_75_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_75_io_push_ready        ), //o
    .io_push_payload (fifoGroup_75_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_75_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_75_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_75_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_75_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_75_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_76 (
    .io_push_valid   (fifoGroup_76_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_76_io_push_ready        ), //o
    .io_push_payload (fifoGroup_76_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_76_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_76_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_76_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_76_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_76_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_77 (
    .io_push_valid   (fifoGroup_77_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_77_io_push_ready        ), //o
    .io_push_payload (fifoGroup_77_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_77_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_77_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_77_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_77_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_77_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_78 (
    .io_push_valid   (fifoGroup_78_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_78_io_push_ready        ), //o
    .io_push_payload (fifoGroup_78_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_78_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_78_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_78_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_78_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_78_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_79 (
    .io_push_valid   (fifoGroup_79_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_79_io_push_ready        ), //o
    .io_push_payload (fifoGroup_79_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_79_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_79_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_79_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_79_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_79_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_80 (
    .io_push_valid   (fifoGroup_80_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_80_io_push_ready        ), //o
    .io_push_payload (fifoGroup_80_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_80_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_80_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_80_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_80_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_80_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_81 (
    .io_push_valid   (fifoGroup_81_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_81_io_push_ready        ), //o
    .io_push_payload (fifoGroup_81_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_81_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_81_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_81_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_81_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_81_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_82 (
    .io_push_valid   (fifoGroup_82_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_82_io_push_ready        ), //o
    .io_push_payload (fifoGroup_82_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_82_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_82_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_82_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_82_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_82_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_83 (
    .io_push_valid   (fifoGroup_83_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_83_io_push_ready        ), //o
    .io_push_payload (fifoGroup_83_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_83_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_83_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_83_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_83_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_83_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_84 (
    .io_push_valid   (fifoGroup_84_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_84_io_push_ready        ), //o
    .io_push_payload (fifoGroup_84_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_84_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_84_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_84_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_84_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_84_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_85 (
    .io_push_valid   (fifoGroup_85_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_85_io_push_ready        ), //o
    .io_push_payload (fifoGroup_85_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_85_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_85_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_85_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_85_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_85_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_86 (
    .io_push_valid   (fifoGroup_86_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_86_io_push_ready        ), //o
    .io_push_payload (fifoGroup_86_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_86_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_86_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_86_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_86_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_86_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_87 (
    .io_push_valid   (fifoGroup_87_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_87_io_push_ready        ), //o
    .io_push_payload (fifoGroup_87_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_87_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_87_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_87_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_87_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_87_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_88 (
    .io_push_valid   (fifoGroup_88_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_88_io_push_ready        ), //o
    .io_push_payload (fifoGroup_88_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_88_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_88_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_88_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_88_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_88_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_89 (
    .io_push_valid   (fifoGroup_89_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_89_io_push_ready        ), //o
    .io_push_payload (fifoGroup_89_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_89_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_89_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_89_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_89_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_89_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_90 (
    .io_push_valid   (fifoGroup_90_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_90_io_push_ready        ), //o
    .io_push_payload (fifoGroup_90_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_90_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_90_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_90_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_90_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_90_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_91 (
    .io_push_valid   (fifoGroup_91_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_91_io_push_ready        ), //o
    .io_push_payload (fifoGroup_91_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_91_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_91_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_91_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_91_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_91_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_92 (
    .io_push_valid   (fifoGroup_92_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_92_io_push_ready        ), //o
    .io_push_payload (fifoGroup_92_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_92_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_92_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_92_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_92_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_92_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_93 (
    .io_push_valid   (fifoGroup_93_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_93_io_push_ready        ), //o
    .io_push_payload (fifoGroup_93_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_93_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_93_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_93_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_93_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_93_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_94 (
    .io_push_valid   (fifoGroup_94_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_94_io_push_ready        ), //o
    .io_push_payload (fifoGroup_94_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_94_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_94_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_94_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_94_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_94_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_95 (
    .io_push_valid   (fifoGroup_95_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_95_io_push_ready        ), //o
    .io_push_payload (fifoGroup_95_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_95_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_95_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_95_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_95_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_95_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_96 (
    .io_push_valid   (fifoGroup_96_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_96_io_push_ready        ), //o
    .io_push_payload (fifoGroup_96_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_96_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_96_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_96_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_96_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_96_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_97 (
    .io_push_valid   (fifoGroup_97_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_97_io_push_ready        ), //o
    .io_push_payload (fifoGroup_97_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_97_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_97_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_97_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_97_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_97_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_98 (
    .io_push_valid   (fifoGroup_98_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_98_io_push_ready        ), //o
    .io_push_payload (fifoGroup_98_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_98_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_98_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_98_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_98_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_98_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_99 (
    .io_push_valid   (fifoGroup_99_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_99_io_push_ready        ), //o
    .io_push_payload (fifoGroup_99_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_99_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_99_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_99_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                              ), //i
    .io_occupancy    (fifoGroup_99_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_99_io_availability[6:0] ), //o
    .clk             (clk                               ), //i
    .resetn          (resetn                            )  //i
  );
  StreamFifo fifoGroup_100 (
    .io_push_valid   (fifoGroup_100_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_100_io_push_ready        ), //o
    .io_push_payload (fifoGroup_100_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_100_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_100_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_100_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_100_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_100_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_101 (
    .io_push_valid   (fifoGroup_101_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_101_io_push_ready        ), //o
    .io_push_payload (fifoGroup_101_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_101_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_101_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_101_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_101_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_101_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_102 (
    .io_push_valid   (fifoGroup_102_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_102_io_push_ready        ), //o
    .io_push_payload (fifoGroup_102_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_102_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_102_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_102_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_102_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_102_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_103 (
    .io_push_valid   (fifoGroup_103_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_103_io_push_ready        ), //o
    .io_push_payload (fifoGroup_103_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_103_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_103_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_103_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_103_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_103_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_104 (
    .io_push_valid   (fifoGroup_104_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_104_io_push_ready        ), //o
    .io_push_payload (fifoGroup_104_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_104_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_104_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_104_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_104_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_104_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_105 (
    .io_push_valid   (fifoGroup_105_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_105_io_push_ready        ), //o
    .io_push_payload (fifoGroup_105_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_105_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_105_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_105_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_105_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_105_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_106 (
    .io_push_valid   (fifoGroup_106_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_106_io_push_ready        ), //o
    .io_push_payload (fifoGroup_106_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_106_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_106_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_106_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_106_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_106_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_107 (
    .io_push_valid   (fifoGroup_107_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_107_io_push_ready        ), //o
    .io_push_payload (fifoGroup_107_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_107_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_107_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_107_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_107_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_107_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_108 (
    .io_push_valid   (fifoGroup_108_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_108_io_push_ready        ), //o
    .io_push_payload (fifoGroup_108_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_108_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_108_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_108_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_108_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_108_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo fifoGroup_109 (
    .io_push_valid   (fifoGroup_109_io_push_valid        ), //i
    .io_push_ready   (fifoGroup_109_io_push_ready        ), //o
    .io_push_payload (fifoGroup_109_io_push_payload[31:0]), //i
    .io_pop_valid    (fifoGroup_109_io_pop_valid         ), //o
    .io_pop_ready    (fifoGroup_109_io_pop_ready         ), //i
    .io_pop_payload  (fifoGroup_109_io_pop_payload[31:0] ), //o
    .io_flush        (1'b0                               ), //i
    .io_occupancy    (fifoGroup_109_io_occupancy[6:0]    ), //o
    .io_availability (fifoGroup_109_io_availability[6:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  always @(*) begin
    case(selectWriteFifo)
      7'b0000000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_0_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_0_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_0_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_0_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_0_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_0_io_occupancy;
      end
      7'b0000001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_1_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_1_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_1_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_1_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_1_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_1_io_occupancy;
      end
      7'b0000010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_2_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_2_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_2_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_2_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_2_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_2_io_occupancy;
      end
      7'b0000011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_3_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_3_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_3_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_3_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_3_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_3_io_occupancy;
      end
      7'b0000100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_4_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_4_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_4_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_4_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_4_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_4_io_occupancy;
      end
      7'b0000101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_5_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_5_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_5_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_5_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_5_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_5_io_occupancy;
      end
      7'b0000110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_6_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_6_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_6_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_6_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_6_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_6_io_occupancy;
      end
      7'b0000111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_7_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_7_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_7_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_7_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_7_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_7_io_occupancy;
      end
      7'b0001000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_8_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_8_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_8_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_8_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_8_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_8_io_occupancy;
      end
      7'b0001001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_9_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_9_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_9_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_9_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_9_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_9_io_occupancy;
      end
      7'b0001010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_10_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_10_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_10_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_10_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_10_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_10_io_occupancy;
      end
      7'b0001011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_11_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_11_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_11_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_11_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_11_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_11_io_occupancy;
      end
      7'b0001100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_12_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_12_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_12_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_12_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_12_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_12_io_occupancy;
      end
      7'b0001101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_13_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_13_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_13_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_13_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_13_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_13_io_occupancy;
      end
      7'b0001110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_14_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_14_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_14_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_14_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_14_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_14_io_occupancy;
      end
      7'b0001111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_15_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_15_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_15_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_15_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_15_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_15_io_occupancy;
      end
      7'b0010000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_16_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_16_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_16_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_16_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_16_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_16_io_occupancy;
      end
      7'b0010001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_17_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_17_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_17_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_17_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_17_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_17_io_occupancy;
      end
      7'b0010010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_18_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_18_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_18_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_18_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_18_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_18_io_occupancy;
      end
      7'b0010011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_19_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_19_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_19_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_19_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_19_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_19_io_occupancy;
      end
      7'b0010100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_20_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_20_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_20_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_20_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_20_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_20_io_occupancy;
      end
      7'b0010101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_21_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_21_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_21_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_21_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_21_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_21_io_occupancy;
      end
      7'b0010110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_22_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_22_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_22_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_22_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_22_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_22_io_occupancy;
      end
      7'b0010111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_23_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_23_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_23_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_23_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_23_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_23_io_occupancy;
      end
      7'b0011000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_24_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_24_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_24_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_24_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_24_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_24_io_occupancy;
      end
      7'b0011001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_25_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_25_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_25_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_25_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_25_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_25_io_occupancy;
      end
      7'b0011010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_26_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_26_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_26_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_26_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_26_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_26_io_occupancy;
      end
      7'b0011011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_27_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_27_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_27_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_27_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_27_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_27_io_occupancy;
      end
      7'b0011100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_28_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_28_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_28_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_28_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_28_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_28_io_occupancy;
      end
      7'b0011101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_29_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_29_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_29_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_29_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_29_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_29_io_occupancy;
      end
      7'b0011110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_30_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_30_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_30_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_30_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_30_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_30_io_occupancy;
      end
      7'b0011111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_31_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_31_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_31_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_31_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_31_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_31_io_occupancy;
      end
      7'b0100000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_32_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_32_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_32_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_32_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_32_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_32_io_occupancy;
      end
      7'b0100001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_33_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_33_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_33_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_33_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_33_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_33_io_occupancy;
      end
      7'b0100010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_34_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_34_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_34_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_34_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_34_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_34_io_occupancy;
      end
      7'b0100011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_35_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_35_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_35_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_35_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_35_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_35_io_occupancy;
      end
      7'b0100100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_36_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_36_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_36_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_36_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_36_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_36_io_occupancy;
      end
      7'b0100101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_37_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_37_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_37_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_37_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_37_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_37_io_occupancy;
      end
      7'b0100110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_38_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_38_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_38_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_38_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_38_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_38_io_occupancy;
      end
      7'b0100111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_39_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_39_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_39_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_39_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_39_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_39_io_occupancy;
      end
      7'b0101000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_40_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_40_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_40_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_40_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_40_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_40_io_occupancy;
      end
      7'b0101001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_41_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_41_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_41_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_41_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_41_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_41_io_occupancy;
      end
      7'b0101010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_42_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_42_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_42_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_42_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_42_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_42_io_occupancy;
      end
      7'b0101011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_43_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_43_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_43_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_43_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_43_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_43_io_occupancy;
      end
      7'b0101100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_44_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_44_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_44_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_44_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_44_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_44_io_occupancy;
      end
      7'b0101101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_45_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_45_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_45_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_45_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_45_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_45_io_occupancy;
      end
      7'b0101110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_46_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_46_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_46_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_46_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_46_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_46_io_occupancy;
      end
      7'b0101111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_47_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_47_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_47_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_47_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_47_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_47_io_occupancy;
      end
      7'b0110000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_48_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_48_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_48_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_48_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_48_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_48_io_occupancy;
      end
      7'b0110001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_49_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_49_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_49_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_49_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_49_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_49_io_occupancy;
      end
      7'b0110010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_50_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_50_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_50_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_50_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_50_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_50_io_occupancy;
      end
      7'b0110011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_51_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_51_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_51_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_51_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_51_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_51_io_occupancy;
      end
      7'b0110100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_52_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_52_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_52_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_52_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_52_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_52_io_occupancy;
      end
      7'b0110101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_53_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_53_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_53_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_53_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_53_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_53_io_occupancy;
      end
      7'b0110110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_54_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_54_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_54_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_54_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_54_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_54_io_occupancy;
      end
      7'b0110111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_55_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_55_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_55_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_55_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_55_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_55_io_occupancy;
      end
      7'b0111000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_56_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_56_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_56_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_56_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_56_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_56_io_occupancy;
      end
      7'b0111001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_57_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_57_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_57_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_57_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_57_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_57_io_occupancy;
      end
      7'b0111010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_58_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_58_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_58_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_58_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_58_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_58_io_occupancy;
      end
      7'b0111011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_59_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_59_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_59_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_59_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_59_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_59_io_occupancy;
      end
      7'b0111100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_60_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_60_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_60_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_60_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_60_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_60_io_occupancy;
      end
      7'b0111101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_61_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_61_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_61_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_61_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_61_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_61_io_occupancy;
      end
      7'b0111110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_62_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_62_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_62_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_62_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_62_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_62_io_occupancy;
      end
      7'b0111111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_63_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_63_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_63_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_63_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_63_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_63_io_occupancy;
      end
      7'b1000000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_64_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_64_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_64_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_64_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_64_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_64_io_occupancy;
      end
      7'b1000001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_65_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_65_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_65_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_65_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_65_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_65_io_occupancy;
      end
      7'b1000010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_66_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_66_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_66_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_66_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_66_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_66_io_occupancy;
      end
      7'b1000011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_67_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_67_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_67_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_67_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_67_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_67_io_occupancy;
      end
      7'b1000100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_68_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_68_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_68_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_68_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_68_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_68_io_occupancy;
      end
      7'b1000101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_69_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_69_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_69_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_69_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_69_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_69_io_occupancy;
      end
      7'b1000110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_70_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_70_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_70_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_70_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_70_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_70_io_occupancy;
      end
      7'b1000111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_71_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_71_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_71_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_71_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_71_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_71_io_occupancy;
      end
      7'b1001000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_72_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_72_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_72_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_72_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_72_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_72_io_occupancy;
      end
      7'b1001001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_73_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_73_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_73_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_73_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_73_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_73_io_occupancy;
      end
      7'b1001010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_74_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_74_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_74_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_74_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_74_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_74_io_occupancy;
      end
      7'b1001011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_75_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_75_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_75_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_75_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_75_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_75_io_occupancy;
      end
      7'b1001100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_76_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_76_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_76_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_76_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_76_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_76_io_occupancy;
      end
      7'b1001101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_77_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_77_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_77_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_77_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_77_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_77_io_occupancy;
      end
      7'b1001110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_78_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_78_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_78_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_78_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_78_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_78_io_occupancy;
      end
      7'b1001111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_79_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_79_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_79_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_79_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_79_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_79_io_occupancy;
      end
      7'b1010000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_80_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_80_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_80_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_80_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_80_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_80_io_occupancy;
      end
      7'b1010001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_81_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_81_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_81_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_81_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_81_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_81_io_occupancy;
      end
      7'b1010010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_82_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_82_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_82_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_82_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_82_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_82_io_occupancy;
      end
      7'b1010011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_83_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_83_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_83_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_83_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_83_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_83_io_occupancy;
      end
      7'b1010100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_84_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_84_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_84_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_84_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_84_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_84_io_occupancy;
      end
      7'b1010101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_85_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_85_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_85_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_85_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_85_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_85_io_occupancy;
      end
      7'b1010110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_86_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_86_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_86_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_86_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_86_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_86_io_occupancy;
      end
      7'b1010111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_87_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_87_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_87_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_87_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_87_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_87_io_occupancy;
      end
      7'b1011000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_88_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_88_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_88_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_88_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_88_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_88_io_occupancy;
      end
      7'b1011001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_89_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_89_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_89_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_89_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_89_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_89_io_occupancy;
      end
      7'b1011010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_90_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_90_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_90_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_90_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_90_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_90_io_occupancy;
      end
      7'b1011011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_91_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_91_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_91_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_91_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_91_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_91_io_occupancy;
      end
      7'b1011100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_92_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_92_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_92_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_92_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_92_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_92_io_occupancy;
      end
      7'b1011101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_93_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_93_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_93_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_93_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_93_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_93_io_occupancy;
      end
      7'b1011110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_94_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_94_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_94_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_94_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_94_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_94_io_occupancy;
      end
      7'b1011111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_95_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_95_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_95_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_95_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_95_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_95_io_occupancy;
      end
      7'b1100000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_96_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_96_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_96_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_96_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_96_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_96_io_occupancy;
      end
      7'b1100001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_97_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_97_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_97_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_97_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_97_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_97_io_occupancy;
      end
      7'b1100010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_98_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_98_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_98_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_98_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_98_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_98_io_occupancy;
      end
      7'b1100011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_99_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_99_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_99_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_99_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_99_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_99_io_occupancy;
      end
      7'b1100100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_100_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_100_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_100_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_100_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_100_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_100_io_occupancy;
      end
      7'b1100101 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_101_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_101_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_101_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_101_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_101_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_101_io_occupancy;
      end
      7'b1100110 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_102_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_102_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_102_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_102_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_102_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_102_io_occupancy;
      end
      7'b1100111 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_103_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_103_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_103_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_103_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_103_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_103_io_occupancy;
      end
      7'b1101000 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_104_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_104_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_104_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_104_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_104_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_104_io_occupancy;
      end
      7'b1101001 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_105_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_105_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_105_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_105_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_105_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_105_io_occupancy;
      end
      7'b1101010 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_106_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_106_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_106_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_106_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_106_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_106_io_occupancy;
      end
      7'b1101011 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_107_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_107_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_107_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_107_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_107_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_107_io_occupancy;
      end
      7'b1101100 : begin
        _zz_when_ArraySlice_l204 = fifoGroup_108_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_108_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_108_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_108_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_108_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_108_io_occupancy;
      end
      default : begin
        _zz_when_ArraySlice_l204 = fifoGroup_109_io_occupancy;
        _zz_inputStreamArrayData_ready = fifoGroup_109_io_push_ready;
        _zz_when_ArraySlice_l208 = fifoGroup_109_io_occupancy;
        _zz_when_ArraySlice_l337 = fifoGroup_109_io_occupancy;
        _zz_inputStreamArrayData_ready_1 = fifoGroup_109_io_push_ready;
        _zz_when_ArraySlice_l341 = fifoGroup_109_io_occupancy;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_1)
      7'b0000000 : _zz_when_ArraySlice_l377 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_0_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_0_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_0_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_0_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_0_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_0_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_0_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_0_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_0_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_0_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_0_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_0_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_0_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_0_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_0_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_0_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_0_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_0_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_0_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_0_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_0_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_0_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_0_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_0_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_0_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_0_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_0_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_0_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_0_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_0_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_0_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_0_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_0_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_0_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_0_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_0_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_0_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_0_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_0_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_0_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_0_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_0_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_0_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_0_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_0_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_0_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_0_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_0_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_0_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_0_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_0_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_0_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_0_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_0_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_0_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_0_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_0_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_0_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_0_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_0_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_0_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_0_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_0_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_0_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_0_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_0_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_0_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_0_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_0_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_0_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_0_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_0_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_0_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_0_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_0_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_0_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_0_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_0_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_0_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_0_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_0_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_0_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_0_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_0_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_0_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_0_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_0_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_0_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_0_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_0_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_0_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_0_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_0_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_0_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_0_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_0_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_0_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_0_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_0_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_0_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_0_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_0_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_0_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_0_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_0_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_0_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_0_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_0_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_0_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_0_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_0_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_1)
      7'b0000000 : _zz_when_ArraySlice_l383 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_1)
      7'b0000000 : _zz_when_ArraySlice_l392 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_1)
      7'b0000000 : _zz_when_ArraySlice_l417 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_1_2)
      7'b0000000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_1_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_1_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_1_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_1_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_1_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_1_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_1_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_1_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_1_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_1_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_1_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_1_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_1_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_1_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_1_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_1_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_1_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_1_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_1_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_1_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_1_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_1_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_1_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_1_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_1_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_1_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_1_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_1_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_1_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_1_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_1_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_1_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_1_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_1_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_1_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_1_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_1_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_1_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_1_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_1_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_1_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_1_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_1_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_1_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_1_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_1_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_1_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_1_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_1_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_1_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_1_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_1_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_1_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_1_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_1_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_1_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_1_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_1_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_1_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_1_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_1_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_1_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_1_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_1_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_1_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_1_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_1_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_1_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_1_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_1_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_1_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_1_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_1_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_1_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_1_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_1_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_1_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_1_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_1_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_1_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_1_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_1_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_1_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_1_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_1_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_1_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_1_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_1_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_1_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_1_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_1_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_1_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_1_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_1_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_1_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_1_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_1_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_1_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_1_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_1_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_1_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_1_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_1_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_1_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_1_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_1_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_1_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_1_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_1_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_1_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_1_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_1_2)
      7'b0000000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_1_2)
      7'b0000000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_1_2)
      7'b0000000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_2_2)
      7'b0000000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_2_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_2_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_2_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_2_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_2_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_2_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_2_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_2_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_2_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_2_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_2_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_2_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_2_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_2_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_2_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_2_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_2_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_2_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_2_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_2_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_2_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_2_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_2_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_2_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_2_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_2_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_2_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_2_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_2_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_2_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_2_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_2_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_2_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_2_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_2_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_2_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_2_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_2_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_2_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_2_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_2_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_2_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_2_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_2_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_2_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_2_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_2_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_2_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_2_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_2_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_2_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_2_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_2_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_2_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_2_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_2_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_2_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_2_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_2_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_2_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_2_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_2_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_2_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_2_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_2_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_2_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_2_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_2_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_2_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_2_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_2_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_2_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_2_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_2_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_2_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_2_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_2_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_2_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_2_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_2_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_2_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_2_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_2_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_2_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_2_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_2_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_2_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_2_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_2_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_2_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_2_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_2_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_2_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_2_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_2_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_2_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_2_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_2_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_2_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_2_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_2_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_2_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_2_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_2_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_2_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_2_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_2_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_2_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_2_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_2_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_2_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_2_2)
      7'b0000000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_2_2)
      7'b0000000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_2_2)
      7'b0000000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_3_2)
      7'b0000000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_3_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_3_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_3_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_3_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_3_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_3_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_3_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_3_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_3_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_3_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_3_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_3_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_3_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_3_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_3_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_3_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_3_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_3_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_3_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_3_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_3_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_3_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_3_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_3_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_3_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_3_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_3_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_3_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_3_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_3_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_3_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_3_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_3_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_3_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_3_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_3_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_3_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_3_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_3_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_3_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_3_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_3_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_3_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_3_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_3_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_3_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_3_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_3_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_3_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_3_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_3_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_3_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_3_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_3_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_3_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_3_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_3_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_3_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_3_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_3_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_3_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_3_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_3_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_3_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_3_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_3_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_3_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_3_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_3_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_3_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_3_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_3_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_3_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_3_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_3_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_3_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_3_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_3_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_3_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_3_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_3_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_3_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_3_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_3_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_3_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_3_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_3_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_3_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_3_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_3_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_3_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_3_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_3_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_3_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_3_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_3_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_3_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_3_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_3_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_3_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_3_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_3_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_3_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_3_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_3_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_3_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_3_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_3_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_3_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_3_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_3_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_3_2)
      7'b0000000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_3_2)
      7'b0000000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_3_2)
      7'b0000000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_4_2)
      7'b0000000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_4_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_4_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_4_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_4_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_4_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_4_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_4_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_4_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_4_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_4_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_4_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_4_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_4_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_4_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_4_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_4_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_4_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_4_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_4_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_4_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_4_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_4_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_4_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_4_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_4_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_4_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_4_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_4_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_4_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_4_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_4_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_4_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_4_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_4_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_4_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_4_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_4_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_4_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_4_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_4_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_4_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_4_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_4_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_4_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_4_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_4_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_4_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_4_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_4_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_4_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_4_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_4_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_4_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_4_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_4_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_4_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_4_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_4_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_4_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_4_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_4_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_4_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_4_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_4_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_4_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_4_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_4_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_4_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_4_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_4_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_4_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_4_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_4_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_4_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_4_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_4_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_4_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_4_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_4_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_4_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_4_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_4_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_4_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_4_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_4_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_4_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_4_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_4_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_4_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_4_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_4_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_4_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_4_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_4_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_4_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_4_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_4_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_4_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_4_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_4_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_4_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_4_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_4_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_4_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_4_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_4_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_4_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_4_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_4_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_4_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_4_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_4_2)
      7'b0000000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_4_2)
      7'b0000000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_4_2)
      7'b0000000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_5_1)
      7'b0000000 : _zz_when_ArraySlice_l377_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_5_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_5_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_5_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_5_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_5_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_5_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_5_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_5_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_5_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_5_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_5_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_5_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_5_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_5_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_5_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_5_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_5_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_5_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_5_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_5_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_5_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_5_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_5_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_5_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_5_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_5_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_5_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_5_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_5_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_5_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_5_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_5_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_5_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_5_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_5_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_5_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_5_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_5_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_5_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_5_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_5_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_5_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_5_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_5_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_5_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_5_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_5_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_5_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_5_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_5_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_5_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_5_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_5_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_5_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_5_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_5_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_5_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_5_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_5_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_5_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_5_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_5_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_5_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_5_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_5_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_5_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_5_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_5_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_5_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_5_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_5_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_5_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_5_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_5_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_5_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_5_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_5_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_5_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_5_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_5_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_5_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_5_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_5_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_5_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_5_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_5_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_5_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_5_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_5_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_5_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_5_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_5_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_5_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_5_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_5_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_5_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_5_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_5_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_5_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_5_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_5_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_5_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_5_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_5_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_5_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_5_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_5_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_5_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_5_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_5_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_5_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_5_1)
      7'b0000000 : _zz_when_ArraySlice_l383_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_5_1)
      7'b0000000 : _zz_when_ArraySlice_l392_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_5_1)
      7'b0000000 : _zz_when_ArraySlice_l417_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_6_1)
      7'b0000000 : _zz_when_ArraySlice_l377_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_6_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_6_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_6_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_6_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_6_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_6_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_6_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_6_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_6_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_6_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_6_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_6_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_6_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_6_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_6_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_6_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_6_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_6_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_6_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_6_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_6_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_6_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_6_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_6_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_6_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_6_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_6_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_6_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_6_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_6_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_6_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_6_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_6_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_6_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_6_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_6_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_6_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_6_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_6_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_6_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_6_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_6_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_6_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_6_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_6_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_6_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_6_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_6_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_6_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_6_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_6_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_6_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_6_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_6_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_6_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_6_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_6_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_6_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_6_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_6_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_6_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_6_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_6_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_6_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_6_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_6_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_6_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_6_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_6_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_6_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_6_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_6_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_6_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_6_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_6_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_6_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_6_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_6_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_6_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_6_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_6_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_6_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_6_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_6_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_6_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_6_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_6_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_6_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_6_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_6_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_6_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_6_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_6_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_6_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_6_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_6_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_6_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_6_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_6_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_6_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_6_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_6_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_6_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_6_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_6_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_6_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_6_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_6_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_6_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_6_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_6_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_6_1)
      7'b0000000 : _zz_when_ArraySlice_l383_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_6_1)
      7'b0000000 : _zz_when_ArraySlice_l392_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_6_1)
      7'b0000000 : _zz_when_ArraySlice_l417_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l377_7_1)
      7'b0000000 : _zz_when_ArraySlice_l377_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l377_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l377_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l377_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l377_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l377_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l377_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l377_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l377_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l377_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l377_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l377_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l377_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l377_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l377_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l377_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l377_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l377_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l377_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l377_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l377_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l377_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l377_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l377_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l377_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l377_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l377_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l377_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l377_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l377_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l377_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l377_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l377_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l377_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l377_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l377_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l377_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l377_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l377_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l377_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l377_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l377_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l377_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l377_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l377_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l377_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l377_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l377_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l377_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l377_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l377_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l377_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l377_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l377_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l377_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l377_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l377_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l377_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l377_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l377_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l377_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l377_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l377_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l377_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l377_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l377_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l377_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l377_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l377_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l377_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l377_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l377_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l377_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l377_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l377_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l377_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l377_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l377_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l377_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l377_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l377_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l377_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l377_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l377_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l377_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l377_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l377_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l377_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l377_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l377_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l377_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l377_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l377_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l377_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l377_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l377_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l377_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l377_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l377_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l377_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l377_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l377_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l377_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l377_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l377_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l377_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l377_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l377_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l377_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l377_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_valid_3)
      7'b0000000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_7_valid_2 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_payload_1)
      7'b0000000 : _zz_outputStreamArrayData_7_payload = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_7_payload = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_7_payload = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_7_payload = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_7_payload = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_7_payload = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_7_payload = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_7_payload = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_7_payload = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_7_payload = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_7_payload = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_7_payload = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_7_payload = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_7_payload = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_7_payload = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_7_payload = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_7_payload = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_7_payload = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_7_payload = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_7_payload = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_7_payload = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_7_payload = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_7_payload = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_7_payload = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_7_payload = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_7_payload = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_7_payload = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_7_payload = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_7_payload = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_7_payload = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_7_payload = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_7_payload = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_7_payload = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_7_payload = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_7_payload = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_7_payload = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_7_payload = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_7_payload = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_7_payload = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_7_payload = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_7_payload = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_7_payload = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_7_payload = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_7_payload = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_7_payload = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_7_payload = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_7_payload = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_7_payload = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_7_payload = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_7_payload = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_7_payload = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_7_payload = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_7_payload = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_7_payload = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_7_payload = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_7_payload = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_7_payload = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_7_payload = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_7_payload = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_7_payload = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_7_payload = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_7_payload = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_7_payload = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_7_payload = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_7_payload = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_7_payload = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_7_payload = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_7_payload = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_7_payload = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_7_payload = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_7_payload = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_7_payload = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_7_payload = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_7_payload = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_7_payload = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_7_payload = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_7_payload = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_7_payload = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_7_payload = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_7_payload = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_7_payload = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_7_payload = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_7_payload = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_7_payload = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_7_payload = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_7_payload = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_7_payload = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_7_payload = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_7_payload = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_7_payload = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_7_payload = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_7_payload = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_7_payload = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_7_payload = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_7_payload = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_7_payload = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_7_payload = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_7_payload = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_7_payload = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_7_payload = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_7_payload = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_7_payload = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_7_payload = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_7_payload = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_7_payload = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_7_payload = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_7_payload = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_7_payload = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_7_payload = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_7_payload = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l383_7_1)
      7'b0000000 : _zz_when_ArraySlice_l383_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l383_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l383_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l383_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l383_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l383_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l383_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l383_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l383_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l383_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l383_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l383_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l383_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l383_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l383_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l383_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l383_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l383_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l383_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l383_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l383_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l383_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l383_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l383_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l383_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l383_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l383_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l383_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l383_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l383_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l383_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l383_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l383_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l383_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l383_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l383_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l383_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l383_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l383_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l383_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l383_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l383_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l383_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l383_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l383_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l383_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l383_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l383_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l383_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l383_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l383_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l383_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l383_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l383_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l383_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l383_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l383_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l383_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l383_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l383_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l383_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l383_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l383_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l383_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l383_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l383_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l383_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l383_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l383_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l383_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l383_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l383_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l383_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l383_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l383_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l383_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l383_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l383_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l383_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l383_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l383_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l383_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l383_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l383_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l383_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l383_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l383_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l383_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l383_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l383_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l383_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l383_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l383_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l383_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l383_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l383_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l383_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l383_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l383_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l383_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l383_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l383_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l383_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l383_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l383_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l383_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l383_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l383_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l383_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l383_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l392_7_1)
      7'b0000000 : _zz_when_ArraySlice_l392_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l392_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l392_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l392_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l392_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l392_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l392_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l392_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l392_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l392_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l392_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l392_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l392_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l392_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l392_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l392_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l392_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l392_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l392_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l392_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l392_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l392_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l392_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l392_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l392_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l392_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l392_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l392_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l392_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l392_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l392_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l392_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l392_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l392_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l392_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l392_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l392_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l392_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l392_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l392_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l392_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l392_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l392_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l392_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l392_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l392_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l392_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l392_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l392_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l392_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l392_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l392_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l392_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l392_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l392_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l392_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l392_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l392_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l392_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l392_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l392_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l392_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l392_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l392_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l392_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l392_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l392_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l392_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l392_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l392_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l392_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l392_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l392_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l392_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l392_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l392_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l392_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l392_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l392_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l392_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l392_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l392_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l392_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l392_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l392_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l392_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l392_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l392_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l392_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l392_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l392_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l392_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l392_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l392_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l392_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l392_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l392_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l392_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l392_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l392_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l392_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l392_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l392_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l392_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l392_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l392_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l392_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l392_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l392_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l392_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l417_7_1)
      7'b0000000 : _zz_when_ArraySlice_l417_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l417_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l417_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l417_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l417_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l417_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l417_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l417_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l417_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l417_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l417_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l417_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l417_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l417_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l417_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l417_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l417_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l417_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l417_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l417_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l417_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l417_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l417_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l417_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l417_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l417_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l417_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l417_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l417_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l417_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l417_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l417_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l417_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l417_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l417_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l417_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l417_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l417_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l417_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l417_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l417_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l417_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l417_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l417_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l417_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l417_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l417_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l417_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l417_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l417_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l417_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l417_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l417_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l417_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l417_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l417_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l417_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l417_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l417_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l417_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l417_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l417_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l417_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l417_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l417_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l417_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l417_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l417_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l417_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l417_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l417_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l417_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l417_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l417_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l417_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l417_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l417_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l417_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l417_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l417_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l417_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l417_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l417_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l417_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l417_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l417_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l417_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l417_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l417_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l417_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l417_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l417_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l417_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l417_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l417_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l417_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l417_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l417_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l417_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l417_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l417_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l417_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l417_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l417_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l417_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l417_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l417_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l417_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l417_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l417_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_1)
      7'b0000000 : _zz_when_ArraySlice_l234 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_0_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_0_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_0_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_1)
      7'b0000000 : _zz_when_ArraySlice_l240 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_1)
      7'b0000000 : _zz_when_ArraySlice_l249 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_1)
      7'b0000000 : _zz_when_ArraySlice_l274 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_1_2)
      7'b0000000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_1_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_1_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_1_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_1_2)
      7'b0000000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_1_2)
      7'b0000000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_1_2)
      7'b0000000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_1_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_1_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_2_2)
      7'b0000000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_2_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_2_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_2_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_2_2)
      7'b0000000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_2_2)
      7'b0000000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_2_2)
      7'b0000000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_2_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_2_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_3_2)
      7'b0000000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_3_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_3_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_3_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_3_2)
      7'b0000000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_3_2)
      7'b0000000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_3_2)
      7'b0000000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_3_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_3_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_4_2)
      7'b0000000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_4_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_4_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_4_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_4_2)
      7'b0000000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_4_2)
      7'b0000000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_4_2)
      7'b0000000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_4_1 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_4_1 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_5_1)
      7'b0000000 : _zz_when_ArraySlice_l234_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_5_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_5_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_5_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_5_1)
      7'b0000000 : _zz_when_ArraySlice_l240_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_5_1)
      7'b0000000 : _zz_when_ArraySlice_l249_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_5_1)
      7'b0000000 : _zz_when_ArraySlice_l274_5 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_5 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_5 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_5 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_5 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_5 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_5 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_5 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_5 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_5 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_5 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_5 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_5 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_5 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_5 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_5 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_5 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_5 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_5 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_5 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_5 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_5 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_5 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_5 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_5 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_5 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_5 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_5 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_5 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_5 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_5 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_5 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_5 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_5 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_5 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_5 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_5 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_5 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_5 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_5 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_5 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_5 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_5 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_5 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_5 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_5 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_5 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_5 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_5 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_5 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_5 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_5 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_5 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_5 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_5 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_5 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_5 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_5 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_5 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_5 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_5 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_5 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_5 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_5 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_5 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_5 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_5 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_5 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_5 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_5 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_5 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_5 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_5 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_5 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_5 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_5 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_5 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_5 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_5 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_5 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_5 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_5 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_5 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_5 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_5 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_5 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_5 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_5 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_5 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_5 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_5 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_5 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_5 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_5 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_5 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_5 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_5 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_5 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_5 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_5 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_5 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_5 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_5 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_5 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_5 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_5 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_5 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_5 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_5 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_5 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_6_1)
      7'b0000000 : _zz_when_ArraySlice_l234_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_6_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_6_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_6_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_6_1)
      7'b0000000 : _zz_when_ArraySlice_l240_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_6_1)
      7'b0000000 : _zz_when_ArraySlice_l249_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_6_1)
      7'b0000000 : _zz_when_ArraySlice_l274_6 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_6 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_6 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_6 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_6 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_6 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_6 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_6 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_6 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_6 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_6 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_6 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_6 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_6 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_6 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_6 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_6 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_6 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_6 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_6 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_6 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_6 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_6 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_6 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_6 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_6 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_6 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_6 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_6 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_6 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_6 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_6 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_6 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_6 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_6 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_6 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_6 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_6 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_6 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_6 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_6 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_6 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_6 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_6 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_6 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_6 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_6 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_6 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_6 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_6 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_6 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_6 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_6 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_6 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_6 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_6 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_6 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_6 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_6 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_6 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_6 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_6 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_6 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_6 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_6 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_6 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_6 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_6 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_6 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_6 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_6 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_6 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_6 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_6 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_6 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_6 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_6 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_6 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_6 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_6 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_6 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_6 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_6 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_6 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_6 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_6 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_6 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_6 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_6 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_6 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_6 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_6 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_6 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_6 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_6 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_6 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_6 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_6 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_6 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_6 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_6 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_6 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_6 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_6 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_6 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_6 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_6 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_6 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_6 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_6 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l234_7_1)
      7'b0000000 : _zz_when_ArraySlice_l234_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l234_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l234_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l234_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l234_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l234_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l234_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l234_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l234_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l234_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l234_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l234_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l234_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l234_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l234_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l234_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l234_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l234_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l234_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l234_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l234_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l234_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l234_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l234_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l234_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l234_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l234_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l234_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l234_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l234_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l234_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l234_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l234_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l234_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l234_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l234_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l234_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l234_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l234_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l234_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l234_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l234_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l234_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l234_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l234_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l234_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l234_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l234_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l234_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l234_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l234_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l234_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l234_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l234_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l234_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l234_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l234_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l234_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l234_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l234_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l234_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l234_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l234_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l234_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l234_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l234_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l234_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l234_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l234_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l234_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l234_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l234_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l234_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l234_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l234_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l234_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l234_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l234_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l234_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l234_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l234_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l234_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l234_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l234_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l234_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l234_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l234_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l234_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l234_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l234_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l234_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l234_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l234_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l234_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l234_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l234_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l234_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l234_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l234_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l234_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l234_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l234_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l234_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l234_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l234_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l234_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l234_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l234_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l234_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l234_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_valid_5)
      7'b0000000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_0_io_pop_valid;
      7'b0000001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_1_io_pop_valid;
      7'b0000010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_2_io_pop_valid;
      7'b0000011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_3_io_pop_valid;
      7'b0000100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_4_io_pop_valid;
      7'b0000101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_5_io_pop_valid;
      7'b0000110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_6_io_pop_valid;
      7'b0000111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_7_io_pop_valid;
      7'b0001000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_8_io_pop_valid;
      7'b0001001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_9_io_pop_valid;
      7'b0001010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_10_io_pop_valid;
      7'b0001011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_11_io_pop_valid;
      7'b0001100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_12_io_pop_valid;
      7'b0001101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_13_io_pop_valid;
      7'b0001110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_14_io_pop_valid;
      7'b0001111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_15_io_pop_valid;
      7'b0010000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_16_io_pop_valid;
      7'b0010001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_17_io_pop_valid;
      7'b0010010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_18_io_pop_valid;
      7'b0010011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_19_io_pop_valid;
      7'b0010100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_20_io_pop_valid;
      7'b0010101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_21_io_pop_valid;
      7'b0010110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_22_io_pop_valid;
      7'b0010111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_23_io_pop_valid;
      7'b0011000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_24_io_pop_valid;
      7'b0011001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_25_io_pop_valid;
      7'b0011010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_26_io_pop_valid;
      7'b0011011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_27_io_pop_valid;
      7'b0011100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_28_io_pop_valid;
      7'b0011101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_29_io_pop_valid;
      7'b0011110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_30_io_pop_valid;
      7'b0011111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_31_io_pop_valid;
      7'b0100000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_32_io_pop_valid;
      7'b0100001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_33_io_pop_valid;
      7'b0100010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_34_io_pop_valid;
      7'b0100011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_35_io_pop_valid;
      7'b0100100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_36_io_pop_valid;
      7'b0100101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_37_io_pop_valid;
      7'b0100110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_38_io_pop_valid;
      7'b0100111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_39_io_pop_valid;
      7'b0101000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_40_io_pop_valid;
      7'b0101001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_41_io_pop_valid;
      7'b0101010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_42_io_pop_valid;
      7'b0101011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_43_io_pop_valid;
      7'b0101100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_44_io_pop_valid;
      7'b0101101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_45_io_pop_valid;
      7'b0101110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_46_io_pop_valid;
      7'b0101111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_47_io_pop_valid;
      7'b0110000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_48_io_pop_valid;
      7'b0110001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_49_io_pop_valid;
      7'b0110010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_50_io_pop_valid;
      7'b0110011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_51_io_pop_valid;
      7'b0110100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_52_io_pop_valid;
      7'b0110101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_53_io_pop_valid;
      7'b0110110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_54_io_pop_valid;
      7'b0110111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_55_io_pop_valid;
      7'b0111000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_56_io_pop_valid;
      7'b0111001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_57_io_pop_valid;
      7'b0111010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_58_io_pop_valid;
      7'b0111011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_59_io_pop_valid;
      7'b0111100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_60_io_pop_valid;
      7'b0111101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_61_io_pop_valid;
      7'b0111110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_62_io_pop_valid;
      7'b0111111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_63_io_pop_valid;
      7'b1000000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_64_io_pop_valid;
      7'b1000001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_65_io_pop_valid;
      7'b1000010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_66_io_pop_valid;
      7'b1000011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_67_io_pop_valid;
      7'b1000100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_68_io_pop_valid;
      7'b1000101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_69_io_pop_valid;
      7'b1000110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_70_io_pop_valid;
      7'b1000111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_71_io_pop_valid;
      7'b1001000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_72_io_pop_valid;
      7'b1001001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_73_io_pop_valid;
      7'b1001010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_74_io_pop_valid;
      7'b1001011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_75_io_pop_valid;
      7'b1001100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_76_io_pop_valid;
      7'b1001101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_77_io_pop_valid;
      7'b1001110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_78_io_pop_valid;
      7'b1001111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_79_io_pop_valid;
      7'b1010000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_80_io_pop_valid;
      7'b1010001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_81_io_pop_valid;
      7'b1010010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_82_io_pop_valid;
      7'b1010011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_83_io_pop_valid;
      7'b1010100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_84_io_pop_valid;
      7'b1010101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_85_io_pop_valid;
      7'b1010110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_86_io_pop_valid;
      7'b1010111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_87_io_pop_valid;
      7'b1011000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_88_io_pop_valid;
      7'b1011001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_89_io_pop_valid;
      7'b1011010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_90_io_pop_valid;
      7'b1011011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_91_io_pop_valid;
      7'b1011100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_92_io_pop_valid;
      7'b1011101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_93_io_pop_valid;
      7'b1011110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_94_io_pop_valid;
      7'b1011111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_95_io_pop_valid;
      7'b1100000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_96_io_pop_valid;
      7'b1100001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_97_io_pop_valid;
      7'b1100010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_98_io_pop_valid;
      7'b1100011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_99_io_pop_valid;
      7'b1100100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_100_io_pop_valid;
      7'b1100101 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_101_io_pop_valid;
      7'b1100110 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_102_io_pop_valid;
      7'b1100111 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_103_io_pop_valid;
      7'b1101000 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_104_io_pop_valid;
      7'b1101001 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_105_io_pop_valid;
      7'b1101010 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_106_io_pop_valid;
      7'b1101011 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_107_io_pop_valid;
      7'b1101100 : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_108_io_pop_valid;
      default : _zz_outputStreamArrayData_7_valid_4 = fifoGroup_109_io_pop_valid;
    endcase
  end

  always @(*) begin
    case(_zz_outputStreamArrayData_7_payload_3)
      7'b0000000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_0_io_pop_payload;
      7'b0000001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_1_io_pop_payload;
      7'b0000010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_2_io_pop_payload;
      7'b0000011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_3_io_pop_payload;
      7'b0000100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_4_io_pop_payload;
      7'b0000101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_5_io_pop_payload;
      7'b0000110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_6_io_pop_payload;
      7'b0000111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_7_io_pop_payload;
      7'b0001000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_8_io_pop_payload;
      7'b0001001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_9_io_pop_payload;
      7'b0001010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_10_io_pop_payload;
      7'b0001011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_11_io_pop_payload;
      7'b0001100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_12_io_pop_payload;
      7'b0001101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_13_io_pop_payload;
      7'b0001110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_14_io_pop_payload;
      7'b0001111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_15_io_pop_payload;
      7'b0010000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_16_io_pop_payload;
      7'b0010001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_17_io_pop_payload;
      7'b0010010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_18_io_pop_payload;
      7'b0010011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_19_io_pop_payload;
      7'b0010100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_20_io_pop_payload;
      7'b0010101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_21_io_pop_payload;
      7'b0010110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_22_io_pop_payload;
      7'b0010111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_23_io_pop_payload;
      7'b0011000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_24_io_pop_payload;
      7'b0011001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_25_io_pop_payload;
      7'b0011010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_26_io_pop_payload;
      7'b0011011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_27_io_pop_payload;
      7'b0011100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_28_io_pop_payload;
      7'b0011101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_29_io_pop_payload;
      7'b0011110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_30_io_pop_payload;
      7'b0011111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_31_io_pop_payload;
      7'b0100000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_32_io_pop_payload;
      7'b0100001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_33_io_pop_payload;
      7'b0100010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_34_io_pop_payload;
      7'b0100011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_35_io_pop_payload;
      7'b0100100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_36_io_pop_payload;
      7'b0100101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_37_io_pop_payload;
      7'b0100110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_38_io_pop_payload;
      7'b0100111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_39_io_pop_payload;
      7'b0101000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_40_io_pop_payload;
      7'b0101001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_41_io_pop_payload;
      7'b0101010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_42_io_pop_payload;
      7'b0101011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_43_io_pop_payload;
      7'b0101100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_44_io_pop_payload;
      7'b0101101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_45_io_pop_payload;
      7'b0101110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_46_io_pop_payload;
      7'b0101111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_47_io_pop_payload;
      7'b0110000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_48_io_pop_payload;
      7'b0110001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_49_io_pop_payload;
      7'b0110010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_50_io_pop_payload;
      7'b0110011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_51_io_pop_payload;
      7'b0110100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_52_io_pop_payload;
      7'b0110101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_53_io_pop_payload;
      7'b0110110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_54_io_pop_payload;
      7'b0110111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_55_io_pop_payload;
      7'b0111000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_56_io_pop_payload;
      7'b0111001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_57_io_pop_payload;
      7'b0111010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_58_io_pop_payload;
      7'b0111011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_59_io_pop_payload;
      7'b0111100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_60_io_pop_payload;
      7'b0111101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_61_io_pop_payload;
      7'b0111110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_62_io_pop_payload;
      7'b0111111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_63_io_pop_payload;
      7'b1000000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_64_io_pop_payload;
      7'b1000001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_65_io_pop_payload;
      7'b1000010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_66_io_pop_payload;
      7'b1000011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_67_io_pop_payload;
      7'b1000100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_68_io_pop_payload;
      7'b1000101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_69_io_pop_payload;
      7'b1000110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_70_io_pop_payload;
      7'b1000111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_71_io_pop_payload;
      7'b1001000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_72_io_pop_payload;
      7'b1001001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_73_io_pop_payload;
      7'b1001010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_74_io_pop_payload;
      7'b1001011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_75_io_pop_payload;
      7'b1001100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_76_io_pop_payload;
      7'b1001101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_77_io_pop_payload;
      7'b1001110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_78_io_pop_payload;
      7'b1001111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_79_io_pop_payload;
      7'b1010000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_80_io_pop_payload;
      7'b1010001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_81_io_pop_payload;
      7'b1010010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_82_io_pop_payload;
      7'b1010011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_83_io_pop_payload;
      7'b1010100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_84_io_pop_payload;
      7'b1010101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_85_io_pop_payload;
      7'b1010110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_86_io_pop_payload;
      7'b1010111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_87_io_pop_payload;
      7'b1011000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_88_io_pop_payload;
      7'b1011001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_89_io_pop_payload;
      7'b1011010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_90_io_pop_payload;
      7'b1011011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_91_io_pop_payload;
      7'b1011100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_92_io_pop_payload;
      7'b1011101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_93_io_pop_payload;
      7'b1011110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_94_io_pop_payload;
      7'b1011111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_95_io_pop_payload;
      7'b1100000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_96_io_pop_payload;
      7'b1100001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_97_io_pop_payload;
      7'b1100010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_98_io_pop_payload;
      7'b1100011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_99_io_pop_payload;
      7'b1100100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_100_io_pop_payload;
      7'b1100101 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_101_io_pop_payload;
      7'b1100110 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_102_io_pop_payload;
      7'b1100111 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_103_io_pop_payload;
      7'b1101000 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_104_io_pop_payload;
      7'b1101001 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_105_io_pop_payload;
      7'b1101010 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_106_io_pop_payload;
      7'b1101011 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_107_io_pop_payload;
      7'b1101100 : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_108_io_pop_payload;
      default : _zz_outputStreamArrayData_7_payload_2 = fifoGroup_109_io_pop_payload;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l240_7_1)
      7'b0000000 : _zz_when_ArraySlice_l240_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l240_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l240_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l240_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l240_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l240_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l240_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l240_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l240_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l240_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l240_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l240_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l240_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l240_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l240_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l240_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l240_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l240_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l240_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l240_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l240_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l240_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l240_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l240_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l240_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l240_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l240_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l240_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l240_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l240_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l240_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l240_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l240_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l240_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l240_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l240_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l240_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l240_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l240_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l240_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l240_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l240_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l240_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l240_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l240_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l240_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l240_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l240_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l240_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l240_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l240_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l240_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l240_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l240_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l240_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l240_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l240_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l240_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l240_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l240_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l240_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l240_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l240_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l240_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l240_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l240_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l240_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l240_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l240_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l240_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l240_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l240_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l240_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l240_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l240_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l240_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l240_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l240_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l240_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l240_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l240_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l240_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l240_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l240_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l240_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l240_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l240_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l240_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l240_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l240_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l240_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l240_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l240_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l240_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l240_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l240_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l240_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l240_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l240_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l240_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l240_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l240_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l240_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l240_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l240_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l240_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l240_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l240_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l240_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l240_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l249_7_1)
      7'b0000000 : _zz_when_ArraySlice_l249_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l249_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l249_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l249_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l249_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l249_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l249_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l249_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l249_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l249_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l249_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l249_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l249_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l249_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l249_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l249_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l249_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l249_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l249_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l249_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l249_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l249_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l249_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l249_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l249_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l249_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l249_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l249_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l249_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l249_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l249_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l249_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l249_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l249_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l249_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l249_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l249_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l249_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l249_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l249_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l249_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l249_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l249_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l249_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l249_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l249_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l249_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l249_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l249_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l249_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l249_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l249_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l249_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l249_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l249_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l249_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l249_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l249_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l249_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l249_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l249_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l249_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l249_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l249_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l249_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l249_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l249_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l249_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l249_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l249_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l249_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l249_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l249_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l249_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l249_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l249_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l249_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l249_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l249_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l249_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l249_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l249_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l249_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l249_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l249_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l249_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l249_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l249_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l249_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l249_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l249_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l249_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l249_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l249_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l249_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l249_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l249_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l249_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l249_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l249_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l249_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l249_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l249_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l249_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l249_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l249_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l249_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l249_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l249_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l249_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  always @(*) begin
    case(_zz_when_ArraySlice_l274_7_1)
      7'b0000000 : _zz_when_ArraySlice_l274_7 = fifoGroup_0_io_occupancy;
      7'b0000001 : _zz_when_ArraySlice_l274_7 = fifoGroup_1_io_occupancy;
      7'b0000010 : _zz_when_ArraySlice_l274_7 = fifoGroup_2_io_occupancy;
      7'b0000011 : _zz_when_ArraySlice_l274_7 = fifoGroup_3_io_occupancy;
      7'b0000100 : _zz_when_ArraySlice_l274_7 = fifoGroup_4_io_occupancy;
      7'b0000101 : _zz_when_ArraySlice_l274_7 = fifoGroup_5_io_occupancy;
      7'b0000110 : _zz_when_ArraySlice_l274_7 = fifoGroup_6_io_occupancy;
      7'b0000111 : _zz_when_ArraySlice_l274_7 = fifoGroup_7_io_occupancy;
      7'b0001000 : _zz_when_ArraySlice_l274_7 = fifoGroup_8_io_occupancy;
      7'b0001001 : _zz_when_ArraySlice_l274_7 = fifoGroup_9_io_occupancy;
      7'b0001010 : _zz_when_ArraySlice_l274_7 = fifoGroup_10_io_occupancy;
      7'b0001011 : _zz_when_ArraySlice_l274_7 = fifoGroup_11_io_occupancy;
      7'b0001100 : _zz_when_ArraySlice_l274_7 = fifoGroup_12_io_occupancy;
      7'b0001101 : _zz_when_ArraySlice_l274_7 = fifoGroup_13_io_occupancy;
      7'b0001110 : _zz_when_ArraySlice_l274_7 = fifoGroup_14_io_occupancy;
      7'b0001111 : _zz_when_ArraySlice_l274_7 = fifoGroup_15_io_occupancy;
      7'b0010000 : _zz_when_ArraySlice_l274_7 = fifoGroup_16_io_occupancy;
      7'b0010001 : _zz_when_ArraySlice_l274_7 = fifoGroup_17_io_occupancy;
      7'b0010010 : _zz_when_ArraySlice_l274_7 = fifoGroup_18_io_occupancy;
      7'b0010011 : _zz_when_ArraySlice_l274_7 = fifoGroup_19_io_occupancy;
      7'b0010100 : _zz_when_ArraySlice_l274_7 = fifoGroup_20_io_occupancy;
      7'b0010101 : _zz_when_ArraySlice_l274_7 = fifoGroup_21_io_occupancy;
      7'b0010110 : _zz_when_ArraySlice_l274_7 = fifoGroup_22_io_occupancy;
      7'b0010111 : _zz_when_ArraySlice_l274_7 = fifoGroup_23_io_occupancy;
      7'b0011000 : _zz_when_ArraySlice_l274_7 = fifoGroup_24_io_occupancy;
      7'b0011001 : _zz_when_ArraySlice_l274_7 = fifoGroup_25_io_occupancy;
      7'b0011010 : _zz_when_ArraySlice_l274_7 = fifoGroup_26_io_occupancy;
      7'b0011011 : _zz_when_ArraySlice_l274_7 = fifoGroup_27_io_occupancy;
      7'b0011100 : _zz_when_ArraySlice_l274_7 = fifoGroup_28_io_occupancy;
      7'b0011101 : _zz_when_ArraySlice_l274_7 = fifoGroup_29_io_occupancy;
      7'b0011110 : _zz_when_ArraySlice_l274_7 = fifoGroup_30_io_occupancy;
      7'b0011111 : _zz_when_ArraySlice_l274_7 = fifoGroup_31_io_occupancy;
      7'b0100000 : _zz_when_ArraySlice_l274_7 = fifoGroup_32_io_occupancy;
      7'b0100001 : _zz_when_ArraySlice_l274_7 = fifoGroup_33_io_occupancy;
      7'b0100010 : _zz_when_ArraySlice_l274_7 = fifoGroup_34_io_occupancy;
      7'b0100011 : _zz_when_ArraySlice_l274_7 = fifoGroup_35_io_occupancy;
      7'b0100100 : _zz_when_ArraySlice_l274_7 = fifoGroup_36_io_occupancy;
      7'b0100101 : _zz_when_ArraySlice_l274_7 = fifoGroup_37_io_occupancy;
      7'b0100110 : _zz_when_ArraySlice_l274_7 = fifoGroup_38_io_occupancy;
      7'b0100111 : _zz_when_ArraySlice_l274_7 = fifoGroup_39_io_occupancy;
      7'b0101000 : _zz_when_ArraySlice_l274_7 = fifoGroup_40_io_occupancy;
      7'b0101001 : _zz_when_ArraySlice_l274_7 = fifoGroup_41_io_occupancy;
      7'b0101010 : _zz_when_ArraySlice_l274_7 = fifoGroup_42_io_occupancy;
      7'b0101011 : _zz_when_ArraySlice_l274_7 = fifoGroup_43_io_occupancy;
      7'b0101100 : _zz_when_ArraySlice_l274_7 = fifoGroup_44_io_occupancy;
      7'b0101101 : _zz_when_ArraySlice_l274_7 = fifoGroup_45_io_occupancy;
      7'b0101110 : _zz_when_ArraySlice_l274_7 = fifoGroup_46_io_occupancy;
      7'b0101111 : _zz_when_ArraySlice_l274_7 = fifoGroup_47_io_occupancy;
      7'b0110000 : _zz_when_ArraySlice_l274_7 = fifoGroup_48_io_occupancy;
      7'b0110001 : _zz_when_ArraySlice_l274_7 = fifoGroup_49_io_occupancy;
      7'b0110010 : _zz_when_ArraySlice_l274_7 = fifoGroup_50_io_occupancy;
      7'b0110011 : _zz_when_ArraySlice_l274_7 = fifoGroup_51_io_occupancy;
      7'b0110100 : _zz_when_ArraySlice_l274_7 = fifoGroup_52_io_occupancy;
      7'b0110101 : _zz_when_ArraySlice_l274_7 = fifoGroup_53_io_occupancy;
      7'b0110110 : _zz_when_ArraySlice_l274_7 = fifoGroup_54_io_occupancy;
      7'b0110111 : _zz_when_ArraySlice_l274_7 = fifoGroup_55_io_occupancy;
      7'b0111000 : _zz_when_ArraySlice_l274_7 = fifoGroup_56_io_occupancy;
      7'b0111001 : _zz_when_ArraySlice_l274_7 = fifoGroup_57_io_occupancy;
      7'b0111010 : _zz_when_ArraySlice_l274_7 = fifoGroup_58_io_occupancy;
      7'b0111011 : _zz_when_ArraySlice_l274_7 = fifoGroup_59_io_occupancy;
      7'b0111100 : _zz_when_ArraySlice_l274_7 = fifoGroup_60_io_occupancy;
      7'b0111101 : _zz_when_ArraySlice_l274_7 = fifoGroup_61_io_occupancy;
      7'b0111110 : _zz_when_ArraySlice_l274_7 = fifoGroup_62_io_occupancy;
      7'b0111111 : _zz_when_ArraySlice_l274_7 = fifoGroup_63_io_occupancy;
      7'b1000000 : _zz_when_ArraySlice_l274_7 = fifoGroup_64_io_occupancy;
      7'b1000001 : _zz_when_ArraySlice_l274_7 = fifoGroup_65_io_occupancy;
      7'b1000010 : _zz_when_ArraySlice_l274_7 = fifoGroup_66_io_occupancy;
      7'b1000011 : _zz_when_ArraySlice_l274_7 = fifoGroup_67_io_occupancy;
      7'b1000100 : _zz_when_ArraySlice_l274_7 = fifoGroup_68_io_occupancy;
      7'b1000101 : _zz_when_ArraySlice_l274_7 = fifoGroup_69_io_occupancy;
      7'b1000110 : _zz_when_ArraySlice_l274_7 = fifoGroup_70_io_occupancy;
      7'b1000111 : _zz_when_ArraySlice_l274_7 = fifoGroup_71_io_occupancy;
      7'b1001000 : _zz_when_ArraySlice_l274_7 = fifoGroup_72_io_occupancy;
      7'b1001001 : _zz_when_ArraySlice_l274_7 = fifoGroup_73_io_occupancy;
      7'b1001010 : _zz_when_ArraySlice_l274_7 = fifoGroup_74_io_occupancy;
      7'b1001011 : _zz_when_ArraySlice_l274_7 = fifoGroup_75_io_occupancy;
      7'b1001100 : _zz_when_ArraySlice_l274_7 = fifoGroup_76_io_occupancy;
      7'b1001101 : _zz_when_ArraySlice_l274_7 = fifoGroup_77_io_occupancy;
      7'b1001110 : _zz_when_ArraySlice_l274_7 = fifoGroup_78_io_occupancy;
      7'b1001111 : _zz_when_ArraySlice_l274_7 = fifoGroup_79_io_occupancy;
      7'b1010000 : _zz_when_ArraySlice_l274_7 = fifoGroup_80_io_occupancy;
      7'b1010001 : _zz_when_ArraySlice_l274_7 = fifoGroup_81_io_occupancy;
      7'b1010010 : _zz_when_ArraySlice_l274_7 = fifoGroup_82_io_occupancy;
      7'b1010011 : _zz_when_ArraySlice_l274_7 = fifoGroup_83_io_occupancy;
      7'b1010100 : _zz_when_ArraySlice_l274_7 = fifoGroup_84_io_occupancy;
      7'b1010101 : _zz_when_ArraySlice_l274_7 = fifoGroup_85_io_occupancy;
      7'b1010110 : _zz_when_ArraySlice_l274_7 = fifoGroup_86_io_occupancy;
      7'b1010111 : _zz_when_ArraySlice_l274_7 = fifoGroup_87_io_occupancy;
      7'b1011000 : _zz_when_ArraySlice_l274_7 = fifoGroup_88_io_occupancy;
      7'b1011001 : _zz_when_ArraySlice_l274_7 = fifoGroup_89_io_occupancy;
      7'b1011010 : _zz_when_ArraySlice_l274_7 = fifoGroup_90_io_occupancy;
      7'b1011011 : _zz_when_ArraySlice_l274_7 = fifoGroup_91_io_occupancy;
      7'b1011100 : _zz_when_ArraySlice_l274_7 = fifoGroup_92_io_occupancy;
      7'b1011101 : _zz_when_ArraySlice_l274_7 = fifoGroup_93_io_occupancy;
      7'b1011110 : _zz_when_ArraySlice_l274_7 = fifoGroup_94_io_occupancy;
      7'b1011111 : _zz_when_ArraySlice_l274_7 = fifoGroup_95_io_occupancy;
      7'b1100000 : _zz_when_ArraySlice_l274_7 = fifoGroup_96_io_occupancy;
      7'b1100001 : _zz_when_ArraySlice_l274_7 = fifoGroup_97_io_occupancy;
      7'b1100010 : _zz_when_ArraySlice_l274_7 = fifoGroup_98_io_occupancy;
      7'b1100011 : _zz_when_ArraySlice_l274_7 = fifoGroup_99_io_occupancy;
      7'b1100100 : _zz_when_ArraySlice_l274_7 = fifoGroup_100_io_occupancy;
      7'b1100101 : _zz_when_ArraySlice_l274_7 = fifoGroup_101_io_occupancy;
      7'b1100110 : _zz_when_ArraySlice_l274_7 = fifoGroup_102_io_occupancy;
      7'b1100111 : _zz_when_ArraySlice_l274_7 = fifoGroup_103_io_occupancy;
      7'b1101000 : _zz_when_ArraySlice_l274_7 = fifoGroup_104_io_occupancy;
      7'b1101001 : _zz_when_ArraySlice_l274_7 = fifoGroup_105_io_occupancy;
      7'b1101010 : _zz_when_ArraySlice_l274_7 = fifoGroup_106_io_occupancy;
      7'b1101011 : _zz_when_ArraySlice_l274_7 = fifoGroup_107_io_occupancy;
      7'b1101100 : _zz_when_ArraySlice_l274_7 = fifoGroup_108_io_occupancy;
      default : _zz_when_ArraySlice_l274_7 = fifoGroup_109_io_occupancy;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_BOOT : arraySliceStateMachine_stateReg_string = "BOOT         ";
      arraySliceStateMachine_enumDef_writeDataOnly : arraySliceStateMachine_stateReg_string = "writeDataOnly";
      arraySliceStateMachine_enumDef_readDataOnly : arraySliceStateMachine_stateReg_string = "readDataOnly ";
      arraySliceStateMachine_enumDef_readWriteData : arraySliceStateMachine_stateReg_string = "readWriteData";
      default : arraySliceStateMachine_stateReg_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(arraySliceStateMachine_stateNext)
      arraySliceStateMachine_enumDef_BOOT : arraySliceStateMachine_stateNext_string = "BOOT         ";
      arraySliceStateMachine_enumDef_writeDataOnly : arraySliceStateMachine_stateNext_string = "writeDataOnly";
      arraySliceStateMachine_enumDef_readDataOnly : arraySliceStateMachine_stateNext_string = "readDataOnly ";
      arraySliceStateMachine_enumDef_readWriteData : arraySliceStateMachine_stateNext_string = "readWriteData";
      default : arraySliceStateMachine_stateNext_string = "?????????????";
    endcase
  end
  `endif

  always @(*) begin
    handshakeTimes_0_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_0_fire_6) begin
          if(!when_ArraySlice_l468) begin
            handshakeTimes_0_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_0_fire_13) begin
          if(!when_ArraySlice_l325) begin
            handshakeTimes_0_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_0_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_0_fire_6) begin
          if(when_ArraySlice_l468) begin
            handshakeTimes_0_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_0_fire_13) begin
          if(when_ArraySlice_l325) begin
            handshakeTimes_0_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_0_willOverflowIfInc = (handshakeTimes_0_value == 13'h1bee);
  assign handshakeTimes_0_willOverflow = (handshakeTimes_0_willOverflowIfInc && handshakeTimes_0_willIncrement);
  always @(*) begin
    if(handshakeTimes_0_willOverflow) begin
      handshakeTimes_0_valueNext = 13'h0;
    end else begin
      handshakeTimes_0_valueNext = (handshakeTimes_0_value + _zz_handshakeTimes_0_valueNext);
    end
    if(handshakeTimes_0_willClear) begin
      handshakeTimes_0_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_1_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_1_fire_6) begin
          if(!when_ArraySlice_l468_1) begin
            handshakeTimes_1_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_1_fire_13) begin
          if(!when_ArraySlice_l325_1) begin
            handshakeTimes_1_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_1_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_1_fire_6) begin
          if(when_ArraySlice_l468_1) begin
            handshakeTimes_1_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_1_fire_13) begin
          if(when_ArraySlice_l325_1) begin
            handshakeTimes_1_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_1_willOverflowIfInc = (handshakeTimes_1_value == 13'h1bee);
  assign handshakeTimes_1_willOverflow = (handshakeTimes_1_willOverflowIfInc && handshakeTimes_1_willIncrement);
  always @(*) begin
    if(handshakeTimes_1_willOverflow) begin
      handshakeTimes_1_valueNext = 13'h0;
    end else begin
      handshakeTimes_1_valueNext = (handshakeTimes_1_value + _zz_handshakeTimes_1_valueNext);
    end
    if(handshakeTimes_1_willClear) begin
      handshakeTimes_1_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_2_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_2_fire_6) begin
          if(!when_ArraySlice_l468_2) begin
            handshakeTimes_2_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_2_fire_13) begin
          if(!when_ArraySlice_l325_2) begin
            handshakeTimes_2_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_2_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_2_fire_6) begin
          if(when_ArraySlice_l468_2) begin
            handshakeTimes_2_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_2_fire_13) begin
          if(when_ArraySlice_l325_2) begin
            handshakeTimes_2_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_2_willOverflowIfInc = (handshakeTimes_2_value == 13'h1bee);
  assign handshakeTimes_2_willOverflow = (handshakeTimes_2_willOverflowIfInc && handshakeTimes_2_willIncrement);
  always @(*) begin
    if(handshakeTimes_2_willOverflow) begin
      handshakeTimes_2_valueNext = 13'h0;
    end else begin
      handshakeTimes_2_valueNext = (handshakeTimes_2_value + _zz_handshakeTimes_2_valueNext);
    end
    if(handshakeTimes_2_willClear) begin
      handshakeTimes_2_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_3_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_3_fire_6) begin
          if(!when_ArraySlice_l468_3) begin
            handshakeTimes_3_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_3_fire_13) begin
          if(!when_ArraySlice_l325_3) begin
            handshakeTimes_3_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_3_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_3_fire_6) begin
          if(when_ArraySlice_l468_3) begin
            handshakeTimes_3_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_3_fire_13) begin
          if(when_ArraySlice_l325_3) begin
            handshakeTimes_3_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_3_willOverflowIfInc = (handshakeTimes_3_value == 13'h1bee);
  assign handshakeTimes_3_willOverflow = (handshakeTimes_3_willOverflowIfInc && handshakeTimes_3_willIncrement);
  always @(*) begin
    if(handshakeTimes_3_willOverflow) begin
      handshakeTimes_3_valueNext = 13'h0;
    end else begin
      handshakeTimes_3_valueNext = (handshakeTimes_3_value + _zz_handshakeTimes_3_valueNext);
    end
    if(handshakeTimes_3_willClear) begin
      handshakeTimes_3_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_4_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_4_fire_6) begin
          if(!when_ArraySlice_l468_4) begin
            handshakeTimes_4_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_4_fire_13) begin
          if(!when_ArraySlice_l325_4) begin
            handshakeTimes_4_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_4_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_4_fire_6) begin
          if(when_ArraySlice_l468_4) begin
            handshakeTimes_4_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_4_fire_13) begin
          if(when_ArraySlice_l325_4) begin
            handshakeTimes_4_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_4_willOverflowIfInc = (handshakeTimes_4_value == 13'h1bee);
  assign handshakeTimes_4_willOverflow = (handshakeTimes_4_willOverflowIfInc && handshakeTimes_4_willIncrement);
  always @(*) begin
    if(handshakeTimes_4_willOverflow) begin
      handshakeTimes_4_valueNext = 13'h0;
    end else begin
      handshakeTimes_4_valueNext = (handshakeTimes_4_value + _zz_handshakeTimes_4_valueNext);
    end
    if(handshakeTimes_4_willClear) begin
      handshakeTimes_4_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_5_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_5_fire_6) begin
          if(!when_ArraySlice_l468_5) begin
            handshakeTimes_5_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_5_fire_13) begin
          if(!when_ArraySlice_l325_5) begin
            handshakeTimes_5_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_5_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_5_fire_6) begin
          if(when_ArraySlice_l468_5) begin
            handshakeTimes_5_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_5_fire_13) begin
          if(when_ArraySlice_l325_5) begin
            handshakeTimes_5_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_5_willOverflowIfInc = (handshakeTimes_5_value == 13'h1bee);
  assign handshakeTimes_5_willOverflow = (handshakeTimes_5_willOverflowIfInc && handshakeTimes_5_willIncrement);
  always @(*) begin
    if(handshakeTimes_5_willOverflow) begin
      handshakeTimes_5_valueNext = 13'h0;
    end else begin
      handshakeTimes_5_valueNext = (handshakeTimes_5_value + _zz_handshakeTimes_5_valueNext);
    end
    if(handshakeTimes_5_willClear) begin
      handshakeTimes_5_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_6_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_6_fire_6) begin
          if(!when_ArraySlice_l468_6) begin
            handshakeTimes_6_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_6_fire_13) begin
          if(!when_ArraySlice_l325_6) begin
            handshakeTimes_6_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_6_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_6_fire_6) begin
          if(when_ArraySlice_l468_6) begin
            handshakeTimes_6_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_6_fire_13) begin
          if(when_ArraySlice_l325_6) begin
            handshakeTimes_6_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_6_willOverflowIfInc = (handshakeTimes_6_value == 13'h1bee);
  assign handshakeTimes_6_willOverflow = (handshakeTimes_6_willOverflowIfInc && handshakeTimes_6_willIncrement);
  always @(*) begin
    if(handshakeTimes_6_willOverflow) begin
      handshakeTimes_6_valueNext = 13'h0;
    end else begin
      handshakeTimes_6_valueNext = (handshakeTimes_6_value + _zz_handshakeTimes_6_valueNext);
    end
    if(handshakeTimes_6_willClear) begin
      handshakeTimes_6_valueNext = 13'h0;
    end
  end

  always @(*) begin
    handshakeTimes_7_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_7_fire_6) begin
          if(!when_ArraySlice_l468_7) begin
            handshakeTimes_7_willIncrement = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_7_fire_13) begin
          if(!when_ArraySlice_l325_7) begin
            handshakeTimes_7_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    handshakeTimes_7_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(outputStreamArrayData_7_fire_6) begin
          if(when_ArraySlice_l468_7) begin
            handshakeTimes_7_willClear = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(outputStreamArrayData_7_fire_13) begin
          if(when_ArraySlice_l325_7) begin
            handshakeTimes_7_willClear = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign handshakeTimes_7_willOverflowIfInc = (handshakeTimes_7_value == 13'h1bee);
  assign handshakeTimes_7_willOverflow = (handshakeTimes_7_willOverflowIfInc && handshakeTimes_7_willIncrement);
  always @(*) begin
    if(handshakeTimes_7_willOverflow) begin
      handshakeTimes_7_valueNext = 13'h0;
    end else begin
      handshakeTimes_7_valueNext = (handshakeTimes_7_value + _zz_handshakeTimes_7_valueNext);
    end
    if(handshakeTimes_7_willClear) begin
      handshakeTimes_7_valueNext = 13'h0;
    end
  end

  always @(*) begin
    outSliceNumb_0_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l382) begin
            if(when_ArraySlice_l383) begin
              if(when_ArraySlice_l384) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392) begin
              if(when_ArraySlice_l393) begin
                if(when_ArraySlice_l395) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417) begin
              if(when_ArraySlice_l418) begin
                if(when_ArraySlice_l420) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447) begin
            if(when_ArraySlice_l449) begin
              if(when_ArraySlice_l450) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l239) begin
            if(when_ArraySlice_l240) begin
              if(when_ArraySlice_l241) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249) begin
              if(when_ArraySlice_l250) begin
                if(when_ArraySlice_l252) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274) begin
              if(when_ArraySlice_l275) begin
                if(when_ArraySlice_l277) begin
                  outSliceNumb_0_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304) begin
            if(when_ArraySlice_l306) begin
              if(when_ArraySlice_l307) begin
                outSliceNumb_0_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_0_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l382) begin
            if(when_ArraySlice_l392) begin
              if(when_ArraySlice_l393) begin
                if(!when_ArraySlice_l395) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417) begin
              if(when_ArraySlice_l418) begin
                if(!when_ArraySlice_l420) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447) begin
            if(when_ArraySlice_l449) begin
              if(!when_ArraySlice_l450) begin
                outSliceNumb_0_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l239) begin
            if(when_ArraySlice_l249) begin
              if(when_ArraySlice_l250) begin
                if(!when_ArraySlice_l252) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274) begin
              if(when_ArraySlice_l275) begin
                if(!when_ArraySlice_l277) begin
                  outSliceNumb_0_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304) begin
            if(when_ArraySlice_l306) begin
              if(!when_ArraySlice_l307) begin
                outSliceNumb_0_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_0_willOverflowIfInc = (outSliceNumb_0_value == 7'h41);
  assign outSliceNumb_0_willOverflow = (outSliceNumb_0_willOverflowIfInc && outSliceNumb_0_willIncrement);
  always @(*) begin
    if(outSliceNumb_0_willOverflow) begin
      outSliceNumb_0_valueNext = 7'h0;
    end else begin
      outSliceNumb_0_valueNext = (outSliceNumb_0_value + _zz_outSliceNumb_0_valueNext);
    end
    if(outSliceNumb_0_willClear) begin
      outSliceNumb_0_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_1_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l382_1) begin
            if(when_ArraySlice_l383_1) begin
              if(when_ArraySlice_l384_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_1) begin
              if(when_ArraySlice_l393_1) begin
                if(when_ArraySlice_l395_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_1) begin
              if(when_ArraySlice_l418_1) begin
                if(when_ArraySlice_l420_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_1) begin
            if(when_ArraySlice_l449_1) begin
              if(when_ArraySlice_l450_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l239_1) begin
            if(when_ArraySlice_l240_1) begin
              if(when_ArraySlice_l241_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_1) begin
              if(when_ArraySlice_l250_1) begin
                if(when_ArraySlice_l252_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_1) begin
              if(when_ArraySlice_l275_1) begin
                if(when_ArraySlice_l277_1) begin
                  outSliceNumb_1_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_1) begin
            if(when_ArraySlice_l306_1) begin
              if(when_ArraySlice_l307_1) begin
                outSliceNumb_1_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_1_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l382_1) begin
            if(when_ArraySlice_l392_1) begin
              if(when_ArraySlice_l393_1) begin
                if(!when_ArraySlice_l395_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_1) begin
              if(when_ArraySlice_l418_1) begin
                if(!when_ArraySlice_l420_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_1) begin
            if(when_ArraySlice_l449_1) begin
              if(!when_ArraySlice_l450_1) begin
                outSliceNumb_1_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l239_1) begin
            if(when_ArraySlice_l249_1) begin
              if(when_ArraySlice_l250_1) begin
                if(!when_ArraySlice_l252_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_1) begin
              if(when_ArraySlice_l275_1) begin
                if(!when_ArraySlice_l277_1) begin
                  outSliceNumb_1_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_1) begin
            if(when_ArraySlice_l306_1) begin
              if(!when_ArraySlice_l307_1) begin
                outSliceNumb_1_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_1_willOverflowIfInc = (outSliceNumb_1_value == 7'h41);
  assign outSliceNumb_1_willOverflow = (outSliceNumb_1_willOverflowIfInc && outSliceNumb_1_willIncrement);
  always @(*) begin
    if(outSliceNumb_1_willOverflow) begin
      outSliceNumb_1_valueNext = 7'h0;
    end else begin
      outSliceNumb_1_valueNext = (outSliceNumb_1_value + _zz_outSliceNumb_1_valueNext);
    end
    if(outSliceNumb_1_willClear) begin
      outSliceNumb_1_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_2_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l382_2) begin
            if(when_ArraySlice_l383_2) begin
              if(when_ArraySlice_l384_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_2) begin
              if(when_ArraySlice_l393_2) begin
                if(when_ArraySlice_l395_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_2) begin
              if(when_ArraySlice_l418_2) begin
                if(when_ArraySlice_l420_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_2) begin
            if(when_ArraySlice_l449_2) begin
              if(when_ArraySlice_l450_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l239_2) begin
            if(when_ArraySlice_l240_2) begin
              if(when_ArraySlice_l241_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_2) begin
              if(when_ArraySlice_l250_2) begin
                if(when_ArraySlice_l252_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_2) begin
              if(when_ArraySlice_l275_2) begin
                if(when_ArraySlice_l277_2) begin
                  outSliceNumb_2_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_2) begin
            if(when_ArraySlice_l306_2) begin
              if(when_ArraySlice_l307_2) begin
                outSliceNumb_2_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_2_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l382_2) begin
            if(when_ArraySlice_l392_2) begin
              if(when_ArraySlice_l393_2) begin
                if(!when_ArraySlice_l395_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_2) begin
              if(when_ArraySlice_l418_2) begin
                if(!when_ArraySlice_l420_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_2) begin
            if(when_ArraySlice_l449_2) begin
              if(!when_ArraySlice_l450_2) begin
                outSliceNumb_2_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l239_2) begin
            if(when_ArraySlice_l249_2) begin
              if(when_ArraySlice_l250_2) begin
                if(!when_ArraySlice_l252_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_2) begin
              if(when_ArraySlice_l275_2) begin
                if(!when_ArraySlice_l277_2) begin
                  outSliceNumb_2_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_2) begin
            if(when_ArraySlice_l306_2) begin
              if(!when_ArraySlice_l307_2) begin
                outSliceNumb_2_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_2_willOverflowIfInc = (outSliceNumb_2_value == 7'h41);
  assign outSliceNumb_2_willOverflow = (outSliceNumb_2_willOverflowIfInc && outSliceNumb_2_willIncrement);
  always @(*) begin
    if(outSliceNumb_2_willOverflow) begin
      outSliceNumb_2_valueNext = 7'h0;
    end else begin
      outSliceNumb_2_valueNext = (outSliceNumb_2_value + _zz_outSliceNumb_2_valueNext);
    end
    if(outSliceNumb_2_willClear) begin
      outSliceNumb_2_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_3_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l382_3) begin
            if(when_ArraySlice_l383_3) begin
              if(when_ArraySlice_l384_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_3) begin
              if(when_ArraySlice_l393_3) begin
                if(when_ArraySlice_l395_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_3) begin
              if(when_ArraySlice_l418_3) begin
                if(when_ArraySlice_l420_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_3) begin
            if(when_ArraySlice_l449_3) begin
              if(when_ArraySlice_l450_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l239_3) begin
            if(when_ArraySlice_l240_3) begin
              if(when_ArraySlice_l241_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_3) begin
              if(when_ArraySlice_l250_3) begin
                if(when_ArraySlice_l252_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_3) begin
              if(when_ArraySlice_l275_3) begin
                if(when_ArraySlice_l277_3) begin
                  outSliceNumb_3_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_3) begin
            if(when_ArraySlice_l306_3) begin
              if(when_ArraySlice_l307_3) begin
                outSliceNumb_3_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_3_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l382_3) begin
            if(when_ArraySlice_l392_3) begin
              if(when_ArraySlice_l393_3) begin
                if(!when_ArraySlice_l395_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_3) begin
              if(when_ArraySlice_l418_3) begin
                if(!when_ArraySlice_l420_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_3) begin
            if(when_ArraySlice_l449_3) begin
              if(!when_ArraySlice_l450_3) begin
                outSliceNumb_3_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l239_3) begin
            if(when_ArraySlice_l249_3) begin
              if(when_ArraySlice_l250_3) begin
                if(!when_ArraySlice_l252_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_3) begin
              if(when_ArraySlice_l275_3) begin
                if(!when_ArraySlice_l277_3) begin
                  outSliceNumb_3_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_3) begin
            if(when_ArraySlice_l306_3) begin
              if(!when_ArraySlice_l307_3) begin
                outSliceNumb_3_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_3_willOverflowIfInc = (outSliceNumb_3_value == 7'h41);
  assign outSliceNumb_3_willOverflow = (outSliceNumb_3_willOverflowIfInc && outSliceNumb_3_willIncrement);
  always @(*) begin
    if(outSliceNumb_3_willOverflow) begin
      outSliceNumb_3_valueNext = 7'h0;
    end else begin
      outSliceNumb_3_valueNext = (outSliceNumb_3_value + _zz_outSliceNumb_3_valueNext);
    end
    if(outSliceNumb_3_willClear) begin
      outSliceNumb_3_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_4_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l382_4) begin
            if(when_ArraySlice_l383_4) begin
              if(when_ArraySlice_l384_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_4) begin
              if(when_ArraySlice_l393_4) begin
                if(when_ArraySlice_l395_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_4) begin
              if(when_ArraySlice_l418_4) begin
                if(when_ArraySlice_l420_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_4) begin
            if(when_ArraySlice_l449_4) begin
              if(when_ArraySlice_l450_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l239_4) begin
            if(when_ArraySlice_l240_4) begin
              if(when_ArraySlice_l241_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_4) begin
              if(when_ArraySlice_l250_4) begin
                if(when_ArraySlice_l252_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_4) begin
              if(when_ArraySlice_l275_4) begin
                if(when_ArraySlice_l277_4) begin
                  outSliceNumb_4_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_4) begin
            if(when_ArraySlice_l306_4) begin
              if(when_ArraySlice_l307_4) begin
                outSliceNumb_4_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_4_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l382_4) begin
            if(when_ArraySlice_l392_4) begin
              if(when_ArraySlice_l393_4) begin
                if(!when_ArraySlice_l395_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_4) begin
              if(when_ArraySlice_l418_4) begin
                if(!when_ArraySlice_l420_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_4) begin
            if(when_ArraySlice_l449_4) begin
              if(!when_ArraySlice_l450_4) begin
                outSliceNumb_4_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l239_4) begin
            if(when_ArraySlice_l249_4) begin
              if(when_ArraySlice_l250_4) begin
                if(!when_ArraySlice_l252_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_4) begin
              if(when_ArraySlice_l275_4) begin
                if(!when_ArraySlice_l277_4) begin
                  outSliceNumb_4_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_4) begin
            if(when_ArraySlice_l306_4) begin
              if(!when_ArraySlice_l307_4) begin
                outSliceNumb_4_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_4_willOverflowIfInc = (outSliceNumb_4_value == 7'h41);
  assign outSliceNumb_4_willOverflow = (outSliceNumb_4_willOverflowIfInc && outSliceNumb_4_willIncrement);
  always @(*) begin
    if(outSliceNumb_4_willOverflow) begin
      outSliceNumb_4_valueNext = 7'h0;
    end else begin
      outSliceNumb_4_valueNext = (outSliceNumb_4_value + _zz_outSliceNumb_4_valueNext);
    end
    if(outSliceNumb_4_willClear) begin
      outSliceNumb_4_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_5_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l382_5) begin
            if(when_ArraySlice_l383_5) begin
              if(when_ArraySlice_l384_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_5) begin
              if(when_ArraySlice_l393_5) begin
                if(when_ArraySlice_l395_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_5) begin
              if(when_ArraySlice_l418_5) begin
                if(when_ArraySlice_l420_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_5) begin
            if(when_ArraySlice_l449_5) begin
              if(when_ArraySlice_l450_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l239_5) begin
            if(when_ArraySlice_l240_5) begin
              if(when_ArraySlice_l241_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_5) begin
              if(when_ArraySlice_l250_5) begin
                if(when_ArraySlice_l252_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_5) begin
              if(when_ArraySlice_l275_5) begin
                if(when_ArraySlice_l277_5) begin
                  outSliceNumb_5_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_5) begin
            if(when_ArraySlice_l306_5) begin
              if(when_ArraySlice_l307_5) begin
                outSliceNumb_5_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_5_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l382_5) begin
            if(when_ArraySlice_l392_5) begin
              if(when_ArraySlice_l393_5) begin
                if(!when_ArraySlice_l395_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_5) begin
              if(when_ArraySlice_l418_5) begin
                if(!when_ArraySlice_l420_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_5) begin
            if(when_ArraySlice_l449_5) begin
              if(!when_ArraySlice_l450_5) begin
                outSliceNumb_5_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l239_5) begin
            if(when_ArraySlice_l249_5) begin
              if(when_ArraySlice_l250_5) begin
                if(!when_ArraySlice_l252_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_5) begin
              if(when_ArraySlice_l275_5) begin
                if(!when_ArraySlice_l277_5) begin
                  outSliceNumb_5_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_5) begin
            if(when_ArraySlice_l306_5) begin
              if(!when_ArraySlice_l307_5) begin
                outSliceNumb_5_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_5_willOverflowIfInc = (outSliceNumb_5_value == 7'h41);
  assign outSliceNumb_5_willOverflow = (outSliceNumb_5_willOverflowIfInc && outSliceNumb_5_willIncrement);
  always @(*) begin
    if(outSliceNumb_5_willOverflow) begin
      outSliceNumb_5_valueNext = 7'h0;
    end else begin
      outSliceNumb_5_valueNext = (outSliceNumb_5_value + _zz_outSliceNumb_5_valueNext);
    end
    if(outSliceNumb_5_willClear) begin
      outSliceNumb_5_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_6_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l382_6) begin
            if(when_ArraySlice_l383_6) begin
              if(when_ArraySlice_l384_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_6) begin
              if(when_ArraySlice_l393_6) begin
                if(when_ArraySlice_l395_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_6) begin
              if(when_ArraySlice_l418_6) begin
                if(when_ArraySlice_l420_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_6) begin
            if(when_ArraySlice_l449_6) begin
              if(when_ArraySlice_l450_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l239_6) begin
            if(when_ArraySlice_l240_6) begin
              if(when_ArraySlice_l241_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_6) begin
              if(when_ArraySlice_l250_6) begin
                if(when_ArraySlice_l252_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_6) begin
              if(when_ArraySlice_l275_6) begin
                if(when_ArraySlice_l277_6) begin
                  outSliceNumb_6_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_6) begin
            if(when_ArraySlice_l306_6) begin
              if(when_ArraySlice_l307_6) begin
                outSliceNumb_6_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_6_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l382_6) begin
            if(when_ArraySlice_l392_6) begin
              if(when_ArraySlice_l393_6) begin
                if(!when_ArraySlice_l395_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_6) begin
              if(when_ArraySlice_l418_6) begin
                if(!when_ArraySlice_l420_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_6) begin
            if(when_ArraySlice_l449_6) begin
              if(!when_ArraySlice_l450_6) begin
                outSliceNumb_6_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l239_6) begin
            if(when_ArraySlice_l249_6) begin
              if(when_ArraySlice_l250_6) begin
                if(!when_ArraySlice_l252_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_6) begin
              if(when_ArraySlice_l275_6) begin
                if(!when_ArraySlice_l277_6) begin
                  outSliceNumb_6_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_6) begin
            if(when_ArraySlice_l306_6) begin
              if(!when_ArraySlice_l307_6) begin
                outSliceNumb_6_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_6_willOverflowIfInc = (outSliceNumb_6_value == 7'h41);
  assign outSliceNumb_6_willOverflow = (outSliceNumb_6_willOverflowIfInc && outSliceNumb_6_willIncrement);
  always @(*) begin
    if(outSliceNumb_6_willOverflow) begin
      outSliceNumb_6_valueNext = 7'h0;
    end else begin
      outSliceNumb_6_valueNext = (outSliceNumb_6_value + _zz_outSliceNumb_6_valueNext);
    end
    if(outSliceNumb_6_willClear) begin
      outSliceNumb_6_valueNext = 7'h0;
    end
  end

  always @(*) begin
    outSliceNumb_7_willIncrement = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l382_7) begin
            if(when_ArraySlice_l383_7) begin
              if(when_ArraySlice_l384_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l392_7) begin
              if(when_ArraySlice_l393_7) begin
                if(when_ArraySlice_l395_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_7) begin
              if(when_ArraySlice_l418_7) begin
                if(when_ArraySlice_l420_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_7) begin
            if(when_ArraySlice_l449_7) begin
              if(when_ArraySlice_l450_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l239_7) begin
            if(when_ArraySlice_l240_7) begin
              if(when_ArraySlice_l241_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
            if(when_ArraySlice_l249_7) begin
              if(when_ArraySlice_l250_7) begin
                if(when_ArraySlice_l252_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_7) begin
              if(when_ArraySlice_l275_7) begin
                if(when_ArraySlice_l277_7) begin
                  outSliceNumb_7_willIncrement = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_7) begin
            if(when_ArraySlice_l306_7) begin
              if(when_ArraySlice_l307_7) begin
                outSliceNumb_7_willIncrement = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outSliceNumb_7_willClear = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l382_7) begin
            if(when_ArraySlice_l392_7) begin
              if(when_ArraySlice_l393_7) begin
                if(!when_ArraySlice_l395_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l417_7) begin
              if(when_ArraySlice_l418_7) begin
                if(!when_ArraySlice_l420_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l447_7) begin
            if(when_ArraySlice_l449_7) begin
              if(!when_ArraySlice_l450_7) begin
                outSliceNumb_7_willClear = 1'b1;
              end
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l239_7) begin
            if(when_ArraySlice_l249_7) begin
              if(when_ArraySlice_l250_7) begin
                if(!when_ArraySlice_l252_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
            if(when_ArraySlice_l274_7) begin
              if(when_ArraySlice_l275_7) begin
                if(!when_ArraySlice_l277_7) begin
                  outSliceNumb_7_willClear = 1'b1;
                end
              end
            end
          end
        end else begin
          if(when_ArraySlice_l304_7) begin
            if(when_ArraySlice_l306_7) begin
              if(!when_ArraySlice_l307_7) begin
                outSliceNumb_7_willClear = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign outSliceNumb_7_willOverflowIfInc = (outSliceNumb_7_value == 7'h41);
  assign outSliceNumb_7_willOverflow = (outSliceNumb_7_willOverflowIfInc && outSliceNumb_7_willIncrement);
  always @(*) begin
    if(outSliceNumb_7_willOverflow) begin
      outSliceNumb_7_valueNext = 7'h0;
    end else begin
      outSliceNumb_7_valueNext = (outSliceNumb_7_value + _zz_outSliceNumb_7_valueNext);
    end
    if(outSliceNumb_7_willClear) begin
      outSliceNumb_7_valueNext = 7'h0;
    end
  end

  always @(*) begin
    inputStreamArrayData_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          inputStreamArrayData_ready = _zz_inputStreamArrayData_ready;
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            inputStreamArrayData_ready = _zz_inputStreamArrayData_ready_1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_0_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            outputStreamArrayData_0_valid = _zz_outputStreamArrayData_0_valid_2;
          end
          if(when_ArraySlice_l382) begin
            if(when_ArraySlice_l417) begin
              outputStreamArrayData_0_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447) begin
            outputStreamArrayData_0_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            outputStreamArrayData_0_valid = _zz_outputStreamArrayData_0_valid_4;
          end
          if(when_ArraySlice_l239) begin
            if(when_ArraySlice_l274) begin
              outputStreamArrayData_0_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304) begin
            outputStreamArrayData_0_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_0_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            outputStreamArrayData_0_payload = _zz_outputStreamArrayData_0_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            outputStreamArrayData_0_payload = _zz_outputStreamArrayData_0_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_1_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            outputStreamArrayData_1_valid = _zz_outputStreamArrayData_1_valid_2;
          end
          if(when_ArraySlice_l382_1) begin
            if(when_ArraySlice_l417_1) begin
              outputStreamArrayData_1_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_1) begin
            outputStreamArrayData_1_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            outputStreamArrayData_1_valid = _zz_outputStreamArrayData_1_valid_4;
          end
          if(when_ArraySlice_l239_1) begin
            if(when_ArraySlice_l274_1) begin
              outputStreamArrayData_1_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_1) begin
            outputStreamArrayData_1_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_1_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            outputStreamArrayData_1_payload = _zz_outputStreamArrayData_1_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            outputStreamArrayData_1_payload = _zz_outputStreamArrayData_1_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_2_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            outputStreamArrayData_2_valid = _zz_outputStreamArrayData_2_valid_2;
          end
          if(when_ArraySlice_l382_2) begin
            if(when_ArraySlice_l417_2) begin
              outputStreamArrayData_2_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_2) begin
            outputStreamArrayData_2_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            outputStreamArrayData_2_valid = _zz_outputStreamArrayData_2_valid_4;
          end
          if(when_ArraySlice_l239_2) begin
            if(when_ArraySlice_l274_2) begin
              outputStreamArrayData_2_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_2) begin
            outputStreamArrayData_2_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_2_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            outputStreamArrayData_2_payload = _zz_outputStreamArrayData_2_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            outputStreamArrayData_2_payload = _zz_outputStreamArrayData_2_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_3_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            outputStreamArrayData_3_valid = _zz_outputStreamArrayData_3_valid_2;
          end
          if(when_ArraySlice_l382_3) begin
            if(when_ArraySlice_l417_3) begin
              outputStreamArrayData_3_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_3) begin
            outputStreamArrayData_3_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            outputStreamArrayData_3_valid = _zz_outputStreamArrayData_3_valid_4;
          end
          if(when_ArraySlice_l239_3) begin
            if(when_ArraySlice_l274_3) begin
              outputStreamArrayData_3_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_3) begin
            outputStreamArrayData_3_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_3_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            outputStreamArrayData_3_payload = _zz_outputStreamArrayData_3_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            outputStreamArrayData_3_payload = _zz_outputStreamArrayData_3_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_4_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            outputStreamArrayData_4_valid = _zz_outputStreamArrayData_4_valid_2;
          end
          if(when_ArraySlice_l382_4) begin
            if(when_ArraySlice_l417_4) begin
              outputStreamArrayData_4_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_4) begin
            outputStreamArrayData_4_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            outputStreamArrayData_4_valid = _zz_outputStreamArrayData_4_valid_4;
          end
          if(when_ArraySlice_l239_4) begin
            if(when_ArraySlice_l274_4) begin
              outputStreamArrayData_4_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_4) begin
            outputStreamArrayData_4_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_4_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            outputStreamArrayData_4_payload = _zz_outputStreamArrayData_4_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            outputStreamArrayData_4_payload = _zz_outputStreamArrayData_4_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_5_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            outputStreamArrayData_5_valid = _zz_outputStreamArrayData_5_valid_2;
          end
          if(when_ArraySlice_l382_5) begin
            if(when_ArraySlice_l417_5) begin
              outputStreamArrayData_5_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_5) begin
            outputStreamArrayData_5_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            outputStreamArrayData_5_valid = _zz_outputStreamArrayData_5_valid_4;
          end
          if(when_ArraySlice_l239_5) begin
            if(when_ArraySlice_l274_5) begin
              outputStreamArrayData_5_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_5) begin
            outputStreamArrayData_5_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_5_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            outputStreamArrayData_5_payload = _zz_outputStreamArrayData_5_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            outputStreamArrayData_5_payload = _zz_outputStreamArrayData_5_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_6_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            outputStreamArrayData_6_valid = _zz_outputStreamArrayData_6_valid_2;
          end
          if(when_ArraySlice_l382_6) begin
            if(when_ArraySlice_l417_6) begin
              outputStreamArrayData_6_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_6) begin
            outputStreamArrayData_6_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            outputStreamArrayData_6_valid = _zz_outputStreamArrayData_6_valid_4;
          end
          if(when_ArraySlice_l239_6) begin
            if(when_ArraySlice_l274_6) begin
              outputStreamArrayData_6_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_6) begin
            outputStreamArrayData_6_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_6_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            outputStreamArrayData_6_payload = _zz_outputStreamArrayData_6_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            outputStreamArrayData_6_payload = _zz_outputStreamArrayData_6_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_7_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            outputStreamArrayData_7_valid = _zz_outputStreamArrayData_7_valid_2;
          end
          if(when_ArraySlice_l382_7) begin
            if(when_ArraySlice_l417_7) begin
              outputStreamArrayData_7_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l447_7) begin
            outputStreamArrayData_7_valid = 1'b1;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            outputStreamArrayData_7_valid = _zz_outputStreamArrayData_7_valid_4;
          end
          if(when_ArraySlice_l239_7) begin
            if(when_ArraySlice_l274_7) begin
              outputStreamArrayData_7_valid = 1'b1;
            end
          end
        end else begin
          if(when_ArraySlice_l304_7) begin
            outputStreamArrayData_7_valid = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputStreamArrayData_7_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            outputStreamArrayData_7_payload = _zz_outputStreamArrayData_7_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            outputStreamArrayData_7_payload = _zz_outputStreamArrayData_7_payload_2;
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[0]) begin
            fifoGroup_0_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[0]) begin
              fifoGroup_0_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[0]) begin
            fifoGroup_0_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[0]) begin
              fifoGroup_0_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_0_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[0]) begin
              fifoGroup_0_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[1]) begin
            fifoGroup_1_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[1]) begin
              fifoGroup_1_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[1]) begin
            fifoGroup_1_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[1]) begin
              fifoGroup_1_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_1_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[1]) begin
              fifoGroup_1_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[2]) begin
            fifoGroup_2_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[2]) begin
              fifoGroup_2_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[2]) begin
            fifoGroup_2_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[2]) begin
              fifoGroup_2_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_2_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[2]) begin
              fifoGroup_2_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[3]) begin
            fifoGroup_3_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[3]) begin
              fifoGroup_3_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[3]) begin
            fifoGroup_3_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[3]) begin
              fifoGroup_3_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_3_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[3]) begin
              fifoGroup_3_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[4]) begin
            fifoGroup_4_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[4]) begin
              fifoGroup_4_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[4]) begin
            fifoGroup_4_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[4]) begin
              fifoGroup_4_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_4_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[4]) begin
              fifoGroup_4_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[5]) begin
            fifoGroup_5_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[5]) begin
              fifoGroup_5_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[5]) begin
            fifoGroup_5_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[5]) begin
              fifoGroup_5_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_5_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[5]) begin
              fifoGroup_5_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[6]) begin
            fifoGroup_6_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[6]) begin
              fifoGroup_6_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[6]) begin
            fifoGroup_6_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[6]) begin
              fifoGroup_6_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_6_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[6]) begin
              fifoGroup_6_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[7]) begin
            fifoGroup_7_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[7]) begin
              fifoGroup_7_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[7]) begin
            fifoGroup_7_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[7]) begin
              fifoGroup_7_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_7_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[7]) begin
              fifoGroup_7_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[8]) begin
            fifoGroup_8_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[8]) begin
              fifoGroup_8_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[8]) begin
            fifoGroup_8_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[8]) begin
              fifoGroup_8_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_8_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[8]) begin
              fifoGroup_8_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[9]) begin
            fifoGroup_9_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[9]) begin
              fifoGroup_9_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[9]) begin
            fifoGroup_9_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[9]) begin
              fifoGroup_9_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_9_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[9]) begin
              fifoGroup_9_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[10]) begin
            fifoGroup_10_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[10]) begin
              fifoGroup_10_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[10]) begin
            fifoGroup_10_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[10]) begin
              fifoGroup_10_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_10_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[10]) begin
              fifoGroup_10_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[11]) begin
            fifoGroup_11_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[11]) begin
              fifoGroup_11_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[11]) begin
            fifoGroup_11_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[11]) begin
              fifoGroup_11_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_11_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[11]) begin
              fifoGroup_11_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[12]) begin
            fifoGroup_12_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[12]) begin
              fifoGroup_12_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[12]) begin
            fifoGroup_12_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[12]) begin
              fifoGroup_12_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_12_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[12]) begin
              fifoGroup_12_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[13]) begin
            fifoGroup_13_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[13]) begin
              fifoGroup_13_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[13]) begin
            fifoGroup_13_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[13]) begin
              fifoGroup_13_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_13_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[13]) begin
              fifoGroup_13_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[14]) begin
            fifoGroup_14_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[14]) begin
              fifoGroup_14_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[14]) begin
            fifoGroup_14_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[14]) begin
              fifoGroup_14_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_14_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[14]) begin
              fifoGroup_14_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[15]) begin
            fifoGroup_15_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[15]) begin
              fifoGroup_15_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[15]) begin
            fifoGroup_15_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[15]) begin
              fifoGroup_15_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_15_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[15]) begin
              fifoGroup_15_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[16]) begin
            fifoGroup_16_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[16]) begin
              fifoGroup_16_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[16]) begin
            fifoGroup_16_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[16]) begin
              fifoGroup_16_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_16_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[16]) begin
              fifoGroup_16_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[17]) begin
            fifoGroup_17_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[17]) begin
              fifoGroup_17_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[17]) begin
            fifoGroup_17_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[17]) begin
              fifoGroup_17_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_17_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[17]) begin
              fifoGroup_17_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[18]) begin
            fifoGroup_18_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[18]) begin
              fifoGroup_18_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[18]) begin
            fifoGroup_18_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[18]) begin
              fifoGroup_18_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_18_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[18]) begin
              fifoGroup_18_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[19]) begin
            fifoGroup_19_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[19]) begin
              fifoGroup_19_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[19]) begin
            fifoGroup_19_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[19]) begin
              fifoGroup_19_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_19_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[19]) begin
              fifoGroup_19_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[20]) begin
            fifoGroup_20_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[20]) begin
              fifoGroup_20_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[20]) begin
            fifoGroup_20_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[20]) begin
              fifoGroup_20_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_20_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[20]) begin
              fifoGroup_20_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[21]) begin
            fifoGroup_21_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[21]) begin
              fifoGroup_21_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[21]) begin
            fifoGroup_21_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[21]) begin
              fifoGroup_21_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_21_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[21]) begin
              fifoGroup_21_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[22]) begin
            fifoGroup_22_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[22]) begin
              fifoGroup_22_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[22]) begin
            fifoGroup_22_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[22]) begin
              fifoGroup_22_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_22_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[22]) begin
              fifoGroup_22_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[23]) begin
            fifoGroup_23_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[23]) begin
              fifoGroup_23_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[23]) begin
            fifoGroup_23_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[23]) begin
              fifoGroup_23_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_23_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[23]) begin
              fifoGroup_23_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[24]) begin
            fifoGroup_24_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[24]) begin
              fifoGroup_24_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[24]) begin
            fifoGroup_24_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[24]) begin
              fifoGroup_24_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_24_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[24]) begin
              fifoGroup_24_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[25]) begin
            fifoGroup_25_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[25]) begin
              fifoGroup_25_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[25]) begin
            fifoGroup_25_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[25]) begin
              fifoGroup_25_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_25_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[25]) begin
              fifoGroup_25_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[26]) begin
            fifoGroup_26_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[26]) begin
              fifoGroup_26_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[26]) begin
            fifoGroup_26_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[26]) begin
              fifoGroup_26_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_26_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[26]) begin
              fifoGroup_26_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[27]) begin
            fifoGroup_27_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[27]) begin
              fifoGroup_27_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[27]) begin
            fifoGroup_27_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[27]) begin
              fifoGroup_27_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_27_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[27]) begin
              fifoGroup_27_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[28]) begin
            fifoGroup_28_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[28]) begin
              fifoGroup_28_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[28]) begin
            fifoGroup_28_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[28]) begin
              fifoGroup_28_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_28_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[28]) begin
              fifoGroup_28_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[29]) begin
            fifoGroup_29_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[29]) begin
              fifoGroup_29_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[29]) begin
            fifoGroup_29_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[29]) begin
              fifoGroup_29_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_29_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[29]) begin
              fifoGroup_29_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[30]) begin
            fifoGroup_30_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[30]) begin
              fifoGroup_30_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[30]) begin
            fifoGroup_30_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[30]) begin
              fifoGroup_30_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_30_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[30]) begin
              fifoGroup_30_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[31]) begin
            fifoGroup_31_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[31]) begin
              fifoGroup_31_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[31]) begin
            fifoGroup_31_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[31]) begin
              fifoGroup_31_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_31_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[31]) begin
              fifoGroup_31_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[32]) begin
            fifoGroup_32_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[32]) begin
              fifoGroup_32_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[32]) begin
            fifoGroup_32_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[32]) begin
              fifoGroup_32_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_32_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[32]) begin
              fifoGroup_32_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[33]) begin
            fifoGroup_33_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[33]) begin
              fifoGroup_33_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[33]) begin
            fifoGroup_33_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[33]) begin
              fifoGroup_33_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_33_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[33]) begin
              fifoGroup_33_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[34]) begin
            fifoGroup_34_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[34]) begin
              fifoGroup_34_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[34]) begin
            fifoGroup_34_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[34]) begin
              fifoGroup_34_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_34_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[34]) begin
              fifoGroup_34_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[35]) begin
            fifoGroup_35_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[35]) begin
              fifoGroup_35_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[35]) begin
            fifoGroup_35_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[35]) begin
              fifoGroup_35_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_35_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[35]) begin
              fifoGroup_35_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[36]) begin
            fifoGroup_36_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[36]) begin
              fifoGroup_36_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[36]) begin
            fifoGroup_36_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[36]) begin
              fifoGroup_36_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_36_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[36]) begin
              fifoGroup_36_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[37]) begin
            fifoGroup_37_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[37]) begin
              fifoGroup_37_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[37]) begin
            fifoGroup_37_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[37]) begin
              fifoGroup_37_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_37_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[37]) begin
              fifoGroup_37_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[38]) begin
            fifoGroup_38_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[38]) begin
              fifoGroup_38_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[38]) begin
            fifoGroup_38_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[38]) begin
              fifoGroup_38_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_38_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[38]) begin
              fifoGroup_38_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[39]) begin
            fifoGroup_39_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[39]) begin
              fifoGroup_39_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[39]) begin
            fifoGroup_39_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[39]) begin
              fifoGroup_39_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_39_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[39]) begin
              fifoGroup_39_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[40]) begin
            fifoGroup_40_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[40]) begin
              fifoGroup_40_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[40]) begin
            fifoGroup_40_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[40]) begin
              fifoGroup_40_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_40_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[40]) begin
              fifoGroup_40_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[41]) begin
            fifoGroup_41_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[41]) begin
              fifoGroup_41_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[41]) begin
            fifoGroup_41_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[41]) begin
              fifoGroup_41_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_41_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[41]) begin
              fifoGroup_41_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[42]) begin
            fifoGroup_42_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[42]) begin
              fifoGroup_42_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[42]) begin
            fifoGroup_42_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[42]) begin
              fifoGroup_42_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_42_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[42]) begin
              fifoGroup_42_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[43]) begin
            fifoGroup_43_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[43]) begin
              fifoGroup_43_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[43]) begin
            fifoGroup_43_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[43]) begin
              fifoGroup_43_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_43_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[43]) begin
              fifoGroup_43_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[44]) begin
            fifoGroup_44_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[44]) begin
              fifoGroup_44_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[44]) begin
            fifoGroup_44_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[44]) begin
              fifoGroup_44_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_44_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[44]) begin
              fifoGroup_44_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[45]) begin
            fifoGroup_45_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[45]) begin
              fifoGroup_45_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[45]) begin
            fifoGroup_45_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[45]) begin
              fifoGroup_45_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_45_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[45]) begin
              fifoGroup_45_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[46]) begin
            fifoGroup_46_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[46]) begin
              fifoGroup_46_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[46]) begin
            fifoGroup_46_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[46]) begin
              fifoGroup_46_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_46_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[46]) begin
              fifoGroup_46_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[47]) begin
            fifoGroup_47_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[47]) begin
              fifoGroup_47_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[47]) begin
            fifoGroup_47_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[47]) begin
              fifoGroup_47_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_47_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[47]) begin
              fifoGroup_47_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[48]) begin
            fifoGroup_48_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[48]) begin
              fifoGroup_48_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[48]) begin
            fifoGroup_48_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[48]) begin
              fifoGroup_48_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_48_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[48]) begin
              fifoGroup_48_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[49]) begin
            fifoGroup_49_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[49]) begin
              fifoGroup_49_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[49]) begin
            fifoGroup_49_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[49]) begin
              fifoGroup_49_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_49_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[49]) begin
              fifoGroup_49_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[50]) begin
            fifoGroup_50_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[50]) begin
              fifoGroup_50_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[50]) begin
            fifoGroup_50_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[50]) begin
              fifoGroup_50_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_50_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[50]) begin
              fifoGroup_50_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[51]) begin
            fifoGroup_51_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[51]) begin
              fifoGroup_51_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[51]) begin
            fifoGroup_51_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[51]) begin
              fifoGroup_51_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_51_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[51]) begin
              fifoGroup_51_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[52]) begin
            fifoGroup_52_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[52]) begin
              fifoGroup_52_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[52]) begin
            fifoGroup_52_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[52]) begin
              fifoGroup_52_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_52_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[52]) begin
              fifoGroup_52_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[53]) begin
            fifoGroup_53_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[53]) begin
              fifoGroup_53_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[53]) begin
            fifoGroup_53_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[53]) begin
              fifoGroup_53_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_53_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[53]) begin
              fifoGroup_53_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[54]) begin
            fifoGroup_54_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[54]) begin
              fifoGroup_54_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[54]) begin
            fifoGroup_54_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[54]) begin
              fifoGroup_54_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_54_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[54]) begin
              fifoGroup_54_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[55]) begin
            fifoGroup_55_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[55]) begin
              fifoGroup_55_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[55]) begin
            fifoGroup_55_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[55]) begin
              fifoGroup_55_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_55_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[55]) begin
              fifoGroup_55_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[56]) begin
            fifoGroup_56_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[56]) begin
              fifoGroup_56_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[56]) begin
            fifoGroup_56_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[56]) begin
              fifoGroup_56_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_56_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[56]) begin
              fifoGroup_56_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[57]) begin
            fifoGroup_57_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[57]) begin
              fifoGroup_57_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[57]) begin
            fifoGroup_57_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[57]) begin
              fifoGroup_57_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_57_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[57]) begin
              fifoGroup_57_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[58]) begin
            fifoGroup_58_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[58]) begin
              fifoGroup_58_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[58]) begin
            fifoGroup_58_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[58]) begin
              fifoGroup_58_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_58_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[58]) begin
              fifoGroup_58_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[59]) begin
            fifoGroup_59_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[59]) begin
              fifoGroup_59_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[59]) begin
            fifoGroup_59_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[59]) begin
              fifoGroup_59_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_59_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[59]) begin
              fifoGroup_59_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[60]) begin
            fifoGroup_60_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[60]) begin
              fifoGroup_60_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[60]) begin
            fifoGroup_60_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[60]) begin
              fifoGroup_60_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_60_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[60]) begin
              fifoGroup_60_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[61]) begin
            fifoGroup_61_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[61]) begin
              fifoGroup_61_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[61]) begin
            fifoGroup_61_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[61]) begin
              fifoGroup_61_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_61_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[61]) begin
              fifoGroup_61_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[62]) begin
            fifoGroup_62_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[62]) begin
              fifoGroup_62_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[62]) begin
            fifoGroup_62_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[62]) begin
              fifoGroup_62_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_62_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[62]) begin
              fifoGroup_62_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[63]) begin
            fifoGroup_63_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[63]) begin
              fifoGroup_63_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[63]) begin
            fifoGroup_63_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[63]) begin
              fifoGroup_63_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_63_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[63]) begin
              fifoGroup_63_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_64_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[64]) begin
            fifoGroup_64_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[64]) begin
              fifoGroup_64_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_64_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[64]) begin
            fifoGroup_64_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[64]) begin
              fifoGroup_64_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_64_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[64]) begin
              fifoGroup_64_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_65_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[65]) begin
            fifoGroup_65_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[65]) begin
              fifoGroup_65_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_65_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[65]) begin
            fifoGroup_65_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[65]) begin
              fifoGroup_65_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_65_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[65]) begin
              fifoGroup_65_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_66_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[66]) begin
            fifoGroup_66_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[66]) begin
              fifoGroup_66_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_66_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[66]) begin
            fifoGroup_66_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[66]) begin
              fifoGroup_66_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_66_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[66]) begin
              fifoGroup_66_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_67_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[67]) begin
            fifoGroup_67_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[67]) begin
              fifoGroup_67_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_67_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[67]) begin
            fifoGroup_67_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[67]) begin
              fifoGroup_67_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_67_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[67]) begin
              fifoGroup_67_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_68_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[68]) begin
            fifoGroup_68_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[68]) begin
              fifoGroup_68_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_68_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[68]) begin
            fifoGroup_68_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[68]) begin
              fifoGroup_68_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_68_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[68]) begin
              fifoGroup_68_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_69_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[69]) begin
            fifoGroup_69_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[69]) begin
              fifoGroup_69_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_69_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[69]) begin
            fifoGroup_69_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[69]) begin
              fifoGroup_69_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_69_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[69]) begin
              fifoGroup_69_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_70_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[70]) begin
            fifoGroup_70_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[70]) begin
              fifoGroup_70_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_70_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[70]) begin
            fifoGroup_70_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[70]) begin
              fifoGroup_70_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_70_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[70]) begin
              fifoGroup_70_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_71_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[71]) begin
            fifoGroup_71_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[71]) begin
              fifoGroup_71_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_71_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[71]) begin
            fifoGroup_71_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[71]) begin
              fifoGroup_71_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_71_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[71]) begin
              fifoGroup_71_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_72_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[72]) begin
            fifoGroup_72_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[72]) begin
              fifoGroup_72_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_72_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[72]) begin
            fifoGroup_72_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[72]) begin
              fifoGroup_72_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_72_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[72]) begin
              fifoGroup_72_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_73_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[73]) begin
            fifoGroup_73_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[73]) begin
              fifoGroup_73_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_73_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[73]) begin
            fifoGroup_73_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[73]) begin
              fifoGroup_73_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_73_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[73]) begin
              fifoGroup_73_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_74_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[74]) begin
            fifoGroup_74_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[74]) begin
              fifoGroup_74_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_74_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[74]) begin
            fifoGroup_74_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[74]) begin
              fifoGroup_74_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_74_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[74]) begin
              fifoGroup_74_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_75_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[75]) begin
            fifoGroup_75_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[75]) begin
              fifoGroup_75_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_75_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[75]) begin
            fifoGroup_75_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[75]) begin
              fifoGroup_75_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_75_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[75]) begin
              fifoGroup_75_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_76_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[76]) begin
            fifoGroup_76_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[76]) begin
              fifoGroup_76_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_76_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[76]) begin
            fifoGroup_76_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[76]) begin
              fifoGroup_76_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_76_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[76]) begin
              fifoGroup_76_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_77_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[77]) begin
            fifoGroup_77_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[77]) begin
              fifoGroup_77_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_77_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[77]) begin
            fifoGroup_77_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[77]) begin
              fifoGroup_77_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_77_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[77]) begin
              fifoGroup_77_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_78_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[78]) begin
            fifoGroup_78_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[78]) begin
              fifoGroup_78_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_78_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[78]) begin
            fifoGroup_78_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[78]) begin
              fifoGroup_78_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_78_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[78]) begin
              fifoGroup_78_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_79_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[79]) begin
            fifoGroup_79_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[79]) begin
              fifoGroup_79_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_79_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[79]) begin
            fifoGroup_79_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[79]) begin
              fifoGroup_79_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_79_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[79]) begin
              fifoGroup_79_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_80_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[80]) begin
            fifoGroup_80_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[80]) begin
              fifoGroup_80_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_80_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[80]) begin
            fifoGroup_80_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[80]) begin
              fifoGroup_80_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_80_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[80]) begin
              fifoGroup_80_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_81_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[81]) begin
            fifoGroup_81_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[81]) begin
              fifoGroup_81_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_81_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[81]) begin
            fifoGroup_81_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[81]) begin
              fifoGroup_81_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_81_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[81]) begin
              fifoGroup_81_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_82_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[82]) begin
            fifoGroup_82_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[82]) begin
              fifoGroup_82_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_82_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[82]) begin
            fifoGroup_82_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[82]) begin
              fifoGroup_82_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_82_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[82]) begin
              fifoGroup_82_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_83_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[83]) begin
            fifoGroup_83_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[83]) begin
              fifoGroup_83_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_83_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[83]) begin
            fifoGroup_83_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[83]) begin
              fifoGroup_83_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_83_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[83]) begin
              fifoGroup_83_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_84_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[84]) begin
            fifoGroup_84_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[84]) begin
              fifoGroup_84_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_84_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[84]) begin
            fifoGroup_84_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[84]) begin
              fifoGroup_84_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_84_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[84]) begin
              fifoGroup_84_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_85_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[85]) begin
            fifoGroup_85_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[85]) begin
              fifoGroup_85_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_85_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[85]) begin
            fifoGroup_85_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[85]) begin
              fifoGroup_85_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_85_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[85]) begin
              fifoGroup_85_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_86_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[86]) begin
            fifoGroup_86_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[86]) begin
              fifoGroup_86_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_86_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[86]) begin
            fifoGroup_86_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[86]) begin
              fifoGroup_86_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_86_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[86]) begin
              fifoGroup_86_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_87_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[87]) begin
            fifoGroup_87_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[87]) begin
              fifoGroup_87_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_87_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[87]) begin
            fifoGroup_87_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[87]) begin
              fifoGroup_87_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_87_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[87]) begin
              fifoGroup_87_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_88_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[88]) begin
            fifoGroup_88_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[88]) begin
              fifoGroup_88_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_88_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[88]) begin
            fifoGroup_88_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[88]) begin
              fifoGroup_88_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_88_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[88]) begin
              fifoGroup_88_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_89_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[89]) begin
            fifoGroup_89_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[89]) begin
              fifoGroup_89_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_89_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[89]) begin
            fifoGroup_89_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[89]) begin
              fifoGroup_89_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_89_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[89]) begin
              fifoGroup_89_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_90_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[90]) begin
            fifoGroup_90_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[90]) begin
              fifoGroup_90_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_90_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[90]) begin
            fifoGroup_90_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[90]) begin
              fifoGroup_90_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_90_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[90]) begin
              fifoGroup_90_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_91_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[91]) begin
            fifoGroup_91_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[91]) begin
              fifoGroup_91_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_91_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[91]) begin
            fifoGroup_91_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[91]) begin
              fifoGroup_91_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_91_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[91]) begin
              fifoGroup_91_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_92_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[92]) begin
            fifoGroup_92_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[92]) begin
              fifoGroup_92_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_92_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[92]) begin
            fifoGroup_92_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[92]) begin
              fifoGroup_92_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_92_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[92]) begin
              fifoGroup_92_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_93_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[93]) begin
            fifoGroup_93_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[93]) begin
              fifoGroup_93_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_93_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[93]) begin
            fifoGroup_93_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[93]) begin
              fifoGroup_93_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_93_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[93]) begin
              fifoGroup_93_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_94_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[94]) begin
            fifoGroup_94_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[94]) begin
              fifoGroup_94_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_94_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[94]) begin
            fifoGroup_94_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[94]) begin
              fifoGroup_94_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_94_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[94]) begin
              fifoGroup_94_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_95_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[95]) begin
            fifoGroup_95_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[95]) begin
              fifoGroup_95_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_95_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[95]) begin
            fifoGroup_95_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[95]) begin
              fifoGroup_95_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_95_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[95]) begin
              fifoGroup_95_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_96_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[96]) begin
            fifoGroup_96_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[96]) begin
              fifoGroup_96_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_96_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[96]) begin
            fifoGroup_96_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[96]) begin
              fifoGroup_96_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_96_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[96]) begin
              fifoGroup_96_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_97_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[97]) begin
            fifoGroup_97_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[97]) begin
              fifoGroup_97_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_97_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[97]) begin
            fifoGroup_97_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[97]) begin
              fifoGroup_97_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_97_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[97]) begin
              fifoGroup_97_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_98_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[98]) begin
            fifoGroup_98_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[98]) begin
              fifoGroup_98_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_98_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[98]) begin
            fifoGroup_98_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[98]) begin
              fifoGroup_98_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_98_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[98]) begin
              fifoGroup_98_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_99_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[99]) begin
            fifoGroup_99_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[99]) begin
              fifoGroup_99_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_99_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[99]) begin
            fifoGroup_99_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[99]) begin
              fifoGroup_99_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_99_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[99]) begin
              fifoGroup_99_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_100_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[100]) begin
            fifoGroup_100_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[100]) begin
              fifoGroup_100_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_100_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[100]) begin
            fifoGroup_100_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[100]) begin
              fifoGroup_100_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_100_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[100]) begin
              fifoGroup_100_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_101_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[101]) begin
            fifoGroup_101_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[101]) begin
              fifoGroup_101_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_101_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[101]) begin
            fifoGroup_101_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[101]) begin
              fifoGroup_101_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_101_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[101]) begin
              fifoGroup_101_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_102_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[102]) begin
            fifoGroup_102_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[102]) begin
              fifoGroup_102_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_102_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[102]) begin
            fifoGroup_102_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[102]) begin
              fifoGroup_102_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_102_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[102]) begin
              fifoGroup_102_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_103_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[103]) begin
            fifoGroup_103_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[103]) begin
              fifoGroup_103_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_103_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[103]) begin
            fifoGroup_103_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[103]) begin
              fifoGroup_103_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_103_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[103]) begin
              fifoGroup_103_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_104_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[104]) begin
            fifoGroup_104_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[104]) begin
              fifoGroup_104_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_104_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[104]) begin
            fifoGroup_104_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[104]) begin
              fifoGroup_104_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_104_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[104]) begin
              fifoGroup_104_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_105_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[105]) begin
            fifoGroup_105_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[105]) begin
              fifoGroup_105_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_105_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[105]) begin
            fifoGroup_105_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[105]) begin
              fifoGroup_105_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_105_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[105]) begin
              fifoGroup_105_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_106_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[106]) begin
            fifoGroup_106_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[106]) begin
              fifoGroup_106_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_106_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[106]) begin
            fifoGroup_106_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[106]) begin
              fifoGroup_106_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_106_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[106]) begin
              fifoGroup_106_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_107_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[107]) begin
            fifoGroup_107_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[107]) begin
              fifoGroup_107_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_107_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[107]) begin
            fifoGroup_107_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[107]) begin
              fifoGroup_107_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_107_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[107]) begin
              fifoGroup_107_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_108_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[108]) begin
            fifoGroup_108_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[108]) begin
              fifoGroup_108_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_108_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[108]) begin
            fifoGroup_108_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[108]) begin
              fifoGroup_108_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_108_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[108]) begin
              fifoGroup_108_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_109_io_push_valid = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_1[109]) begin
            fifoGroup_109_io_push_valid = _zz_io_push_valid;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_19[109]) begin
              fifoGroup_109_io_push_valid = _zz_io_push_valid_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_109_io_push_payload = 32'h0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l204) begin
          if(_zz_2[109]) begin
            fifoGroup_109_io_push_payload = _zz_io_push_payload;
          end
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l336) begin
          if(when_ArraySlice_l337) begin
            if(_zz_20[109]) begin
              fifoGroup_109_io_push_payload = _zz_io_push_payload_1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifoGroup_109_io_pop_ready = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l376) begin
          if(when_ArraySlice_l377) begin
            if(_zz_3[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready;
            end
          end
        end
        if(when_ArraySlice_l376_1) begin
          if(when_ArraySlice_l377_1) begin
            if(_zz_4[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_1;
            end
          end
        end
        if(when_ArraySlice_l376_2) begin
          if(when_ArraySlice_l377_2) begin
            if(_zz_5[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_2;
            end
          end
        end
        if(when_ArraySlice_l376_3) begin
          if(when_ArraySlice_l377_3) begin
            if(_zz_6[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_3;
            end
          end
        end
        if(when_ArraySlice_l376_4) begin
          if(when_ArraySlice_l377_4) begin
            if(_zz_7[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_4;
            end
          end
        end
        if(when_ArraySlice_l376_5) begin
          if(when_ArraySlice_l377_5) begin
            if(_zz_8[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_5;
            end
          end
        end
        if(when_ArraySlice_l376_6) begin
          if(when_ArraySlice_l377_6) begin
            if(_zz_9[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_6;
            end
          end
        end
        if(when_ArraySlice_l376_7) begin
          if(when_ArraySlice_l377_7) begin
            if(_zz_10[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_7;
            end
          end
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l233) begin
          if(when_ArraySlice_l234) begin
            if(_zz_11[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_8;
            end
          end
        end
        if(when_ArraySlice_l233_1) begin
          if(when_ArraySlice_l234_1) begin
            if(_zz_12[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_9;
            end
          end
        end
        if(when_ArraySlice_l233_2) begin
          if(when_ArraySlice_l234_2) begin
            if(_zz_13[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_10;
            end
          end
        end
        if(when_ArraySlice_l233_3) begin
          if(when_ArraySlice_l234_3) begin
            if(_zz_14[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_11;
            end
          end
        end
        if(when_ArraySlice_l233_4) begin
          if(when_ArraySlice_l234_4) begin
            if(_zz_15[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_12;
            end
          end
        end
        if(when_ArraySlice_l233_5) begin
          if(when_ArraySlice_l234_5) begin
            if(_zz_16[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_13;
            end
          end
        end
        if(when_ArraySlice_l233_6) begin
          if(when_ArraySlice_l234_6) begin
            if(_zz_17[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_14;
            end
          end
        end
        if(when_ArraySlice_l233_7) begin
          if(when_ArraySlice_l234_7) begin
            if(_zz_18[109]) begin
              fifoGroup_109_io_pop_ready = _zz_io_pop_ready_15;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign arraySliceStateMachine_wantExit = 1'b0;
  always @(*) begin
    arraySliceStateMachine_wantStart = 1'b0;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
      end
      default : begin
        arraySliceStateMachine_wantStart = 1'b1;
      end
    endcase
  end

  assign arraySliceStateMachine_wantKill = 1'b0;
  always @(*) begin
    arraySliceStateMachine_stateNext = arraySliceStateMachine_stateReg;
    case(arraySliceStateMachine_stateReg)
      arraySliceStateMachine_enumDef_writeDataOnly : begin
        if(when_ArraySlice_l216) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readWriteData;
        end
      end
      arraySliceStateMachine_enumDef_readDataOnly : begin
        if(when_ArraySlice_l478) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readWriteData;
        end
      end
      arraySliceStateMachine_enumDef_readWriteData : begin
        if(when_ArraySlice_l357) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_writeDataOnly;
        end
        if(when_ArraySlice_l361) begin
          arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_readDataOnly;
        end
      end
      default : begin
      end
    endcase
    if(arraySliceStateMachine_wantStart) begin
      arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_writeDataOnly;
    end
    if(arraySliceStateMachine_wantKill) begin
      arraySliceStateMachine_stateNext = arraySliceStateMachine_enumDef_BOOT;
    end
  end

  assign when_ArraySlice_l204 = (_zz_when_ArraySlice_l204 < hReg);
  assign _zz_1 = ({127'd0,1'b1} <<< selectWriteFifo);
  assign _zz_2 = ({127'd0,1'b1} <<< selectWriteFifo);
  assign _zz_io_push_valid = inputStreamArrayData_valid;
  assign _zz_io_push_payload = inputStreamArrayData_payload;
  assign inputStreamArrayData_fire = (inputStreamArrayData_valid && inputStreamArrayData_ready);
  assign when_ArraySlice_l208 = ((_zz_when_ArraySlice_l208 == _zz_when_ArraySlice_l208_1) && inputStreamArrayData_fire);
  assign when_ArraySlice_l209 = (selectWriteFifo == _zz_when_ArraySlice_l209);
  always @(*) begin
    debug_0 = 1'b0;
    if(when_ArraySlice_l158) begin
      if(when_ArraySlice_l159) begin
        debug_0 = 1'b1;
      end else begin
        debug_0 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166) begin
        debug_0 = 1'b1;
      end else begin
        debug_0 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1 = 1'b0;
    if(when_ArraySlice_l158_1) begin
      if(when_ArraySlice_l159_1) begin
        debug_1 = 1'b1;
      end else begin
        debug_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_1) begin
        debug_1 = 1'b1;
      end else begin
        debug_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2 = 1'b0;
    if(when_ArraySlice_l158_2) begin
      if(when_ArraySlice_l159_2) begin
        debug_2 = 1'b1;
      end else begin
        debug_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_2) begin
        debug_2 = 1'b1;
      end else begin
        debug_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3 = 1'b0;
    if(when_ArraySlice_l158_3) begin
      if(when_ArraySlice_l159_3) begin
        debug_3 = 1'b1;
      end else begin
        debug_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_3) begin
        debug_3 = 1'b1;
      end else begin
        debug_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4 = 1'b0;
    if(when_ArraySlice_l158_4) begin
      if(when_ArraySlice_l159_4) begin
        debug_4 = 1'b1;
      end else begin
        debug_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_4) begin
        debug_4 = 1'b1;
      end else begin
        debug_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5 = 1'b0;
    if(when_ArraySlice_l158_5) begin
      if(when_ArraySlice_l159_5) begin
        debug_5 = 1'b1;
      end else begin
        debug_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_5) begin
        debug_5 = 1'b1;
      end else begin
        debug_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6 = 1'b0;
    if(when_ArraySlice_l158_6) begin
      if(when_ArraySlice_l159_6) begin
        debug_6 = 1'b1;
      end else begin
        debug_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_6) begin
        debug_6 = 1'b1;
      end else begin
        debug_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7 = 1'b0;
    if(when_ArraySlice_l158_7) begin
      if(when_ArraySlice_l159_7) begin
        debug_7 = 1'b1;
      end else begin
        debug_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_7) begin
        debug_7 = 1'b1;
      end else begin
        debug_7 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158 = (_zz_when_ArraySlice_l158 <= _zz_when_ArraySlice_l158_3);
  assign when_ArraySlice_l159 = (_zz_when_ArraySlice_l159 <= _zz_when_ArraySlice_l159_1);
  assign _zz_realValue_0 = (_zz__zz_realValue_0 % _zz__zz_realValue_0_1);
  assign when_ArraySlice_l110 = (_zz_realValue_0 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110) begin
      realValue_0 = (_zz_realValue_0_416 - _zz_realValue_0);
    end else begin
      realValue_0 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166 = (_zz_when_ArraySlice_l166 <= _zz_when_ArraySlice_l166_1);
  assign when_ArraySlice_l158_1 = (_zz_when_ArraySlice_l158_1_1 <= _zz_when_ArraySlice_l158_1_4);
  assign when_ArraySlice_l159_1 = (_zz_when_ArraySlice_l159_1_1 <= _zz_when_ArraySlice_l159_1_3);
  assign _zz_realValue_0_1 = (_zz__zz_realValue_0_1_1 % _zz__zz_realValue_0_1_2);
  assign when_ArraySlice_l110_1 = (_zz_realValue_0_1 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_1) begin
      realValue_0_1 = (_zz_realValue_0_1_1 - _zz_realValue_0_1);
    end else begin
      realValue_0_1 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_1 = (_zz_when_ArraySlice_l166_1_1 <= _zz_when_ArraySlice_l166_1_3);
  assign when_ArraySlice_l158_2 = (_zz_when_ArraySlice_l158_2_1 <= _zz_when_ArraySlice_l158_2_4);
  assign when_ArraySlice_l159_2 = (_zz_when_ArraySlice_l159_2_1 <= _zz_when_ArraySlice_l159_2_3);
  assign _zz_realValue_0_2 = (_zz__zz_realValue_0_2 % _zz__zz_realValue_0_2_1);
  assign when_ArraySlice_l110_2 = (_zz_realValue_0_2 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_2) begin
      realValue_0_2 = (_zz_realValue_0_2_1 - _zz_realValue_0_2);
    end else begin
      realValue_0_2 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_2 = (_zz_when_ArraySlice_l166_2_1 <= _zz_when_ArraySlice_l166_2_3);
  assign when_ArraySlice_l158_3 = (_zz_when_ArraySlice_l158_3_1 <= _zz_when_ArraySlice_l158_3_4);
  assign when_ArraySlice_l159_3 = (_zz_when_ArraySlice_l159_3_1 <= _zz_when_ArraySlice_l159_3_3);
  assign _zz_realValue_0_3 = (_zz__zz_realValue_0_3 % _zz__zz_realValue_0_3_1);
  assign when_ArraySlice_l110_3 = (_zz_realValue_0_3 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_3) begin
      realValue_0_3 = (_zz_realValue_0_3_1 - _zz_realValue_0_3);
    end else begin
      realValue_0_3 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_3 = (_zz_when_ArraySlice_l166_3_1 <= _zz_when_ArraySlice_l166_3_3);
  assign when_ArraySlice_l158_4 = (_zz_when_ArraySlice_l158_4 <= _zz_when_ArraySlice_l158_4_3);
  assign when_ArraySlice_l159_4 = (_zz_when_ArraySlice_l159_4_1 <= _zz_when_ArraySlice_l159_4_3);
  assign _zz_realValue_0_4 = (_zz__zz_realValue_0_4 % _zz__zz_realValue_0_4_1);
  assign when_ArraySlice_l110_4 = (_zz_realValue_0_4 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_4) begin
      realValue_0_4 = (_zz_realValue_0_4_1 - _zz_realValue_0_4);
    end else begin
      realValue_0_4 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_4 = (_zz_when_ArraySlice_l166_4_1 <= _zz_when_ArraySlice_l166_4_3);
  assign when_ArraySlice_l158_5 = (_zz_when_ArraySlice_l158_5 <= _zz_when_ArraySlice_l158_5_3);
  assign when_ArraySlice_l159_5 = (_zz_when_ArraySlice_l159_5_1 <= _zz_when_ArraySlice_l159_5_3);
  assign _zz_realValue_0_5 = (_zz__zz_realValue_0_5 % _zz__zz_realValue_0_5_1);
  assign when_ArraySlice_l110_5 = (_zz_realValue_0_5 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_5) begin
      realValue_0_5 = (_zz_realValue_0_5_1 - _zz_realValue_0_5);
    end else begin
      realValue_0_5 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_5 = (_zz_when_ArraySlice_l166_5_1 <= _zz_when_ArraySlice_l166_5_3);
  assign when_ArraySlice_l158_6 = (_zz_when_ArraySlice_l158_6 <= _zz_when_ArraySlice_l158_6_3);
  assign when_ArraySlice_l159_6 = (_zz_when_ArraySlice_l159_6 <= _zz_when_ArraySlice_l159_6_2);
  assign _zz_realValue_0_6 = (_zz__zz_realValue_0_6 % _zz__zz_realValue_0_6_1);
  assign when_ArraySlice_l110_6 = (_zz_realValue_0_6 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_6) begin
      realValue_0_6 = (_zz_realValue_0_6_1 - _zz_realValue_0_6);
    end else begin
      realValue_0_6 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_6 = (_zz_when_ArraySlice_l166_6_1 <= _zz_when_ArraySlice_l166_6_3);
  assign when_ArraySlice_l158_7 = (_zz_when_ArraySlice_l158_7 <= _zz_when_ArraySlice_l158_7_3);
  assign when_ArraySlice_l159_7 = (_zz_when_ArraySlice_l159_7 <= _zz_when_ArraySlice_l159_7_2);
  assign _zz_realValue_0_7 = (_zz__zz_realValue_0_7 % _zz__zz_realValue_0_7_1);
  assign when_ArraySlice_l110_7 = (_zz_realValue_0_7 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_7) begin
      realValue_0_7 = (_zz_realValue_0_7_1 - _zz_realValue_0_7);
    end else begin
      realValue_0_7 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_7 = (_zz_when_ArraySlice_l166_7 <= _zz_when_ArraySlice_l166_7_2);
  assign when_ArraySlice_l216 = ((((((((debug_0 == 1'b1) && (debug_1 == 1'b1)) && (debug_2 == 1'b1)) && (debug_3 == 1'b1)) && (debug_4 == 1'b1)) && (debug_5 == 1'b1)) && (debug_6 == 1'b1)) && (debug_7 == 1'b1));
  assign when_ArraySlice_l222 = (! allowPadding_0);
  assign when_ArraySlice_l222_1 = (! allowPadding_1);
  assign when_ArraySlice_l222_2 = (! allowPadding_2);
  assign when_ArraySlice_l222_3 = (! allowPadding_3);
  assign when_ArraySlice_l222_4 = (! allowPadding_4);
  assign when_ArraySlice_l222_5 = (! allowPadding_5);
  assign when_ArraySlice_l222_6 = (! allowPadding_6);
  assign when_ArraySlice_l222_7 = (! allowPadding_7);
  assign when_ArraySlice_l376 = (_zz_when_ArraySlice_l376 < _zz_when_ArraySlice_l376_3);
  assign when_ArraySlice_l377 = ((! holdReadOp_0) && (_zz_when_ArraySlice_l377 != 7'h0));
  assign _zz_outputStreamArrayData_0_valid = (selectReadFifo_0 + _zz__zz_outputStreamArrayData_0_valid);
  assign _zz_3 = ({127'd0,1'b1} <<< _zz__zz_3);
  assign _zz_io_pop_ready = outputStreamArrayData_0_ready;
  assign when_ArraySlice_l382 = (! holdReadOp_0);
  assign outputStreamArrayData_0_fire = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l383 = ((7'h01 < _zz_when_ArraySlice_l383) && outputStreamArrayData_0_fire);
  assign when_ArraySlice_l384 = (handshakeTimes_0_value == _zz_when_ArraySlice_l384);
  assign when_ArraySlice_l387 = (_zz_when_ArraySlice_l387 == 13'h0);
  assign outputStreamArrayData_0_fire_1 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l392 = ((_zz_when_ArraySlice_l392 == 7'h01) && outputStreamArrayData_0_fire_1);
  assign when_ArraySlice_l393 = (handshakeTimes_0_value == _zz_when_ArraySlice_l393);
  assign _zz_realValue1_0 = (_zz__zz_realValue1_0 % _zz__zz_realValue1_0_1);
  assign when_ArraySlice_l95 = (_zz_realValue1_0 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95) begin
      realValue1_0 = (_zz_realValue1_0_48 - _zz_realValue1_0);
    end else begin
      realValue1_0 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395 = (_zz_when_ArraySlice_l395 < _zz_when_ArraySlice_l395_2);
  always @(*) begin
    debug_0_1 = 1'b0;
    if(when_ArraySlice_l158_8) begin
      if(when_ArraySlice_l159_8) begin
        debug_0_1 = 1'b1;
      end else begin
        debug_0_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_8) begin
        debug_0_1 = 1'b1;
      end else begin
        debug_0_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_1 = 1'b0;
    if(when_ArraySlice_l158_9) begin
      if(when_ArraySlice_l159_9) begin
        debug_1_1 = 1'b1;
      end else begin
        debug_1_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_9) begin
        debug_1_1 = 1'b1;
      end else begin
        debug_1_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_1 = 1'b0;
    if(when_ArraySlice_l158_10) begin
      if(when_ArraySlice_l159_10) begin
        debug_2_1 = 1'b1;
      end else begin
        debug_2_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_10) begin
        debug_2_1 = 1'b1;
      end else begin
        debug_2_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_1 = 1'b0;
    if(when_ArraySlice_l158_11) begin
      if(when_ArraySlice_l159_11) begin
        debug_3_1 = 1'b1;
      end else begin
        debug_3_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_11) begin
        debug_3_1 = 1'b1;
      end else begin
        debug_3_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_1 = 1'b0;
    if(when_ArraySlice_l158_12) begin
      if(when_ArraySlice_l159_12) begin
        debug_4_1 = 1'b1;
      end else begin
        debug_4_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_12) begin
        debug_4_1 = 1'b1;
      end else begin
        debug_4_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_1 = 1'b0;
    if(when_ArraySlice_l158_13) begin
      if(when_ArraySlice_l159_13) begin
        debug_5_1 = 1'b1;
      end else begin
        debug_5_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_13) begin
        debug_5_1 = 1'b1;
      end else begin
        debug_5_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_1 = 1'b0;
    if(when_ArraySlice_l158_14) begin
      if(when_ArraySlice_l159_14) begin
        debug_6_1 = 1'b1;
      end else begin
        debug_6_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_14) begin
        debug_6_1 = 1'b1;
      end else begin
        debug_6_1 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_1 = 1'b0;
    if(when_ArraySlice_l158_15) begin
      if(when_ArraySlice_l159_15) begin
        debug_7_1 = 1'b1;
      end else begin
        debug_7_1 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_15) begin
        debug_7_1 = 1'b1;
      end else begin
        debug_7_1 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_8 = (_zz_when_ArraySlice_l158_8 <= _zz_when_ArraySlice_l158_8_3);
  assign when_ArraySlice_l159_8 = (_zz_when_ArraySlice_l159_8 <= _zz_when_ArraySlice_l159_8_1);
  assign _zz_realValue_0_8 = (_zz__zz_realValue_0_8 % _zz__zz_realValue_0_8_1);
  assign when_ArraySlice_l110_8 = (_zz_realValue_0_8 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_8) begin
      realValue_0_8 = (_zz_realValue_0_8_1 - _zz_realValue_0_8);
    end else begin
      realValue_0_8 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_8 = (_zz_when_ArraySlice_l166_8 <= _zz_when_ArraySlice_l166_8_1);
  assign when_ArraySlice_l158_9 = (_zz_when_ArraySlice_l158_9 <= _zz_when_ArraySlice_l158_9_3);
  assign when_ArraySlice_l159_9 = (_zz_when_ArraySlice_l159_9 <= _zz_when_ArraySlice_l159_9_2);
  assign _zz_realValue_0_9 = (_zz__zz_realValue_0_9 % _zz__zz_realValue_0_9_1);
  assign when_ArraySlice_l110_9 = (_zz_realValue_0_9 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_9) begin
      realValue_0_9 = (_zz_realValue_0_9_1 - _zz_realValue_0_9);
    end else begin
      realValue_0_9 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_9 = (_zz_when_ArraySlice_l166_9 <= _zz_when_ArraySlice_l166_9_2);
  assign when_ArraySlice_l158_10 = (_zz_when_ArraySlice_l158_10 <= _zz_when_ArraySlice_l158_10_3);
  assign when_ArraySlice_l159_10 = (_zz_when_ArraySlice_l159_10 <= _zz_when_ArraySlice_l159_10_2);
  assign _zz_realValue_0_10 = (_zz__zz_realValue_0_10 % _zz__zz_realValue_0_10_1);
  assign when_ArraySlice_l110_10 = (_zz_realValue_0_10 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_10) begin
      realValue_0_10 = (_zz_realValue_0_10_1 - _zz_realValue_0_10);
    end else begin
      realValue_0_10 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_10 = (_zz_when_ArraySlice_l166_10 <= _zz_when_ArraySlice_l166_10_2);
  assign when_ArraySlice_l158_11 = (_zz_when_ArraySlice_l158_11 <= _zz_when_ArraySlice_l158_11_3);
  assign when_ArraySlice_l159_11 = (_zz_when_ArraySlice_l159_11 <= _zz_when_ArraySlice_l159_11_2);
  assign _zz_realValue_0_11 = (_zz__zz_realValue_0_11 % _zz__zz_realValue_0_11_1);
  assign when_ArraySlice_l110_11 = (_zz_realValue_0_11 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_11) begin
      realValue_0_11 = (_zz_realValue_0_11_1 - _zz_realValue_0_11);
    end else begin
      realValue_0_11 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_11 = (_zz_when_ArraySlice_l166_11 <= _zz_when_ArraySlice_l166_11_2);
  assign when_ArraySlice_l158_12 = (_zz_when_ArraySlice_l158_12 <= _zz_when_ArraySlice_l158_12_3);
  assign when_ArraySlice_l159_12 = (_zz_when_ArraySlice_l159_12 <= _zz_when_ArraySlice_l159_12_2);
  assign _zz_realValue_0_12 = (_zz__zz_realValue_0_12 % _zz__zz_realValue_0_12_1);
  assign when_ArraySlice_l110_12 = (_zz_realValue_0_12 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_12) begin
      realValue_0_12 = (_zz_realValue_0_12_1 - _zz_realValue_0_12);
    end else begin
      realValue_0_12 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_12 = (_zz_when_ArraySlice_l166_12 <= _zz_when_ArraySlice_l166_12_2);
  assign when_ArraySlice_l158_13 = (_zz_when_ArraySlice_l158_13 <= _zz_when_ArraySlice_l158_13_3);
  assign when_ArraySlice_l159_13 = (_zz_when_ArraySlice_l159_13 <= _zz_when_ArraySlice_l159_13_2);
  assign _zz_realValue_0_13 = (_zz__zz_realValue_0_13 % _zz__zz_realValue_0_13_1);
  assign when_ArraySlice_l110_13 = (_zz_realValue_0_13 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_13) begin
      realValue_0_13 = (_zz_realValue_0_13_1 - _zz_realValue_0_13);
    end else begin
      realValue_0_13 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_13 = (_zz_when_ArraySlice_l166_13 <= _zz_when_ArraySlice_l166_13_2);
  assign when_ArraySlice_l158_14 = (_zz_when_ArraySlice_l158_14 <= _zz_when_ArraySlice_l158_14_3);
  assign when_ArraySlice_l159_14 = (_zz_when_ArraySlice_l159_14 <= _zz_when_ArraySlice_l159_14_2);
  assign _zz_realValue_0_14 = (_zz__zz_realValue_0_14 % _zz__zz_realValue_0_14_1);
  assign when_ArraySlice_l110_14 = (_zz_realValue_0_14 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_14) begin
      realValue_0_14 = (_zz_realValue_0_14_1 - _zz_realValue_0_14);
    end else begin
      realValue_0_14 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_14 = (_zz_when_ArraySlice_l166_14 <= _zz_when_ArraySlice_l166_14_2);
  assign when_ArraySlice_l158_15 = (_zz_when_ArraySlice_l158_15 <= _zz_when_ArraySlice_l158_15_3);
  assign when_ArraySlice_l159_15 = (_zz_when_ArraySlice_l159_15 <= _zz_when_ArraySlice_l159_15_2);
  assign _zz_realValue_0_15 = (_zz__zz_realValue_0_15 % _zz__zz_realValue_0_15_1);
  assign when_ArraySlice_l110_15 = (_zz_realValue_0_15 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_15) begin
      realValue_0_15 = (_zz_realValue_0_15_1 - _zz_realValue_0_15);
    end else begin
      realValue_0_15 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_15 = (_zz_when_ArraySlice_l166_15 <= _zz_when_ArraySlice_l166_15_2);
  assign when_ArraySlice_l400 = (! (((((_zz_when_ArraySlice_l400 && _zz_when_ArraySlice_l400_3) && (holdReadOp_5 == _zz_when_ArraySlice_l400_4)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && ((((_zz_when_ArraySlice_l400_5 && _zz_when_ArraySlice_l400_8) && (debug_5_1 == _zz_when_ArraySlice_l400_9)) && (debug_6_1 == 1'b1)) && (debug_7_1 == 1'b1))));
  assign when_ArraySlice_l403 = (_zz_when_ArraySlice_l403 <= _zz_when_ArraySlice_l403_1);
  assign when_ArraySlice_l406 = (_zz_when_ArraySlice_l406 <= _zz_when_ArraySlice_l406_1);
  assign when_ArraySlice_l413 = (_zz_when_ArraySlice_l413 == 13'h0);
  assign when_ArraySlice_l417 = (_zz_when_ArraySlice_l417 == 7'h0);
  assign outputStreamArrayData_0_fire_2 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l418 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l418) && outputStreamArrayData_0_fire_2);
  assign _zz_realValue1_0_1 = (_zz__zz_realValue1_0_1_1 % _zz__zz_realValue1_0_1_2);
  assign when_ArraySlice_l95_1 = (_zz_realValue1_0_1 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_1) begin
      realValue1_0_1 = (_zz_realValue1_0_1_1 - _zz_realValue1_0_1);
    end else begin
      realValue1_0_1 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420 = (_zz_when_ArraySlice_l420 < _zz_when_ArraySlice_l420_2);
  always @(*) begin
    debug_0_2 = 1'b0;
    if(when_ArraySlice_l158_16) begin
      if(when_ArraySlice_l159_16) begin
        debug_0_2 = 1'b1;
      end else begin
        debug_0_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_16) begin
        debug_0_2 = 1'b1;
      end else begin
        debug_0_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_2 = 1'b0;
    if(when_ArraySlice_l158_17) begin
      if(when_ArraySlice_l159_17) begin
        debug_1_2 = 1'b1;
      end else begin
        debug_1_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_17) begin
        debug_1_2 = 1'b1;
      end else begin
        debug_1_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_2 = 1'b0;
    if(when_ArraySlice_l158_18) begin
      if(when_ArraySlice_l159_18) begin
        debug_2_2 = 1'b1;
      end else begin
        debug_2_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_18) begin
        debug_2_2 = 1'b1;
      end else begin
        debug_2_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_2 = 1'b0;
    if(when_ArraySlice_l158_19) begin
      if(when_ArraySlice_l159_19) begin
        debug_3_2 = 1'b1;
      end else begin
        debug_3_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_19) begin
        debug_3_2 = 1'b1;
      end else begin
        debug_3_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_2 = 1'b0;
    if(when_ArraySlice_l158_20) begin
      if(when_ArraySlice_l159_20) begin
        debug_4_2 = 1'b1;
      end else begin
        debug_4_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_20) begin
        debug_4_2 = 1'b1;
      end else begin
        debug_4_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_2 = 1'b0;
    if(when_ArraySlice_l158_21) begin
      if(when_ArraySlice_l159_21) begin
        debug_5_2 = 1'b1;
      end else begin
        debug_5_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_21) begin
        debug_5_2 = 1'b1;
      end else begin
        debug_5_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_2 = 1'b0;
    if(when_ArraySlice_l158_22) begin
      if(when_ArraySlice_l159_22) begin
        debug_6_2 = 1'b1;
      end else begin
        debug_6_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_22) begin
        debug_6_2 = 1'b1;
      end else begin
        debug_6_2 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_2 = 1'b0;
    if(when_ArraySlice_l158_23) begin
      if(when_ArraySlice_l159_23) begin
        debug_7_2 = 1'b1;
      end else begin
        debug_7_2 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_23) begin
        debug_7_2 = 1'b1;
      end else begin
        debug_7_2 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_16 = (_zz_when_ArraySlice_l158_16 <= _zz_when_ArraySlice_l158_16_3);
  assign when_ArraySlice_l159_16 = (_zz_when_ArraySlice_l159_16 <= _zz_when_ArraySlice_l159_16_1);
  assign _zz_realValue_0_16 = (_zz__zz_realValue_0_16 % _zz__zz_realValue_0_16_1);
  assign when_ArraySlice_l110_16 = (_zz_realValue_0_16 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_16) begin
      realValue_0_16 = (_zz_realValue_0_16_1 - _zz_realValue_0_16);
    end else begin
      realValue_0_16 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_16 = (_zz_when_ArraySlice_l166_16 <= _zz_when_ArraySlice_l166_16_1);
  assign when_ArraySlice_l158_17 = (_zz_when_ArraySlice_l158_17 <= _zz_when_ArraySlice_l158_17_3);
  assign when_ArraySlice_l159_17 = (_zz_when_ArraySlice_l159_17 <= _zz_when_ArraySlice_l159_17_2);
  assign _zz_realValue_0_17 = (_zz__zz_realValue_0_17 % _zz__zz_realValue_0_17_1);
  assign when_ArraySlice_l110_17 = (_zz_realValue_0_17 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_17) begin
      realValue_0_17 = (_zz_realValue_0_17_1 - _zz_realValue_0_17);
    end else begin
      realValue_0_17 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_17 = (_zz_when_ArraySlice_l166_17 <= _zz_when_ArraySlice_l166_17_2);
  assign when_ArraySlice_l158_18 = (_zz_when_ArraySlice_l158_18 <= _zz_when_ArraySlice_l158_18_3);
  assign when_ArraySlice_l159_18 = (_zz_when_ArraySlice_l159_18 <= _zz_when_ArraySlice_l159_18_2);
  assign _zz_realValue_0_18 = (_zz__zz_realValue_0_18 % _zz__zz_realValue_0_18_1);
  assign when_ArraySlice_l110_18 = (_zz_realValue_0_18 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_18) begin
      realValue_0_18 = (_zz_realValue_0_18_1 - _zz_realValue_0_18);
    end else begin
      realValue_0_18 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_18 = (_zz_when_ArraySlice_l166_18 <= _zz_when_ArraySlice_l166_18_2);
  assign when_ArraySlice_l158_19 = (_zz_when_ArraySlice_l158_19 <= _zz_when_ArraySlice_l158_19_3);
  assign when_ArraySlice_l159_19 = (_zz_when_ArraySlice_l159_19 <= _zz_when_ArraySlice_l159_19_2);
  assign _zz_realValue_0_19 = (_zz__zz_realValue_0_19 % _zz__zz_realValue_0_19_1);
  assign when_ArraySlice_l110_19 = (_zz_realValue_0_19 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_19) begin
      realValue_0_19 = (_zz_realValue_0_19_1 - _zz_realValue_0_19);
    end else begin
      realValue_0_19 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_19 = (_zz_when_ArraySlice_l166_19 <= _zz_when_ArraySlice_l166_19_2);
  assign when_ArraySlice_l158_20 = (_zz_when_ArraySlice_l158_20 <= _zz_when_ArraySlice_l158_20_3);
  assign when_ArraySlice_l159_20 = (_zz_when_ArraySlice_l159_20 <= _zz_when_ArraySlice_l159_20_2);
  assign _zz_realValue_0_20 = (_zz__zz_realValue_0_20 % _zz__zz_realValue_0_20_1);
  assign when_ArraySlice_l110_20 = (_zz_realValue_0_20 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_20) begin
      realValue_0_20 = (_zz_realValue_0_20_1 - _zz_realValue_0_20);
    end else begin
      realValue_0_20 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_20 = (_zz_when_ArraySlice_l166_20 <= _zz_when_ArraySlice_l166_20_2);
  assign when_ArraySlice_l158_21 = (_zz_when_ArraySlice_l158_21 <= _zz_when_ArraySlice_l158_21_3);
  assign when_ArraySlice_l159_21 = (_zz_when_ArraySlice_l159_21 <= _zz_when_ArraySlice_l159_21_2);
  assign _zz_realValue_0_21 = (_zz__zz_realValue_0_21 % _zz__zz_realValue_0_21_1);
  assign when_ArraySlice_l110_21 = (_zz_realValue_0_21 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_21) begin
      realValue_0_21 = (_zz_realValue_0_21_1 - _zz_realValue_0_21);
    end else begin
      realValue_0_21 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_21 = (_zz_when_ArraySlice_l166_21 <= _zz_when_ArraySlice_l166_21_2);
  assign when_ArraySlice_l158_22 = (_zz_when_ArraySlice_l158_22 <= _zz_when_ArraySlice_l158_22_3);
  assign when_ArraySlice_l159_22 = (_zz_when_ArraySlice_l159_22 <= _zz_when_ArraySlice_l159_22_2);
  assign _zz_realValue_0_22 = (_zz__zz_realValue_0_22 % _zz__zz_realValue_0_22_1);
  assign when_ArraySlice_l110_22 = (_zz_realValue_0_22 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_22) begin
      realValue_0_22 = (_zz_realValue_0_22_1 - _zz_realValue_0_22);
    end else begin
      realValue_0_22 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_22 = (_zz_when_ArraySlice_l166_22 <= _zz_when_ArraySlice_l166_22_2);
  assign when_ArraySlice_l158_23 = (_zz_when_ArraySlice_l158_23 <= _zz_when_ArraySlice_l158_23_3);
  assign when_ArraySlice_l159_23 = (_zz_when_ArraySlice_l159_23 <= _zz_when_ArraySlice_l159_23_2);
  assign _zz_realValue_0_23 = (_zz__zz_realValue_0_23 % _zz__zz_realValue_0_23_1);
  assign when_ArraySlice_l110_23 = (_zz_realValue_0_23 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_23) begin
      realValue_0_23 = (_zz_realValue_0_23_1 - _zz_realValue_0_23);
    end else begin
      realValue_0_23 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_23 = (_zz_when_ArraySlice_l166_23 <= _zz_when_ArraySlice_l166_23_2);
  assign when_ArraySlice_l425 = (! ((((((_zz_when_ArraySlice_l425 && _zz_when_ArraySlice_l425_1) && (holdReadOp_4 == _zz_when_ArraySlice_l425_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_3 && _zz_when_ArraySlice_l425_4) && (debug_4_2 == _zz_when_ArraySlice_l425_5)) && (debug_5_2 == 1'b1)) && (debug_6_2 == 1'b1)) && (debug_7_2 == 1'b1))));
  assign when_ArraySlice_l428 = (_zz_when_ArraySlice_l428 <= _zz_when_ArraySlice_l428_1);
  assign when_ArraySlice_l431 = (_zz_when_ArraySlice_l431 <= _zz_when_ArraySlice_l431_1);
  assign outputStreamArrayData_0_fire_3 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l438 = ((_zz_when_ArraySlice_l438 == 13'h0) && outputStreamArrayData_0_fire_3);
  assign outputStreamArrayData_0_fire_4 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l449 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l449) && outputStreamArrayData_0_fire_4);
  assign _zz_realValue1_0_2 = (_zz__zz_realValue1_0_2 % _zz__zz_realValue1_0_2_1);
  assign when_ArraySlice_l95_2 = (_zz_realValue1_0_2 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_2) begin
      realValue1_0_2 = (_zz_realValue1_0_2_1 - _zz_realValue1_0_2);
    end else begin
      realValue1_0_2 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450 = (_zz_when_ArraySlice_l450 < _zz_when_ArraySlice_l450_2);
  always @(*) begin
    debug_0_3 = 1'b0;
    if(when_ArraySlice_l158_24) begin
      if(when_ArraySlice_l159_24) begin
        debug_0_3 = 1'b1;
      end else begin
        debug_0_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_24) begin
        debug_0_3 = 1'b1;
      end else begin
        debug_0_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_3 = 1'b0;
    if(when_ArraySlice_l158_25) begin
      if(when_ArraySlice_l159_25) begin
        debug_1_3 = 1'b1;
      end else begin
        debug_1_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_25) begin
        debug_1_3 = 1'b1;
      end else begin
        debug_1_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_3 = 1'b0;
    if(when_ArraySlice_l158_26) begin
      if(when_ArraySlice_l159_26) begin
        debug_2_3 = 1'b1;
      end else begin
        debug_2_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_26) begin
        debug_2_3 = 1'b1;
      end else begin
        debug_2_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_3 = 1'b0;
    if(when_ArraySlice_l158_27) begin
      if(when_ArraySlice_l159_27) begin
        debug_3_3 = 1'b1;
      end else begin
        debug_3_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_27) begin
        debug_3_3 = 1'b1;
      end else begin
        debug_3_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_3 = 1'b0;
    if(when_ArraySlice_l158_28) begin
      if(when_ArraySlice_l159_28) begin
        debug_4_3 = 1'b1;
      end else begin
        debug_4_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_28) begin
        debug_4_3 = 1'b1;
      end else begin
        debug_4_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_3 = 1'b0;
    if(when_ArraySlice_l158_29) begin
      if(when_ArraySlice_l159_29) begin
        debug_5_3 = 1'b1;
      end else begin
        debug_5_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_29) begin
        debug_5_3 = 1'b1;
      end else begin
        debug_5_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_3 = 1'b0;
    if(when_ArraySlice_l158_30) begin
      if(when_ArraySlice_l159_30) begin
        debug_6_3 = 1'b1;
      end else begin
        debug_6_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_30) begin
        debug_6_3 = 1'b1;
      end else begin
        debug_6_3 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_3 = 1'b0;
    if(when_ArraySlice_l158_31) begin
      if(when_ArraySlice_l159_31) begin
        debug_7_3 = 1'b1;
      end else begin
        debug_7_3 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_31) begin
        debug_7_3 = 1'b1;
      end else begin
        debug_7_3 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_24 = (_zz_when_ArraySlice_l158_24 <= _zz_when_ArraySlice_l158_24_3);
  assign when_ArraySlice_l159_24 = (_zz_when_ArraySlice_l159_24 <= _zz_when_ArraySlice_l159_24_1);
  assign _zz_realValue_0_24 = (_zz__zz_realValue_0_24 % _zz__zz_realValue_0_24_1);
  assign when_ArraySlice_l110_24 = (_zz_realValue_0_24 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_24) begin
      realValue_0_24 = (_zz_realValue_0_24_1 - _zz_realValue_0_24);
    end else begin
      realValue_0_24 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_24 = (_zz_when_ArraySlice_l166_24 <= _zz_when_ArraySlice_l166_24_1);
  assign when_ArraySlice_l158_25 = (_zz_when_ArraySlice_l158_25 <= _zz_when_ArraySlice_l158_25_3);
  assign when_ArraySlice_l159_25 = (_zz_when_ArraySlice_l159_25 <= _zz_when_ArraySlice_l159_25_2);
  assign _zz_realValue_0_25 = (_zz__zz_realValue_0_25 % _zz__zz_realValue_0_25_1);
  assign when_ArraySlice_l110_25 = (_zz_realValue_0_25 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_25) begin
      realValue_0_25 = (_zz_realValue_0_25_1 - _zz_realValue_0_25);
    end else begin
      realValue_0_25 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_25 = (_zz_when_ArraySlice_l166_25 <= _zz_when_ArraySlice_l166_25_2);
  assign when_ArraySlice_l158_26 = (_zz_when_ArraySlice_l158_26 <= _zz_when_ArraySlice_l158_26_3);
  assign when_ArraySlice_l159_26 = (_zz_when_ArraySlice_l159_26 <= _zz_when_ArraySlice_l159_26_2);
  assign _zz_realValue_0_26 = (_zz__zz_realValue_0_26 % _zz__zz_realValue_0_26_1);
  assign when_ArraySlice_l110_26 = (_zz_realValue_0_26 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_26) begin
      realValue_0_26 = (_zz_realValue_0_26_1 - _zz_realValue_0_26);
    end else begin
      realValue_0_26 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_26 = (_zz_when_ArraySlice_l166_26 <= _zz_when_ArraySlice_l166_26_2);
  assign when_ArraySlice_l158_27 = (_zz_when_ArraySlice_l158_27 <= _zz_when_ArraySlice_l158_27_3);
  assign when_ArraySlice_l159_27 = (_zz_when_ArraySlice_l159_27 <= _zz_when_ArraySlice_l159_27_2);
  assign _zz_realValue_0_27 = (_zz__zz_realValue_0_27 % _zz__zz_realValue_0_27_1);
  assign when_ArraySlice_l110_27 = (_zz_realValue_0_27 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_27) begin
      realValue_0_27 = (_zz_realValue_0_27_1 - _zz_realValue_0_27);
    end else begin
      realValue_0_27 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_27 = (_zz_when_ArraySlice_l166_27 <= _zz_when_ArraySlice_l166_27_2);
  assign when_ArraySlice_l158_28 = (_zz_when_ArraySlice_l158_28 <= _zz_when_ArraySlice_l158_28_3);
  assign when_ArraySlice_l159_28 = (_zz_when_ArraySlice_l159_28 <= _zz_when_ArraySlice_l159_28_2);
  assign _zz_realValue_0_28 = (_zz__zz_realValue_0_28 % _zz__zz_realValue_0_28_1);
  assign when_ArraySlice_l110_28 = (_zz_realValue_0_28 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_28) begin
      realValue_0_28 = (_zz_realValue_0_28_1 - _zz_realValue_0_28);
    end else begin
      realValue_0_28 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_28 = (_zz_when_ArraySlice_l166_28 <= _zz_when_ArraySlice_l166_28_2);
  assign when_ArraySlice_l158_29 = (_zz_when_ArraySlice_l158_29 <= _zz_when_ArraySlice_l158_29_3);
  assign when_ArraySlice_l159_29 = (_zz_when_ArraySlice_l159_29 <= _zz_when_ArraySlice_l159_29_2);
  assign _zz_realValue_0_29 = (_zz__zz_realValue_0_29 % _zz__zz_realValue_0_29_1);
  assign when_ArraySlice_l110_29 = (_zz_realValue_0_29 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_29) begin
      realValue_0_29 = (_zz_realValue_0_29_1 - _zz_realValue_0_29);
    end else begin
      realValue_0_29 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_29 = (_zz_when_ArraySlice_l166_29 <= _zz_when_ArraySlice_l166_29_2);
  assign when_ArraySlice_l158_30 = (_zz_when_ArraySlice_l158_30 <= _zz_when_ArraySlice_l158_30_3);
  assign when_ArraySlice_l159_30 = (_zz_when_ArraySlice_l159_30 <= _zz_when_ArraySlice_l159_30_2);
  assign _zz_realValue_0_30 = (_zz__zz_realValue_0_30 % _zz__zz_realValue_0_30_1);
  assign when_ArraySlice_l110_30 = (_zz_realValue_0_30 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_30) begin
      realValue_0_30 = (_zz_realValue_0_30_1 - _zz_realValue_0_30);
    end else begin
      realValue_0_30 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_30 = (_zz_when_ArraySlice_l166_30 <= _zz_when_ArraySlice_l166_30_2);
  assign when_ArraySlice_l158_31 = (_zz_when_ArraySlice_l158_31 <= _zz_when_ArraySlice_l158_31_3);
  assign when_ArraySlice_l159_31 = (_zz_when_ArraySlice_l159_31 <= _zz_when_ArraySlice_l159_31_2);
  assign _zz_realValue_0_31 = (_zz__zz_realValue_0_31 % _zz__zz_realValue_0_31_1);
  assign when_ArraySlice_l110_31 = (_zz_realValue_0_31 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_31) begin
      realValue_0_31 = (_zz_realValue_0_31_1 - _zz_realValue_0_31);
    end else begin
      realValue_0_31 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_31 = (_zz_when_ArraySlice_l166_31 <= _zz_when_ArraySlice_l166_31_2);
  assign when_ArraySlice_l457 = (! ((((((_zz_when_ArraySlice_l457 && _zz_when_ArraySlice_l457_1) && (holdReadOp_4 == _zz_when_ArraySlice_l457_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_3 && _zz_when_ArraySlice_l457_4) && (debug_4_3 == _zz_when_ArraySlice_l457_5)) && (debug_5_3 == 1'b1)) && (debug_6_3 == 1'b1)) && (debug_7_3 == 1'b1))));
  assign outputStreamArrayData_0_fire_5 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l461 = ((_zz_when_ArraySlice_l461 == 13'h0) && outputStreamArrayData_0_fire_5);
  assign when_ArraySlice_l447 = (allowPadding_0 && (_zz_when_ArraySlice_l447 <= _zz_when_ArraySlice_l447_1));
  assign outputStreamArrayData_0_fire_6 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l468 = (handshakeTimes_0_value == _zz_when_ArraySlice_l468);
  assign when_ArraySlice_l376_1 = (_zz_when_ArraySlice_l376_1_1 < _zz_when_ArraySlice_l376_1_4);
  assign when_ArraySlice_l377_1 = ((! holdReadOp_1) && (_zz_when_ArraySlice_l377_1_1 != 7'h0));
  assign _zz_outputStreamArrayData_1_valid = (selectReadFifo_1 + _zz__zz_outputStreamArrayData_1_valid);
  assign _zz_4 = ({127'd0,1'b1} <<< _zz__zz_4);
  assign _zz_io_pop_ready_1 = outputStreamArrayData_1_ready;
  assign when_ArraySlice_l382_1 = (! holdReadOp_1);
  assign outputStreamArrayData_1_fire = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l383_1 = ((7'h01 < _zz_when_ArraySlice_l383_1_1) && outputStreamArrayData_1_fire);
  assign when_ArraySlice_l384_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l384_1_1);
  assign when_ArraySlice_l387_1 = (_zz_when_ArraySlice_l387_1_1 == 13'h0);
  assign outputStreamArrayData_1_fire_1 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l392_1 = ((_zz_when_ArraySlice_l392_1_1 == 7'h01) && outputStreamArrayData_1_fire_1);
  assign when_ArraySlice_l393_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l393_1_1);
  assign _zz_realValue1_0_3 = (_zz__zz_realValue1_0_3 % _zz__zz_realValue1_0_3_1);
  assign when_ArraySlice_l95_3 = (_zz_realValue1_0_3 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_3) begin
      realValue1_0_3 = (_zz_realValue1_0_3_1 - _zz_realValue1_0_3);
    end else begin
      realValue1_0_3 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_1 = (_zz_when_ArraySlice_l395_1_1 < _zz_when_ArraySlice_l395_1_3);
  always @(*) begin
    debug_0_4 = 1'b0;
    if(when_ArraySlice_l158_32) begin
      if(when_ArraySlice_l159_32) begin
        debug_0_4 = 1'b1;
      end else begin
        debug_0_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_32) begin
        debug_0_4 = 1'b1;
      end else begin
        debug_0_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_4 = 1'b0;
    if(when_ArraySlice_l158_33) begin
      if(when_ArraySlice_l159_33) begin
        debug_1_4 = 1'b1;
      end else begin
        debug_1_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_33) begin
        debug_1_4 = 1'b1;
      end else begin
        debug_1_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_4 = 1'b0;
    if(when_ArraySlice_l158_34) begin
      if(when_ArraySlice_l159_34) begin
        debug_2_4 = 1'b1;
      end else begin
        debug_2_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_34) begin
        debug_2_4 = 1'b1;
      end else begin
        debug_2_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_4 = 1'b0;
    if(when_ArraySlice_l158_35) begin
      if(when_ArraySlice_l159_35) begin
        debug_3_4 = 1'b1;
      end else begin
        debug_3_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_35) begin
        debug_3_4 = 1'b1;
      end else begin
        debug_3_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_4 = 1'b0;
    if(when_ArraySlice_l158_36) begin
      if(when_ArraySlice_l159_36) begin
        debug_4_4 = 1'b1;
      end else begin
        debug_4_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_36) begin
        debug_4_4 = 1'b1;
      end else begin
        debug_4_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_4 = 1'b0;
    if(when_ArraySlice_l158_37) begin
      if(when_ArraySlice_l159_37) begin
        debug_5_4 = 1'b1;
      end else begin
        debug_5_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_37) begin
        debug_5_4 = 1'b1;
      end else begin
        debug_5_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_4 = 1'b0;
    if(when_ArraySlice_l158_38) begin
      if(when_ArraySlice_l159_38) begin
        debug_6_4 = 1'b1;
      end else begin
        debug_6_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_38) begin
        debug_6_4 = 1'b1;
      end else begin
        debug_6_4 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_4 = 1'b0;
    if(when_ArraySlice_l158_39) begin
      if(when_ArraySlice_l159_39) begin
        debug_7_4 = 1'b1;
      end else begin
        debug_7_4 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_39) begin
        debug_7_4 = 1'b1;
      end else begin
        debug_7_4 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_32 = (_zz_when_ArraySlice_l158_32 <= _zz_when_ArraySlice_l158_32_3);
  assign when_ArraySlice_l159_32 = (_zz_when_ArraySlice_l159_32 <= _zz_when_ArraySlice_l159_32_1);
  assign _zz_realValue_0_32 = (_zz__zz_realValue_0_32 % _zz__zz_realValue_0_32_1);
  assign when_ArraySlice_l110_32 = (_zz_realValue_0_32 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_32) begin
      realValue_0_32 = (_zz_realValue_0_32_1 - _zz_realValue_0_32);
    end else begin
      realValue_0_32 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_32 = (_zz_when_ArraySlice_l166_32 <= _zz_when_ArraySlice_l166_32_1);
  assign when_ArraySlice_l158_33 = (_zz_when_ArraySlice_l158_33 <= _zz_when_ArraySlice_l158_33_3);
  assign when_ArraySlice_l159_33 = (_zz_when_ArraySlice_l159_33 <= _zz_when_ArraySlice_l159_33_2);
  assign _zz_realValue_0_33 = (_zz__zz_realValue_0_33 % _zz__zz_realValue_0_33_1);
  assign when_ArraySlice_l110_33 = (_zz_realValue_0_33 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_33) begin
      realValue_0_33 = (_zz_realValue_0_33_1 - _zz_realValue_0_33);
    end else begin
      realValue_0_33 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_33 = (_zz_when_ArraySlice_l166_33 <= _zz_when_ArraySlice_l166_33_2);
  assign when_ArraySlice_l158_34 = (_zz_when_ArraySlice_l158_34 <= _zz_when_ArraySlice_l158_34_3);
  assign when_ArraySlice_l159_34 = (_zz_when_ArraySlice_l159_34 <= _zz_when_ArraySlice_l159_34_2);
  assign _zz_realValue_0_34 = (_zz__zz_realValue_0_34 % _zz__zz_realValue_0_34_1);
  assign when_ArraySlice_l110_34 = (_zz_realValue_0_34 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_34) begin
      realValue_0_34 = (_zz_realValue_0_34_1 - _zz_realValue_0_34);
    end else begin
      realValue_0_34 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_34 = (_zz_when_ArraySlice_l166_34 <= _zz_when_ArraySlice_l166_34_2);
  assign when_ArraySlice_l158_35 = (_zz_when_ArraySlice_l158_35 <= _zz_when_ArraySlice_l158_35_3);
  assign when_ArraySlice_l159_35 = (_zz_when_ArraySlice_l159_35 <= _zz_when_ArraySlice_l159_35_2);
  assign _zz_realValue_0_35 = (_zz__zz_realValue_0_35 % _zz__zz_realValue_0_35_1);
  assign when_ArraySlice_l110_35 = (_zz_realValue_0_35 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_35) begin
      realValue_0_35 = (_zz_realValue_0_35_1 - _zz_realValue_0_35);
    end else begin
      realValue_0_35 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_35 = (_zz_when_ArraySlice_l166_35 <= _zz_when_ArraySlice_l166_35_2);
  assign when_ArraySlice_l158_36 = (_zz_when_ArraySlice_l158_36 <= _zz_when_ArraySlice_l158_36_3);
  assign when_ArraySlice_l159_36 = (_zz_when_ArraySlice_l159_36 <= _zz_when_ArraySlice_l159_36_2);
  assign _zz_realValue_0_36 = (_zz__zz_realValue_0_36 % _zz__zz_realValue_0_36_1);
  assign when_ArraySlice_l110_36 = (_zz_realValue_0_36 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_36) begin
      realValue_0_36 = (_zz_realValue_0_36_1 - _zz_realValue_0_36);
    end else begin
      realValue_0_36 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_36 = (_zz_when_ArraySlice_l166_36 <= _zz_when_ArraySlice_l166_36_2);
  assign when_ArraySlice_l158_37 = (_zz_when_ArraySlice_l158_37 <= _zz_when_ArraySlice_l158_37_3);
  assign when_ArraySlice_l159_37 = (_zz_when_ArraySlice_l159_37 <= _zz_when_ArraySlice_l159_37_2);
  assign _zz_realValue_0_37 = (_zz__zz_realValue_0_37 % _zz__zz_realValue_0_37_1);
  assign when_ArraySlice_l110_37 = (_zz_realValue_0_37 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_37) begin
      realValue_0_37 = (_zz_realValue_0_37_1 - _zz_realValue_0_37);
    end else begin
      realValue_0_37 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_37 = (_zz_when_ArraySlice_l166_37 <= _zz_when_ArraySlice_l166_37_2);
  assign when_ArraySlice_l158_38 = (_zz_when_ArraySlice_l158_38 <= _zz_when_ArraySlice_l158_38_3);
  assign when_ArraySlice_l159_38 = (_zz_when_ArraySlice_l159_38 <= _zz_when_ArraySlice_l159_38_2);
  assign _zz_realValue_0_38 = (_zz__zz_realValue_0_38 % _zz__zz_realValue_0_38_1);
  assign when_ArraySlice_l110_38 = (_zz_realValue_0_38 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_38) begin
      realValue_0_38 = (_zz_realValue_0_38_1 - _zz_realValue_0_38);
    end else begin
      realValue_0_38 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_38 = (_zz_when_ArraySlice_l166_38 <= _zz_when_ArraySlice_l166_38_2);
  assign when_ArraySlice_l158_39 = (_zz_when_ArraySlice_l158_39 <= _zz_when_ArraySlice_l158_39_3);
  assign when_ArraySlice_l159_39 = (_zz_when_ArraySlice_l159_39 <= _zz_when_ArraySlice_l159_39_2);
  assign _zz_realValue_0_39 = (_zz__zz_realValue_0_39 % _zz__zz_realValue_0_39_1);
  assign when_ArraySlice_l110_39 = (_zz_realValue_0_39 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_39) begin
      realValue_0_39 = (_zz_realValue_0_39_1 - _zz_realValue_0_39);
    end else begin
      realValue_0_39 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_39 = (_zz_when_ArraySlice_l166_39 <= _zz_when_ArraySlice_l166_39_2);
  assign when_ArraySlice_l400_1 = (! ((((((_zz_when_ArraySlice_l400_1_1 && _zz_when_ArraySlice_l400_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_1_4 && _zz_when_ArraySlice_l400_1_5) && (debug_4_4 == _zz_when_ArraySlice_l400_1_6)) && (debug_5_4 == 1'b1)) && (debug_6_4 == 1'b1)) && (debug_7_4 == 1'b1))));
  assign when_ArraySlice_l403_1 = (_zz_when_ArraySlice_l403_1_1 <= _zz_when_ArraySlice_l403_1_2);
  assign when_ArraySlice_l406_1 = (_zz_when_ArraySlice_l406_1_1 <= _zz_when_ArraySlice_l406_1_2);
  assign when_ArraySlice_l413_1 = (_zz_when_ArraySlice_l413_1_1 == 13'h0);
  assign when_ArraySlice_l417_1 = (_zz_when_ArraySlice_l417_1_1 == 7'h0);
  assign outputStreamArrayData_1_fire_2 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l418_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l418_1_1) && outputStreamArrayData_1_fire_2);
  assign _zz_realValue1_0_4 = (_zz__zz_realValue1_0_4 % _zz__zz_realValue1_0_4_1);
  assign when_ArraySlice_l95_4 = (_zz_realValue1_0_4 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_4) begin
      realValue1_0_4 = (_zz_realValue1_0_4_1 - _zz_realValue1_0_4);
    end else begin
      realValue1_0_4 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_1 = (_zz_when_ArraySlice_l420_1_1 < _zz_when_ArraySlice_l420_1_3);
  always @(*) begin
    debug_0_5 = 1'b0;
    if(when_ArraySlice_l158_40) begin
      if(when_ArraySlice_l159_40) begin
        debug_0_5 = 1'b1;
      end else begin
        debug_0_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_40) begin
        debug_0_5 = 1'b1;
      end else begin
        debug_0_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_5 = 1'b0;
    if(when_ArraySlice_l158_41) begin
      if(when_ArraySlice_l159_41) begin
        debug_1_5 = 1'b1;
      end else begin
        debug_1_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_41) begin
        debug_1_5 = 1'b1;
      end else begin
        debug_1_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_5 = 1'b0;
    if(when_ArraySlice_l158_42) begin
      if(when_ArraySlice_l159_42) begin
        debug_2_5 = 1'b1;
      end else begin
        debug_2_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_42) begin
        debug_2_5 = 1'b1;
      end else begin
        debug_2_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_5 = 1'b0;
    if(when_ArraySlice_l158_43) begin
      if(when_ArraySlice_l159_43) begin
        debug_3_5 = 1'b1;
      end else begin
        debug_3_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_43) begin
        debug_3_5 = 1'b1;
      end else begin
        debug_3_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_5 = 1'b0;
    if(when_ArraySlice_l158_44) begin
      if(when_ArraySlice_l159_44) begin
        debug_4_5 = 1'b1;
      end else begin
        debug_4_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_44) begin
        debug_4_5 = 1'b1;
      end else begin
        debug_4_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_5 = 1'b0;
    if(when_ArraySlice_l158_45) begin
      if(when_ArraySlice_l159_45) begin
        debug_5_5 = 1'b1;
      end else begin
        debug_5_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_45) begin
        debug_5_5 = 1'b1;
      end else begin
        debug_5_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_5 = 1'b0;
    if(when_ArraySlice_l158_46) begin
      if(when_ArraySlice_l159_46) begin
        debug_6_5 = 1'b1;
      end else begin
        debug_6_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_46) begin
        debug_6_5 = 1'b1;
      end else begin
        debug_6_5 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_5 = 1'b0;
    if(when_ArraySlice_l158_47) begin
      if(when_ArraySlice_l159_47) begin
        debug_7_5 = 1'b1;
      end else begin
        debug_7_5 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_47) begin
        debug_7_5 = 1'b1;
      end else begin
        debug_7_5 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_40 = (_zz_when_ArraySlice_l158_40 <= _zz_when_ArraySlice_l158_40_3);
  assign when_ArraySlice_l159_40 = (_zz_when_ArraySlice_l159_40 <= _zz_when_ArraySlice_l159_40_1);
  assign _zz_realValue_0_40 = (_zz__zz_realValue_0_40 % _zz__zz_realValue_0_40_1);
  assign when_ArraySlice_l110_40 = (_zz_realValue_0_40 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_40) begin
      realValue_0_40 = (_zz_realValue_0_40_1 - _zz_realValue_0_40);
    end else begin
      realValue_0_40 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_40 = (_zz_when_ArraySlice_l166_40 <= _zz_when_ArraySlice_l166_40_1);
  assign when_ArraySlice_l158_41 = (_zz_when_ArraySlice_l158_41 <= _zz_when_ArraySlice_l158_41_3);
  assign when_ArraySlice_l159_41 = (_zz_when_ArraySlice_l159_41 <= _zz_when_ArraySlice_l159_41_2);
  assign _zz_realValue_0_41 = (_zz__zz_realValue_0_41 % _zz__zz_realValue_0_41_1);
  assign when_ArraySlice_l110_41 = (_zz_realValue_0_41 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_41) begin
      realValue_0_41 = (_zz_realValue_0_41_1 - _zz_realValue_0_41);
    end else begin
      realValue_0_41 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_41 = (_zz_when_ArraySlice_l166_41 <= _zz_when_ArraySlice_l166_41_2);
  assign when_ArraySlice_l158_42 = (_zz_when_ArraySlice_l158_42 <= _zz_when_ArraySlice_l158_42_3);
  assign when_ArraySlice_l159_42 = (_zz_when_ArraySlice_l159_42 <= _zz_when_ArraySlice_l159_42_2);
  assign _zz_realValue_0_42 = (_zz__zz_realValue_0_42 % _zz__zz_realValue_0_42_1);
  assign when_ArraySlice_l110_42 = (_zz_realValue_0_42 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_42) begin
      realValue_0_42 = (_zz_realValue_0_42_1 - _zz_realValue_0_42);
    end else begin
      realValue_0_42 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_42 = (_zz_when_ArraySlice_l166_42 <= _zz_when_ArraySlice_l166_42_2);
  assign when_ArraySlice_l158_43 = (_zz_when_ArraySlice_l158_43 <= _zz_when_ArraySlice_l158_43_3);
  assign when_ArraySlice_l159_43 = (_zz_when_ArraySlice_l159_43 <= _zz_when_ArraySlice_l159_43_2);
  assign _zz_realValue_0_43 = (_zz__zz_realValue_0_43 % _zz__zz_realValue_0_43_1);
  assign when_ArraySlice_l110_43 = (_zz_realValue_0_43 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_43) begin
      realValue_0_43 = (_zz_realValue_0_43_1 - _zz_realValue_0_43);
    end else begin
      realValue_0_43 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_43 = (_zz_when_ArraySlice_l166_43 <= _zz_when_ArraySlice_l166_43_2);
  assign when_ArraySlice_l158_44 = (_zz_when_ArraySlice_l158_44 <= _zz_when_ArraySlice_l158_44_3);
  assign when_ArraySlice_l159_44 = (_zz_when_ArraySlice_l159_44 <= _zz_when_ArraySlice_l159_44_2);
  assign _zz_realValue_0_44 = (_zz__zz_realValue_0_44 % _zz__zz_realValue_0_44_1);
  assign when_ArraySlice_l110_44 = (_zz_realValue_0_44 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_44) begin
      realValue_0_44 = (_zz_realValue_0_44_1 - _zz_realValue_0_44);
    end else begin
      realValue_0_44 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_44 = (_zz_when_ArraySlice_l166_44 <= _zz_when_ArraySlice_l166_44_2);
  assign when_ArraySlice_l158_45 = (_zz_when_ArraySlice_l158_45 <= _zz_when_ArraySlice_l158_45_3);
  assign when_ArraySlice_l159_45 = (_zz_when_ArraySlice_l159_45 <= _zz_when_ArraySlice_l159_45_2);
  assign _zz_realValue_0_45 = (_zz__zz_realValue_0_45 % _zz__zz_realValue_0_45_1);
  assign when_ArraySlice_l110_45 = (_zz_realValue_0_45 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_45) begin
      realValue_0_45 = (_zz_realValue_0_45_1 - _zz_realValue_0_45);
    end else begin
      realValue_0_45 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_45 = (_zz_when_ArraySlice_l166_45 <= _zz_when_ArraySlice_l166_45_2);
  assign when_ArraySlice_l158_46 = (_zz_when_ArraySlice_l158_46 <= _zz_when_ArraySlice_l158_46_3);
  assign when_ArraySlice_l159_46 = (_zz_when_ArraySlice_l159_46 <= _zz_when_ArraySlice_l159_46_2);
  assign _zz_realValue_0_46 = (_zz__zz_realValue_0_46 % _zz__zz_realValue_0_46_1);
  assign when_ArraySlice_l110_46 = (_zz_realValue_0_46 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_46) begin
      realValue_0_46 = (_zz_realValue_0_46_1 - _zz_realValue_0_46);
    end else begin
      realValue_0_46 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_46 = (_zz_when_ArraySlice_l166_46 <= _zz_when_ArraySlice_l166_46_2);
  assign when_ArraySlice_l158_47 = (_zz_when_ArraySlice_l158_47 <= _zz_when_ArraySlice_l158_47_3);
  assign when_ArraySlice_l159_47 = (_zz_when_ArraySlice_l159_47 <= _zz_when_ArraySlice_l159_47_2);
  assign _zz_realValue_0_47 = (_zz__zz_realValue_0_47 % _zz__zz_realValue_0_47_1);
  assign when_ArraySlice_l110_47 = (_zz_realValue_0_47 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_47) begin
      realValue_0_47 = (_zz_realValue_0_47_1 - _zz_realValue_0_47);
    end else begin
      realValue_0_47 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_47 = (_zz_when_ArraySlice_l166_47 <= _zz_when_ArraySlice_l166_47_2);
  assign when_ArraySlice_l425_1 = (! ((((((_zz_when_ArraySlice_l425_1_1 && _zz_when_ArraySlice_l425_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l425_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_1_4 && _zz_when_ArraySlice_l425_1_5) && (debug_4_5 == _zz_when_ArraySlice_l425_1_6)) && (debug_5_5 == 1'b1)) && (debug_6_5 == 1'b1)) && (debug_7_5 == 1'b1))));
  assign when_ArraySlice_l428_1 = (_zz_when_ArraySlice_l428_1_1 <= _zz_when_ArraySlice_l428_1_2);
  assign when_ArraySlice_l431_1 = (_zz_when_ArraySlice_l431_1_1 <= _zz_when_ArraySlice_l431_1_2);
  assign outputStreamArrayData_1_fire_3 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l438_1 = ((_zz_when_ArraySlice_l438_1_1 == 13'h0) && outputStreamArrayData_1_fire_3);
  assign outputStreamArrayData_1_fire_4 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l449_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l449_1_1) && outputStreamArrayData_1_fire_4);
  assign _zz_realValue1_0_5 = (_zz__zz_realValue1_0_5 % _zz__zz_realValue1_0_5_1);
  assign when_ArraySlice_l95_5 = (_zz_realValue1_0_5 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_5) begin
      realValue1_0_5 = (_zz_realValue1_0_5_1 - _zz_realValue1_0_5);
    end else begin
      realValue1_0_5 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_1 = (_zz_when_ArraySlice_l450_1_1 < _zz_when_ArraySlice_l450_1_3);
  always @(*) begin
    debug_0_6 = 1'b0;
    if(when_ArraySlice_l158_48) begin
      if(when_ArraySlice_l159_48) begin
        debug_0_6 = 1'b1;
      end else begin
        debug_0_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_48) begin
        debug_0_6 = 1'b1;
      end else begin
        debug_0_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_6 = 1'b0;
    if(when_ArraySlice_l158_49) begin
      if(when_ArraySlice_l159_49) begin
        debug_1_6 = 1'b1;
      end else begin
        debug_1_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_49) begin
        debug_1_6 = 1'b1;
      end else begin
        debug_1_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_6 = 1'b0;
    if(when_ArraySlice_l158_50) begin
      if(when_ArraySlice_l159_50) begin
        debug_2_6 = 1'b1;
      end else begin
        debug_2_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_50) begin
        debug_2_6 = 1'b1;
      end else begin
        debug_2_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_6 = 1'b0;
    if(when_ArraySlice_l158_51) begin
      if(when_ArraySlice_l159_51) begin
        debug_3_6 = 1'b1;
      end else begin
        debug_3_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_51) begin
        debug_3_6 = 1'b1;
      end else begin
        debug_3_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_6 = 1'b0;
    if(when_ArraySlice_l158_52) begin
      if(when_ArraySlice_l159_52) begin
        debug_4_6 = 1'b1;
      end else begin
        debug_4_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_52) begin
        debug_4_6 = 1'b1;
      end else begin
        debug_4_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_6 = 1'b0;
    if(when_ArraySlice_l158_53) begin
      if(when_ArraySlice_l159_53) begin
        debug_5_6 = 1'b1;
      end else begin
        debug_5_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_53) begin
        debug_5_6 = 1'b1;
      end else begin
        debug_5_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_6 = 1'b0;
    if(when_ArraySlice_l158_54) begin
      if(when_ArraySlice_l159_54) begin
        debug_6_6 = 1'b1;
      end else begin
        debug_6_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_54) begin
        debug_6_6 = 1'b1;
      end else begin
        debug_6_6 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_6 = 1'b0;
    if(when_ArraySlice_l158_55) begin
      if(when_ArraySlice_l159_55) begin
        debug_7_6 = 1'b1;
      end else begin
        debug_7_6 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_55) begin
        debug_7_6 = 1'b1;
      end else begin
        debug_7_6 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_48 = (_zz_when_ArraySlice_l158_48 <= _zz_when_ArraySlice_l158_48_3);
  assign when_ArraySlice_l159_48 = (_zz_when_ArraySlice_l159_48 <= _zz_when_ArraySlice_l159_48_1);
  assign _zz_realValue_0_48 = (_zz__zz_realValue_0_48 % _zz__zz_realValue_0_48_1);
  assign when_ArraySlice_l110_48 = (_zz_realValue_0_48 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_48) begin
      realValue_0_48 = (_zz_realValue_0_48_1 - _zz_realValue_0_48);
    end else begin
      realValue_0_48 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_48 = (_zz_when_ArraySlice_l166_48 <= _zz_when_ArraySlice_l166_48_1);
  assign when_ArraySlice_l158_49 = (_zz_when_ArraySlice_l158_49 <= _zz_when_ArraySlice_l158_49_3);
  assign when_ArraySlice_l159_49 = (_zz_when_ArraySlice_l159_49 <= _zz_when_ArraySlice_l159_49_2);
  assign _zz_realValue_0_49 = (_zz__zz_realValue_0_49 % _zz__zz_realValue_0_49_1);
  assign when_ArraySlice_l110_49 = (_zz_realValue_0_49 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_49) begin
      realValue_0_49 = (_zz_realValue_0_49_1 - _zz_realValue_0_49);
    end else begin
      realValue_0_49 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_49 = (_zz_when_ArraySlice_l166_49 <= _zz_when_ArraySlice_l166_49_2);
  assign when_ArraySlice_l158_50 = (_zz_when_ArraySlice_l158_50 <= _zz_when_ArraySlice_l158_50_3);
  assign when_ArraySlice_l159_50 = (_zz_when_ArraySlice_l159_50 <= _zz_when_ArraySlice_l159_50_2);
  assign _zz_realValue_0_50 = (_zz__zz_realValue_0_50 % _zz__zz_realValue_0_50_1);
  assign when_ArraySlice_l110_50 = (_zz_realValue_0_50 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_50) begin
      realValue_0_50 = (_zz_realValue_0_50_1 - _zz_realValue_0_50);
    end else begin
      realValue_0_50 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_50 = (_zz_when_ArraySlice_l166_50 <= _zz_when_ArraySlice_l166_50_2);
  assign when_ArraySlice_l158_51 = (_zz_when_ArraySlice_l158_51 <= _zz_when_ArraySlice_l158_51_3);
  assign when_ArraySlice_l159_51 = (_zz_when_ArraySlice_l159_51 <= _zz_when_ArraySlice_l159_51_2);
  assign _zz_realValue_0_51 = (_zz__zz_realValue_0_51 % _zz__zz_realValue_0_51_1);
  assign when_ArraySlice_l110_51 = (_zz_realValue_0_51 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_51) begin
      realValue_0_51 = (_zz_realValue_0_51_1 - _zz_realValue_0_51);
    end else begin
      realValue_0_51 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_51 = (_zz_when_ArraySlice_l166_51 <= _zz_when_ArraySlice_l166_51_2);
  assign when_ArraySlice_l158_52 = (_zz_when_ArraySlice_l158_52 <= _zz_when_ArraySlice_l158_52_3);
  assign when_ArraySlice_l159_52 = (_zz_when_ArraySlice_l159_52 <= _zz_when_ArraySlice_l159_52_2);
  assign _zz_realValue_0_52 = (_zz__zz_realValue_0_52 % _zz__zz_realValue_0_52_1);
  assign when_ArraySlice_l110_52 = (_zz_realValue_0_52 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_52) begin
      realValue_0_52 = (_zz_realValue_0_52_1 - _zz_realValue_0_52);
    end else begin
      realValue_0_52 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_52 = (_zz_when_ArraySlice_l166_52 <= _zz_when_ArraySlice_l166_52_2);
  assign when_ArraySlice_l158_53 = (_zz_when_ArraySlice_l158_53 <= _zz_when_ArraySlice_l158_53_3);
  assign when_ArraySlice_l159_53 = (_zz_when_ArraySlice_l159_53 <= _zz_when_ArraySlice_l159_53_2);
  assign _zz_realValue_0_53 = (_zz__zz_realValue_0_53 % _zz__zz_realValue_0_53_1);
  assign when_ArraySlice_l110_53 = (_zz_realValue_0_53 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_53) begin
      realValue_0_53 = (_zz_realValue_0_53_1 - _zz_realValue_0_53);
    end else begin
      realValue_0_53 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_53 = (_zz_when_ArraySlice_l166_53 <= _zz_when_ArraySlice_l166_53_2);
  assign when_ArraySlice_l158_54 = (_zz_when_ArraySlice_l158_54 <= _zz_when_ArraySlice_l158_54_3);
  assign when_ArraySlice_l159_54 = (_zz_when_ArraySlice_l159_54 <= _zz_when_ArraySlice_l159_54_2);
  assign _zz_realValue_0_54 = (_zz__zz_realValue_0_54 % _zz__zz_realValue_0_54_1);
  assign when_ArraySlice_l110_54 = (_zz_realValue_0_54 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_54) begin
      realValue_0_54 = (_zz_realValue_0_54_1 - _zz_realValue_0_54);
    end else begin
      realValue_0_54 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_54 = (_zz_when_ArraySlice_l166_54 <= _zz_when_ArraySlice_l166_54_2);
  assign when_ArraySlice_l158_55 = (_zz_when_ArraySlice_l158_55 <= _zz_when_ArraySlice_l158_55_3);
  assign when_ArraySlice_l159_55 = (_zz_when_ArraySlice_l159_55 <= _zz_when_ArraySlice_l159_55_2);
  assign _zz_realValue_0_55 = (_zz__zz_realValue_0_55 % _zz__zz_realValue_0_55_1);
  assign when_ArraySlice_l110_55 = (_zz_realValue_0_55 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_55) begin
      realValue_0_55 = (_zz_realValue_0_55_1 - _zz_realValue_0_55);
    end else begin
      realValue_0_55 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_55 = (_zz_when_ArraySlice_l166_55 <= _zz_when_ArraySlice_l166_55_2);
  assign when_ArraySlice_l457_1 = (! ((((((_zz_when_ArraySlice_l457_1_1 && _zz_when_ArraySlice_l457_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l457_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_1_4 && _zz_when_ArraySlice_l457_1_5) && (debug_4_6 == _zz_when_ArraySlice_l457_1_6)) && (debug_5_6 == 1'b1)) && (debug_6_6 == 1'b1)) && (debug_7_6 == 1'b1))));
  assign outputStreamArrayData_1_fire_5 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l461_1 = ((_zz_when_ArraySlice_l461_1_1 == 13'h0) && outputStreamArrayData_1_fire_5);
  assign when_ArraySlice_l447_1 = (allowPadding_1 && (_zz_when_ArraySlice_l447_1_1 <= _zz_when_ArraySlice_l447_1_2));
  assign outputStreamArrayData_1_fire_6 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l468_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l468_1_1);
  assign when_ArraySlice_l376_2 = (_zz_when_ArraySlice_l376_2_1 < _zz_when_ArraySlice_l376_2_4);
  assign when_ArraySlice_l377_2 = ((! holdReadOp_2) && (_zz_when_ArraySlice_l377_2_1 != 7'h0));
  assign _zz_outputStreamArrayData_2_valid = (selectReadFifo_2 + _zz__zz_outputStreamArrayData_2_valid);
  assign _zz_5 = ({127'd0,1'b1} <<< _zz__zz_5);
  assign _zz_io_pop_ready_2 = outputStreamArrayData_2_ready;
  assign when_ArraySlice_l382_2 = (! holdReadOp_2);
  assign outputStreamArrayData_2_fire = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l383_2 = ((7'h01 < _zz_when_ArraySlice_l383_2_1) && outputStreamArrayData_2_fire);
  assign when_ArraySlice_l384_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l384_2_1);
  assign when_ArraySlice_l387_2 = (_zz_when_ArraySlice_l387_2 == 13'h0);
  assign outputStreamArrayData_2_fire_1 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l392_2 = ((_zz_when_ArraySlice_l392_2_1 == 7'h01) && outputStreamArrayData_2_fire_1);
  assign when_ArraySlice_l393_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l393_2_1);
  assign _zz_realValue1_0_6 = (_zz__zz_realValue1_0_6 % _zz__zz_realValue1_0_6_1);
  assign when_ArraySlice_l95_6 = (_zz_realValue1_0_6 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_6) begin
      realValue1_0_6 = (_zz_realValue1_0_6_1 - _zz_realValue1_0_6);
    end else begin
      realValue1_0_6 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_2 = (_zz_when_ArraySlice_l395_2_1 < _zz_when_ArraySlice_l395_2_3);
  always @(*) begin
    debug_0_7 = 1'b0;
    if(when_ArraySlice_l158_56) begin
      if(when_ArraySlice_l159_56) begin
        debug_0_7 = 1'b1;
      end else begin
        debug_0_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_56) begin
        debug_0_7 = 1'b1;
      end else begin
        debug_0_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_7 = 1'b0;
    if(when_ArraySlice_l158_57) begin
      if(when_ArraySlice_l159_57) begin
        debug_1_7 = 1'b1;
      end else begin
        debug_1_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_57) begin
        debug_1_7 = 1'b1;
      end else begin
        debug_1_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_7 = 1'b0;
    if(when_ArraySlice_l158_58) begin
      if(when_ArraySlice_l159_58) begin
        debug_2_7 = 1'b1;
      end else begin
        debug_2_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_58) begin
        debug_2_7 = 1'b1;
      end else begin
        debug_2_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_7 = 1'b0;
    if(when_ArraySlice_l158_59) begin
      if(when_ArraySlice_l159_59) begin
        debug_3_7 = 1'b1;
      end else begin
        debug_3_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_59) begin
        debug_3_7 = 1'b1;
      end else begin
        debug_3_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_7 = 1'b0;
    if(when_ArraySlice_l158_60) begin
      if(when_ArraySlice_l159_60) begin
        debug_4_7 = 1'b1;
      end else begin
        debug_4_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_60) begin
        debug_4_7 = 1'b1;
      end else begin
        debug_4_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_7 = 1'b0;
    if(when_ArraySlice_l158_61) begin
      if(when_ArraySlice_l159_61) begin
        debug_5_7 = 1'b1;
      end else begin
        debug_5_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_61) begin
        debug_5_7 = 1'b1;
      end else begin
        debug_5_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_7 = 1'b0;
    if(when_ArraySlice_l158_62) begin
      if(when_ArraySlice_l159_62) begin
        debug_6_7 = 1'b1;
      end else begin
        debug_6_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_62) begin
        debug_6_7 = 1'b1;
      end else begin
        debug_6_7 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_7 = 1'b0;
    if(when_ArraySlice_l158_63) begin
      if(when_ArraySlice_l159_63) begin
        debug_7_7 = 1'b1;
      end else begin
        debug_7_7 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_63) begin
        debug_7_7 = 1'b1;
      end else begin
        debug_7_7 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_56 = (_zz_when_ArraySlice_l158_56 <= _zz_when_ArraySlice_l158_56_3);
  assign when_ArraySlice_l159_56 = (_zz_when_ArraySlice_l159_56 <= _zz_when_ArraySlice_l159_56_1);
  assign _zz_realValue_0_56 = (_zz__zz_realValue_0_56 % _zz__zz_realValue_0_56_1);
  assign when_ArraySlice_l110_56 = (_zz_realValue_0_56 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_56) begin
      realValue_0_56 = (_zz_realValue_0_56_1 - _zz_realValue_0_56);
    end else begin
      realValue_0_56 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_56 = (_zz_when_ArraySlice_l166_56 <= _zz_when_ArraySlice_l166_56_1);
  assign when_ArraySlice_l158_57 = (_zz_when_ArraySlice_l158_57 <= _zz_when_ArraySlice_l158_57_3);
  assign when_ArraySlice_l159_57 = (_zz_when_ArraySlice_l159_57 <= _zz_when_ArraySlice_l159_57_2);
  assign _zz_realValue_0_57 = (_zz__zz_realValue_0_57 % _zz__zz_realValue_0_57_1);
  assign when_ArraySlice_l110_57 = (_zz_realValue_0_57 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_57) begin
      realValue_0_57 = (_zz_realValue_0_57_1 - _zz_realValue_0_57);
    end else begin
      realValue_0_57 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_57 = (_zz_when_ArraySlice_l166_57 <= _zz_when_ArraySlice_l166_57_2);
  assign when_ArraySlice_l158_58 = (_zz_when_ArraySlice_l158_58 <= _zz_when_ArraySlice_l158_58_3);
  assign when_ArraySlice_l159_58 = (_zz_when_ArraySlice_l159_58 <= _zz_when_ArraySlice_l159_58_2);
  assign _zz_realValue_0_58 = (_zz__zz_realValue_0_58 % _zz__zz_realValue_0_58_1);
  assign when_ArraySlice_l110_58 = (_zz_realValue_0_58 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_58) begin
      realValue_0_58 = (_zz_realValue_0_58_1 - _zz_realValue_0_58);
    end else begin
      realValue_0_58 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_58 = (_zz_when_ArraySlice_l166_58 <= _zz_when_ArraySlice_l166_58_2);
  assign when_ArraySlice_l158_59 = (_zz_when_ArraySlice_l158_59 <= _zz_when_ArraySlice_l158_59_3);
  assign when_ArraySlice_l159_59 = (_zz_when_ArraySlice_l159_59 <= _zz_when_ArraySlice_l159_59_2);
  assign _zz_realValue_0_59 = (_zz__zz_realValue_0_59 % _zz__zz_realValue_0_59_1);
  assign when_ArraySlice_l110_59 = (_zz_realValue_0_59 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_59) begin
      realValue_0_59 = (_zz_realValue_0_59_1 - _zz_realValue_0_59);
    end else begin
      realValue_0_59 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_59 = (_zz_when_ArraySlice_l166_59 <= _zz_when_ArraySlice_l166_59_2);
  assign when_ArraySlice_l158_60 = (_zz_when_ArraySlice_l158_60 <= _zz_when_ArraySlice_l158_60_3);
  assign when_ArraySlice_l159_60 = (_zz_when_ArraySlice_l159_60 <= _zz_when_ArraySlice_l159_60_2);
  assign _zz_realValue_0_60 = (_zz__zz_realValue_0_60 % _zz__zz_realValue_0_60_1);
  assign when_ArraySlice_l110_60 = (_zz_realValue_0_60 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_60) begin
      realValue_0_60 = (_zz_realValue_0_60_1 - _zz_realValue_0_60);
    end else begin
      realValue_0_60 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_60 = (_zz_when_ArraySlice_l166_60 <= _zz_when_ArraySlice_l166_60_2);
  assign when_ArraySlice_l158_61 = (_zz_when_ArraySlice_l158_61 <= _zz_when_ArraySlice_l158_61_3);
  assign when_ArraySlice_l159_61 = (_zz_when_ArraySlice_l159_61 <= _zz_when_ArraySlice_l159_61_2);
  assign _zz_realValue_0_61 = (_zz__zz_realValue_0_61 % _zz__zz_realValue_0_61_1);
  assign when_ArraySlice_l110_61 = (_zz_realValue_0_61 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_61) begin
      realValue_0_61 = (_zz_realValue_0_61_1 - _zz_realValue_0_61);
    end else begin
      realValue_0_61 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_61 = (_zz_when_ArraySlice_l166_61 <= _zz_when_ArraySlice_l166_61_2);
  assign when_ArraySlice_l158_62 = (_zz_when_ArraySlice_l158_62 <= _zz_when_ArraySlice_l158_62_3);
  assign when_ArraySlice_l159_62 = (_zz_when_ArraySlice_l159_62 <= _zz_when_ArraySlice_l159_62_2);
  assign _zz_realValue_0_62 = (_zz__zz_realValue_0_62 % _zz__zz_realValue_0_62_1);
  assign when_ArraySlice_l110_62 = (_zz_realValue_0_62 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_62) begin
      realValue_0_62 = (_zz_realValue_0_62_1 - _zz_realValue_0_62);
    end else begin
      realValue_0_62 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_62 = (_zz_when_ArraySlice_l166_62 <= _zz_when_ArraySlice_l166_62_2);
  assign when_ArraySlice_l158_63 = (_zz_when_ArraySlice_l158_63 <= _zz_when_ArraySlice_l158_63_3);
  assign when_ArraySlice_l159_63 = (_zz_when_ArraySlice_l159_63 <= _zz_when_ArraySlice_l159_63_2);
  assign _zz_realValue_0_63 = (_zz__zz_realValue_0_63 % _zz__zz_realValue_0_63_1);
  assign when_ArraySlice_l110_63 = (_zz_realValue_0_63 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_63) begin
      realValue_0_63 = (_zz_realValue_0_63_1 - _zz_realValue_0_63);
    end else begin
      realValue_0_63 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_63 = (_zz_when_ArraySlice_l166_63 <= _zz_when_ArraySlice_l166_63_2);
  assign when_ArraySlice_l400_2 = (! ((((((_zz_when_ArraySlice_l400_2_1 && _zz_when_ArraySlice_l400_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_2_4 && _zz_when_ArraySlice_l400_2_5) && (debug_4_7 == _zz_when_ArraySlice_l400_2_6)) && (debug_5_7 == 1'b1)) && (debug_6_7 == 1'b1)) && (debug_7_7 == 1'b1))));
  assign when_ArraySlice_l403_2 = (_zz_when_ArraySlice_l403_2_1 <= _zz_when_ArraySlice_l403_2_2);
  assign when_ArraySlice_l406_2 = (_zz_when_ArraySlice_l406_2_1 <= _zz_when_ArraySlice_l406_2_2);
  assign when_ArraySlice_l413_2 = (_zz_when_ArraySlice_l413_2 == 13'h0);
  assign when_ArraySlice_l417_2 = (_zz_when_ArraySlice_l417_2_1 == 7'h0);
  assign outputStreamArrayData_2_fire_2 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l418_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l418_2_1) && outputStreamArrayData_2_fire_2);
  assign _zz_realValue1_0_7 = (_zz__zz_realValue1_0_7 % _zz__zz_realValue1_0_7_1);
  assign when_ArraySlice_l95_7 = (_zz_realValue1_0_7 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_7) begin
      realValue1_0_7 = (_zz_realValue1_0_7_1 - _zz_realValue1_0_7);
    end else begin
      realValue1_0_7 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_2 = (_zz_when_ArraySlice_l420_2_1 < _zz_when_ArraySlice_l420_2_3);
  always @(*) begin
    debug_0_8 = 1'b0;
    if(when_ArraySlice_l158_64) begin
      if(when_ArraySlice_l159_64) begin
        debug_0_8 = 1'b1;
      end else begin
        debug_0_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_64) begin
        debug_0_8 = 1'b1;
      end else begin
        debug_0_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_8 = 1'b0;
    if(when_ArraySlice_l158_65) begin
      if(when_ArraySlice_l159_65) begin
        debug_1_8 = 1'b1;
      end else begin
        debug_1_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_65) begin
        debug_1_8 = 1'b1;
      end else begin
        debug_1_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_8 = 1'b0;
    if(when_ArraySlice_l158_66) begin
      if(when_ArraySlice_l159_66) begin
        debug_2_8 = 1'b1;
      end else begin
        debug_2_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_66) begin
        debug_2_8 = 1'b1;
      end else begin
        debug_2_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_8 = 1'b0;
    if(when_ArraySlice_l158_67) begin
      if(when_ArraySlice_l159_67) begin
        debug_3_8 = 1'b1;
      end else begin
        debug_3_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_67) begin
        debug_3_8 = 1'b1;
      end else begin
        debug_3_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_8 = 1'b0;
    if(when_ArraySlice_l158_68) begin
      if(when_ArraySlice_l159_68) begin
        debug_4_8 = 1'b1;
      end else begin
        debug_4_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_68) begin
        debug_4_8 = 1'b1;
      end else begin
        debug_4_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_8 = 1'b0;
    if(when_ArraySlice_l158_69) begin
      if(when_ArraySlice_l159_69) begin
        debug_5_8 = 1'b1;
      end else begin
        debug_5_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_69) begin
        debug_5_8 = 1'b1;
      end else begin
        debug_5_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_8 = 1'b0;
    if(when_ArraySlice_l158_70) begin
      if(when_ArraySlice_l159_70) begin
        debug_6_8 = 1'b1;
      end else begin
        debug_6_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_70) begin
        debug_6_8 = 1'b1;
      end else begin
        debug_6_8 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_8 = 1'b0;
    if(when_ArraySlice_l158_71) begin
      if(when_ArraySlice_l159_71) begin
        debug_7_8 = 1'b1;
      end else begin
        debug_7_8 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_71) begin
        debug_7_8 = 1'b1;
      end else begin
        debug_7_8 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_64 = (_zz_when_ArraySlice_l158_64 <= _zz_when_ArraySlice_l158_64_3);
  assign when_ArraySlice_l159_64 = (_zz_when_ArraySlice_l159_64 <= _zz_when_ArraySlice_l159_64_1);
  assign _zz_realValue_0_64 = (_zz__zz_realValue_0_64 % _zz__zz_realValue_0_64_1);
  assign when_ArraySlice_l110_64 = (_zz_realValue_0_64 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_64) begin
      realValue_0_64 = (_zz_realValue_0_64_1 - _zz_realValue_0_64);
    end else begin
      realValue_0_64 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_64 = (_zz_when_ArraySlice_l166_64 <= _zz_when_ArraySlice_l166_64_1);
  assign when_ArraySlice_l158_65 = (_zz_when_ArraySlice_l158_65 <= _zz_when_ArraySlice_l158_65_3);
  assign when_ArraySlice_l159_65 = (_zz_when_ArraySlice_l159_65 <= _zz_when_ArraySlice_l159_65_2);
  assign _zz_realValue_0_65 = (_zz__zz_realValue_0_65 % _zz__zz_realValue_0_65_1);
  assign when_ArraySlice_l110_65 = (_zz_realValue_0_65 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_65) begin
      realValue_0_65 = (_zz_realValue_0_65_1 - _zz_realValue_0_65);
    end else begin
      realValue_0_65 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_65 = (_zz_when_ArraySlice_l166_65 <= _zz_when_ArraySlice_l166_65_2);
  assign when_ArraySlice_l158_66 = (_zz_when_ArraySlice_l158_66 <= _zz_when_ArraySlice_l158_66_3);
  assign when_ArraySlice_l159_66 = (_zz_when_ArraySlice_l159_66 <= _zz_when_ArraySlice_l159_66_2);
  assign _zz_realValue_0_66 = (_zz__zz_realValue_0_66 % _zz__zz_realValue_0_66_1);
  assign when_ArraySlice_l110_66 = (_zz_realValue_0_66 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_66) begin
      realValue_0_66 = (_zz_realValue_0_66_1 - _zz_realValue_0_66);
    end else begin
      realValue_0_66 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_66 = (_zz_when_ArraySlice_l166_66 <= _zz_when_ArraySlice_l166_66_2);
  assign when_ArraySlice_l158_67 = (_zz_when_ArraySlice_l158_67 <= _zz_when_ArraySlice_l158_67_3);
  assign when_ArraySlice_l159_67 = (_zz_when_ArraySlice_l159_67 <= _zz_when_ArraySlice_l159_67_2);
  assign _zz_realValue_0_67 = (_zz__zz_realValue_0_67 % _zz__zz_realValue_0_67_1);
  assign when_ArraySlice_l110_67 = (_zz_realValue_0_67 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_67) begin
      realValue_0_67 = (_zz_realValue_0_67_1 - _zz_realValue_0_67);
    end else begin
      realValue_0_67 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_67 = (_zz_when_ArraySlice_l166_67 <= _zz_when_ArraySlice_l166_67_2);
  assign when_ArraySlice_l158_68 = (_zz_when_ArraySlice_l158_68 <= _zz_when_ArraySlice_l158_68_3);
  assign when_ArraySlice_l159_68 = (_zz_when_ArraySlice_l159_68 <= _zz_when_ArraySlice_l159_68_2);
  assign _zz_realValue_0_68 = (_zz__zz_realValue_0_68 % _zz__zz_realValue_0_68_1);
  assign when_ArraySlice_l110_68 = (_zz_realValue_0_68 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_68) begin
      realValue_0_68 = (_zz_realValue_0_68_1 - _zz_realValue_0_68);
    end else begin
      realValue_0_68 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_68 = (_zz_when_ArraySlice_l166_68 <= _zz_when_ArraySlice_l166_68_2);
  assign when_ArraySlice_l158_69 = (_zz_when_ArraySlice_l158_69 <= _zz_when_ArraySlice_l158_69_3);
  assign when_ArraySlice_l159_69 = (_zz_when_ArraySlice_l159_69 <= _zz_when_ArraySlice_l159_69_2);
  assign _zz_realValue_0_69 = (_zz__zz_realValue_0_69 % _zz__zz_realValue_0_69_1);
  assign when_ArraySlice_l110_69 = (_zz_realValue_0_69 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_69) begin
      realValue_0_69 = (_zz_realValue_0_69_1 - _zz_realValue_0_69);
    end else begin
      realValue_0_69 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_69 = (_zz_when_ArraySlice_l166_69 <= _zz_when_ArraySlice_l166_69_2);
  assign when_ArraySlice_l158_70 = (_zz_when_ArraySlice_l158_70 <= _zz_when_ArraySlice_l158_70_3);
  assign when_ArraySlice_l159_70 = (_zz_when_ArraySlice_l159_70 <= _zz_when_ArraySlice_l159_70_2);
  assign _zz_realValue_0_70 = (_zz__zz_realValue_0_70 % _zz__zz_realValue_0_70_1);
  assign when_ArraySlice_l110_70 = (_zz_realValue_0_70 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_70) begin
      realValue_0_70 = (_zz_realValue_0_70_1 - _zz_realValue_0_70);
    end else begin
      realValue_0_70 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_70 = (_zz_when_ArraySlice_l166_70 <= _zz_when_ArraySlice_l166_70_2);
  assign when_ArraySlice_l158_71 = (_zz_when_ArraySlice_l158_71 <= _zz_when_ArraySlice_l158_71_3);
  assign when_ArraySlice_l159_71 = (_zz_when_ArraySlice_l159_71 <= _zz_when_ArraySlice_l159_71_2);
  assign _zz_realValue_0_71 = (_zz__zz_realValue_0_71 % _zz__zz_realValue_0_71_1);
  assign when_ArraySlice_l110_71 = (_zz_realValue_0_71 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_71) begin
      realValue_0_71 = (_zz_realValue_0_71_1 - _zz_realValue_0_71);
    end else begin
      realValue_0_71 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_71 = (_zz_when_ArraySlice_l166_71 <= _zz_when_ArraySlice_l166_71_2);
  assign when_ArraySlice_l425_2 = (! ((((((_zz_when_ArraySlice_l425_2_1 && _zz_when_ArraySlice_l425_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l425_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_2_4 && _zz_when_ArraySlice_l425_2_5) && (debug_4_8 == _zz_when_ArraySlice_l425_2_6)) && (debug_5_8 == 1'b1)) && (debug_6_8 == 1'b1)) && (debug_7_8 == 1'b1))));
  assign when_ArraySlice_l428_2 = (_zz_when_ArraySlice_l428_2_1 <= _zz_when_ArraySlice_l428_2_2);
  assign when_ArraySlice_l431_2 = (_zz_when_ArraySlice_l431_2_1 <= _zz_when_ArraySlice_l431_2_2);
  assign outputStreamArrayData_2_fire_3 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l438_2 = ((_zz_when_ArraySlice_l438_2 == 13'h0) && outputStreamArrayData_2_fire_3);
  assign outputStreamArrayData_2_fire_4 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l449_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l449_2_1) && outputStreamArrayData_2_fire_4);
  assign _zz_realValue1_0_8 = (_zz__zz_realValue1_0_8 % _zz__zz_realValue1_0_8_1);
  assign when_ArraySlice_l95_8 = (_zz_realValue1_0_8 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_8) begin
      realValue1_0_8 = (_zz_realValue1_0_8_1 - _zz_realValue1_0_8);
    end else begin
      realValue1_0_8 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_2 = (_zz_when_ArraySlice_l450_2_1 < _zz_when_ArraySlice_l450_2_3);
  always @(*) begin
    debug_0_9 = 1'b0;
    if(when_ArraySlice_l158_72) begin
      if(when_ArraySlice_l159_72) begin
        debug_0_9 = 1'b1;
      end else begin
        debug_0_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_72) begin
        debug_0_9 = 1'b1;
      end else begin
        debug_0_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_9 = 1'b0;
    if(when_ArraySlice_l158_73) begin
      if(when_ArraySlice_l159_73) begin
        debug_1_9 = 1'b1;
      end else begin
        debug_1_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_73) begin
        debug_1_9 = 1'b1;
      end else begin
        debug_1_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_9 = 1'b0;
    if(when_ArraySlice_l158_74) begin
      if(when_ArraySlice_l159_74) begin
        debug_2_9 = 1'b1;
      end else begin
        debug_2_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_74) begin
        debug_2_9 = 1'b1;
      end else begin
        debug_2_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_9 = 1'b0;
    if(when_ArraySlice_l158_75) begin
      if(when_ArraySlice_l159_75) begin
        debug_3_9 = 1'b1;
      end else begin
        debug_3_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_75) begin
        debug_3_9 = 1'b1;
      end else begin
        debug_3_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_9 = 1'b0;
    if(when_ArraySlice_l158_76) begin
      if(when_ArraySlice_l159_76) begin
        debug_4_9 = 1'b1;
      end else begin
        debug_4_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_76) begin
        debug_4_9 = 1'b1;
      end else begin
        debug_4_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_9 = 1'b0;
    if(when_ArraySlice_l158_77) begin
      if(when_ArraySlice_l159_77) begin
        debug_5_9 = 1'b1;
      end else begin
        debug_5_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_77) begin
        debug_5_9 = 1'b1;
      end else begin
        debug_5_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_9 = 1'b0;
    if(when_ArraySlice_l158_78) begin
      if(when_ArraySlice_l159_78) begin
        debug_6_9 = 1'b1;
      end else begin
        debug_6_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_78) begin
        debug_6_9 = 1'b1;
      end else begin
        debug_6_9 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_9 = 1'b0;
    if(when_ArraySlice_l158_79) begin
      if(when_ArraySlice_l159_79) begin
        debug_7_9 = 1'b1;
      end else begin
        debug_7_9 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_79) begin
        debug_7_9 = 1'b1;
      end else begin
        debug_7_9 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_72 = (_zz_when_ArraySlice_l158_72 <= _zz_when_ArraySlice_l158_72_3);
  assign when_ArraySlice_l159_72 = (_zz_when_ArraySlice_l159_72 <= _zz_when_ArraySlice_l159_72_1);
  assign _zz_realValue_0_72 = (_zz__zz_realValue_0_72 % _zz__zz_realValue_0_72_1);
  assign when_ArraySlice_l110_72 = (_zz_realValue_0_72 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_72) begin
      realValue_0_72 = (_zz_realValue_0_72_1 - _zz_realValue_0_72);
    end else begin
      realValue_0_72 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_72 = (_zz_when_ArraySlice_l166_72 <= _zz_when_ArraySlice_l166_72_1);
  assign when_ArraySlice_l158_73 = (_zz_when_ArraySlice_l158_73 <= _zz_when_ArraySlice_l158_73_3);
  assign when_ArraySlice_l159_73 = (_zz_when_ArraySlice_l159_73 <= _zz_when_ArraySlice_l159_73_2);
  assign _zz_realValue_0_73 = (_zz__zz_realValue_0_73 % _zz__zz_realValue_0_73_1);
  assign when_ArraySlice_l110_73 = (_zz_realValue_0_73 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_73) begin
      realValue_0_73 = (_zz_realValue_0_73_1 - _zz_realValue_0_73);
    end else begin
      realValue_0_73 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_73 = (_zz_when_ArraySlice_l166_73 <= _zz_when_ArraySlice_l166_73_2);
  assign when_ArraySlice_l158_74 = (_zz_when_ArraySlice_l158_74 <= _zz_when_ArraySlice_l158_74_3);
  assign when_ArraySlice_l159_74 = (_zz_when_ArraySlice_l159_74 <= _zz_when_ArraySlice_l159_74_2);
  assign _zz_realValue_0_74 = (_zz__zz_realValue_0_74 % _zz__zz_realValue_0_74_1);
  assign when_ArraySlice_l110_74 = (_zz_realValue_0_74 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_74) begin
      realValue_0_74 = (_zz_realValue_0_74_1 - _zz_realValue_0_74);
    end else begin
      realValue_0_74 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_74 = (_zz_when_ArraySlice_l166_74 <= _zz_when_ArraySlice_l166_74_2);
  assign when_ArraySlice_l158_75 = (_zz_when_ArraySlice_l158_75 <= _zz_when_ArraySlice_l158_75_3);
  assign when_ArraySlice_l159_75 = (_zz_when_ArraySlice_l159_75 <= _zz_when_ArraySlice_l159_75_2);
  assign _zz_realValue_0_75 = (_zz__zz_realValue_0_75 % _zz__zz_realValue_0_75_1);
  assign when_ArraySlice_l110_75 = (_zz_realValue_0_75 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_75) begin
      realValue_0_75 = (_zz_realValue_0_75_1 - _zz_realValue_0_75);
    end else begin
      realValue_0_75 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_75 = (_zz_when_ArraySlice_l166_75 <= _zz_when_ArraySlice_l166_75_2);
  assign when_ArraySlice_l158_76 = (_zz_when_ArraySlice_l158_76 <= _zz_when_ArraySlice_l158_76_3);
  assign when_ArraySlice_l159_76 = (_zz_when_ArraySlice_l159_76 <= _zz_when_ArraySlice_l159_76_2);
  assign _zz_realValue_0_76 = (_zz__zz_realValue_0_76 % _zz__zz_realValue_0_76_1);
  assign when_ArraySlice_l110_76 = (_zz_realValue_0_76 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_76) begin
      realValue_0_76 = (_zz_realValue_0_76_1 - _zz_realValue_0_76);
    end else begin
      realValue_0_76 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_76 = (_zz_when_ArraySlice_l166_76 <= _zz_when_ArraySlice_l166_76_2);
  assign when_ArraySlice_l158_77 = (_zz_when_ArraySlice_l158_77 <= _zz_when_ArraySlice_l158_77_3);
  assign when_ArraySlice_l159_77 = (_zz_when_ArraySlice_l159_77 <= _zz_when_ArraySlice_l159_77_2);
  assign _zz_realValue_0_77 = (_zz__zz_realValue_0_77 % _zz__zz_realValue_0_77_1);
  assign when_ArraySlice_l110_77 = (_zz_realValue_0_77 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_77) begin
      realValue_0_77 = (_zz_realValue_0_77_1 - _zz_realValue_0_77);
    end else begin
      realValue_0_77 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_77 = (_zz_when_ArraySlice_l166_77 <= _zz_when_ArraySlice_l166_77_2);
  assign when_ArraySlice_l158_78 = (_zz_when_ArraySlice_l158_78 <= _zz_when_ArraySlice_l158_78_3);
  assign when_ArraySlice_l159_78 = (_zz_when_ArraySlice_l159_78 <= _zz_when_ArraySlice_l159_78_2);
  assign _zz_realValue_0_78 = (_zz__zz_realValue_0_78 % _zz__zz_realValue_0_78_1);
  assign when_ArraySlice_l110_78 = (_zz_realValue_0_78 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_78) begin
      realValue_0_78 = (_zz_realValue_0_78_1 - _zz_realValue_0_78);
    end else begin
      realValue_0_78 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_78 = (_zz_when_ArraySlice_l166_78 <= _zz_when_ArraySlice_l166_78_2);
  assign when_ArraySlice_l158_79 = (_zz_when_ArraySlice_l158_79 <= _zz_when_ArraySlice_l158_79_3);
  assign when_ArraySlice_l159_79 = (_zz_when_ArraySlice_l159_79 <= _zz_when_ArraySlice_l159_79_2);
  assign _zz_realValue_0_79 = (_zz__zz_realValue_0_79 % _zz__zz_realValue_0_79_1);
  assign when_ArraySlice_l110_79 = (_zz_realValue_0_79 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_79) begin
      realValue_0_79 = (_zz_realValue_0_79_1 - _zz_realValue_0_79);
    end else begin
      realValue_0_79 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_79 = (_zz_when_ArraySlice_l166_79 <= _zz_when_ArraySlice_l166_79_2);
  assign when_ArraySlice_l457_2 = (! ((((((_zz_when_ArraySlice_l457_2_1 && _zz_when_ArraySlice_l457_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l457_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_2_4 && _zz_when_ArraySlice_l457_2_5) && (debug_4_9 == _zz_when_ArraySlice_l457_2_6)) && (debug_5_9 == 1'b1)) && (debug_6_9 == 1'b1)) && (debug_7_9 == 1'b1))));
  assign outputStreamArrayData_2_fire_5 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l461_2 = ((_zz_when_ArraySlice_l461_2 == 13'h0) && outputStreamArrayData_2_fire_5);
  assign when_ArraySlice_l447_2 = (allowPadding_2 && (_zz_when_ArraySlice_l447_2_1 <= _zz_when_ArraySlice_l447_2_2));
  assign outputStreamArrayData_2_fire_6 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l468_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l468_2_1);
  assign when_ArraySlice_l376_3 = (_zz_when_ArraySlice_l376_3_1 < _zz_when_ArraySlice_l376_3_4);
  assign when_ArraySlice_l377_3 = ((! holdReadOp_3) && (_zz_when_ArraySlice_l377_3_1 != 7'h0));
  assign _zz_outputStreamArrayData_3_valid = (selectReadFifo_3 + _zz__zz_outputStreamArrayData_3_valid);
  assign _zz_6 = ({127'd0,1'b1} <<< _zz__zz_6);
  assign _zz_io_pop_ready_3 = outputStreamArrayData_3_ready;
  assign when_ArraySlice_l382_3 = (! holdReadOp_3);
  assign outputStreamArrayData_3_fire = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l383_3 = ((7'h01 < _zz_when_ArraySlice_l383_3_1) && outputStreamArrayData_3_fire);
  assign when_ArraySlice_l384_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l384_3);
  assign when_ArraySlice_l387_3 = (_zz_when_ArraySlice_l387_3 == 13'h0);
  assign outputStreamArrayData_3_fire_1 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l392_3 = ((_zz_when_ArraySlice_l392_3_1 == 7'h01) && outputStreamArrayData_3_fire_1);
  assign when_ArraySlice_l393_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l393_3);
  assign _zz_realValue1_0_9 = (_zz__zz_realValue1_0_9 % _zz__zz_realValue1_0_9_1);
  assign when_ArraySlice_l95_9 = (_zz_realValue1_0_9 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_9) begin
      realValue1_0_9 = (_zz_realValue1_0_9_1 - _zz_realValue1_0_9);
    end else begin
      realValue1_0_9 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_3 = (_zz_when_ArraySlice_l395_3 < _zz_when_ArraySlice_l395_3_2);
  always @(*) begin
    debug_0_10 = 1'b0;
    if(when_ArraySlice_l158_80) begin
      if(when_ArraySlice_l159_80) begin
        debug_0_10 = 1'b1;
      end else begin
        debug_0_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_80) begin
        debug_0_10 = 1'b1;
      end else begin
        debug_0_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_10 = 1'b0;
    if(when_ArraySlice_l158_81) begin
      if(when_ArraySlice_l159_81) begin
        debug_1_10 = 1'b1;
      end else begin
        debug_1_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_81) begin
        debug_1_10 = 1'b1;
      end else begin
        debug_1_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_10 = 1'b0;
    if(when_ArraySlice_l158_82) begin
      if(when_ArraySlice_l159_82) begin
        debug_2_10 = 1'b1;
      end else begin
        debug_2_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_82) begin
        debug_2_10 = 1'b1;
      end else begin
        debug_2_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_10 = 1'b0;
    if(when_ArraySlice_l158_83) begin
      if(when_ArraySlice_l159_83) begin
        debug_3_10 = 1'b1;
      end else begin
        debug_3_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_83) begin
        debug_3_10 = 1'b1;
      end else begin
        debug_3_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_10 = 1'b0;
    if(when_ArraySlice_l158_84) begin
      if(when_ArraySlice_l159_84) begin
        debug_4_10 = 1'b1;
      end else begin
        debug_4_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_84) begin
        debug_4_10 = 1'b1;
      end else begin
        debug_4_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_10 = 1'b0;
    if(when_ArraySlice_l158_85) begin
      if(when_ArraySlice_l159_85) begin
        debug_5_10 = 1'b1;
      end else begin
        debug_5_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_85) begin
        debug_5_10 = 1'b1;
      end else begin
        debug_5_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_10 = 1'b0;
    if(when_ArraySlice_l158_86) begin
      if(when_ArraySlice_l159_86) begin
        debug_6_10 = 1'b1;
      end else begin
        debug_6_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_86) begin
        debug_6_10 = 1'b1;
      end else begin
        debug_6_10 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_10 = 1'b0;
    if(when_ArraySlice_l158_87) begin
      if(when_ArraySlice_l159_87) begin
        debug_7_10 = 1'b1;
      end else begin
        debug_7_10 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_87) begin
        debug_7_10 = 1'b1;
      end else begin
        debug_7_10 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_80 = (_zz_when_ArraySlice_l158_80 <= _zz_when_ArraySlice_l158_80_3);
  assign when_ArraySlice_l159_80 = (_zz_when_ArraySlice_l159_80 <= _zz_when_ArraySlice_l159_80_1);
  assign _zz_realValue_0_80 = (_zz__zz_realValue_0_80 % _zz__zz_realValue_0_80_1);
  assign when_ArraySlice_l110_80 = (_zz_realValue_0_80 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_80) begin
      realValue_0_80 = (_zz_realValue_0_80_1 - _zz_realValue_0_80);
    end else begin
      realValue_0_80 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_80 = (_zz_when_ArraySlice_l166_80 <= _zz_when_ArraySlice_l166_80_1);
  assign when_ArraySlice_l158_81 = (_zz_when_ArraySlice_l158_81 <= _zz_when_ArraySlice_l158_81_3);
  assign when_ArraySlice_l159_81 = (_zz_when_ArraySlice_l159_81 <= _zz_when_ArraySlice_l159_81_2);
  assign _zz_realValue_0_81 = (_zz__zz_realValue_0_81 % _zz__zz_realValue_0_81_1);
  assign when_ArraySlice_l110_81 = (_zz_realValue_0_81 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_81) begin
      realValue_0_81 = (_zz_realValue_0_81_1 - _zz_realValue_0_81);
    end else begin
      realValue_0_81 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_81 = (_zz_when_ArraySlice_l166_81 <= _zz_when_ArraySlice_l166_81_2);
  assign when_ArraySlice_l158_82 = (_zz_when_ArraySlice_l158_82 <= _zz_when_ArraySlice_l158_82_3);
  assign when_ArraySlice_l159_82 = (_zz_when_ArraySlice_l159_82 <= _zz_when_ArraySlice_l159_82_2);
  assign _zz_realValue_0_82 = (_zz__zz_realValue_0_82 % _zz__zz_realValue_0_82_1);
  assign when_ArraySlice_l110_82 = (_zz_realValue_0_82 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_82) begin
      realValue_0_82 = (_zz_realValue_0_82_1 - _zz_realValue_0_82);
    end else begin
      realValue_0_82 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_82 = (_zz_when_ArraySlice_l166_82 <= _zz_when_ArraySlice_l166_82_2);
  assign when_ArraySlice_l158_83 = (_zz_when_ArraySlice_l158_83 <= _zz_when_ArraySlice_l158_83_3);
  assign when_ArraySlice_l159_83 = (_zz_when_ArraySlice_l159_83 <= _zz_when_ArraySlice_l159_83_2);
  assign _zz_realValue_0_83 = (_zz__zz_realValue_0_83 % _zz__zz_realValue_0_83_1);
  assign when_ArraySlice_l110_83 = (_zz_realValue_0_83 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_83) begin
      realValue_0_83 = (_zz_realValue_0_83_1 - _zz_realValue_0_83);
    end else begin
      realValue_0_83 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_83 = (_zz_when_ArraySlice_l166_83 <= _zz_when_ArraySlice_l166_83_2);
  assign when_ArraySlice_l158_84 = (_zz_when_ArraySlice_l158_84 <= _zz_when_ArraySlice_l158_84_3);
  assign when_ArraySlice_l159_84 = (_zz_when_ArraySlice_l159_84 <= _zz_when_ArraySlice_l159_84_2);
  assign _zz_realValue_0_84 = (_zz__zz_realValue_0_84 % _zz__zz_realValue_0_84_1);
  assign when_ArraySlice_l110_84 = (_zz_realValue_0_84 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_84) begin
      realValue_0_84 = (_zz_realValue_0_84_1 - _zz_realValue_0_84);
    end else begin
      realValue_0_84 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_84 = (_zz_when_ArraySlice_l166_84 <= _zz_when_ArraySlice_l166_84_2);
  assign when_ArraySlice_l158_85 = (_zz_when_ArraySlice_l158_85 <= _zz_when_ArraySlice_l158_85_3);
  assign when_ArraySlice_l159_85 = (_zz_when_ArraySlice_l159_85 <= _zz_when_ArraySlice_l159_85_2);
  assign _zz_realValue_0_85 = (_zz__zz_realValue_0_85 % _zz__zz_realValue_0_85_1);
  assign when_ArraySlice_l110_85 = (_zz_realValue_0_85 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_85) begin
      realValue_0_85 = (_zz_realValue_0_85_1 - _zz_realValue_0_85);
    end else begin
      realValue_0_85 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_85 = (_zz_when_ArraySlice_l166_85 <= _zz_when_ArraySlice_l166_85_2);
  assign when_ArraySlice_l158_86 = (_zz_when_ArraySlice_l158_86 <= _zz_when_ArraySlice_l158_86_3);
  assign when_ArraySlice_l159_86 = (_zz_when_ArraySlice_l159_86 <= _zz_when_ArraySlice_l159_86_2);
  assign _zz_realValue_0_86 = (_zz__zz_realValue_0_86 % _zz__zz_realValue_0_86_1);
  assign when_ArraySlice_l110_86 = (_zz_realValue_0_86 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_86) begin
      realValue_0_86 = (_zz_realValue_0_86_1 - _zz_realValue_0_86);
    end else begin
      realValue_0_86 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_86 = (_zz_when_ArraySlice_l166_86 <= _zz_when_ArraySlice_l166_86_2);
  assign when_ArraySlice_l158_87 = (_zz_when_ArraySlice_l158_87 <= _zz_when_ArraySlice_l158_87_3);
  assign when_ArraySlice_l159_87 = (_zz_when_ArraySlice_l159_87 <= _zz_when_ArraySlice_l159_87_2);
  assign _zz_realValue_0_87 = (_zz__zz_realValue_0_87 % _zz__zz_realValue_0_87_1);
  assign when_ArraySlice_l110_87 = (_zz_realValue_0_87 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_87) begin
      realValue_0_87 = (_zz_realValue_0_87_1 - _zz_realValue_0_87);
    end else begin
      realValue_0_87 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_87 = (_zz_when_ArraySlice_l166_87 <= _zz_when_ArraySlice_l166_87_2);
  assign when_ArraySlice_l400_3 = (! ((((((_zz_when_ArraySlice_l400_3_1 && _zz_when_ArraySlice_l400_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_3_4 && _zz_when_ArraySlice_l400_3_5) && (debug_4_10 == _zz_when_ArraySlice_l400_3_6)) && (debug_5_10 == 1'b1)) && (debug_6_10 == 1'b1)) && (debug_7_10 == 1'b1))));
  assign when_ArraySlice_l403_3 = (_zz_when_ArraySlice_l403_3_1 <= _zz_when_ArraySlice_l403_3_2);
  assign when_ArraySlice_l406_3 = (_zz_when_ArraySlice_l406_3_1 <= _zz_when_ArraySlice_l406_3_2);
  assign when_ArraySlice_l413_3 = (_zz_when_ArraySlice_l413_3 == 13'h0);
  assign when_ArraySlice_l417_3 = (_zz_when_ArraySlice_l417_3_1 == 7'h0);
  assign outputStreamArrayData_3_fire_2 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l418_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l418_3_1) && outputStreamArrayData_3_fire_2);
  assign _zz_realValue1_0_10 = (_zz__zz_realValue1_0_10 % _zz__zz_realValue1_0_10_1);
  assign when_ArraySlice_l95_10 = (_zz_realValue1_0_10 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_10) begin
      realValue1_0_10 = (_zz_realValue1_0_10_1 - _zz_realValue1_0_10);
    end else begin
      realValue1_0_10 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_3 = (_zz_when_ArraySlice_l420_3 < _zz_when_ArraySlice_l420_3_2);
  always @(*) begin
    debug_0_11 = 1'b0;
    if(when_ArraySlice_l158_88) begin
      if(when_ArraySlice_l159_88) begin
        debug_0_11 = 1'b1;
      end else begin
        debug_0_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_88) begin
        debug_0_11 = 1'b1;
      end else begin
        debug_0_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_11 = 1'b0;
    if(when_ArraySlice_l158_89) begin
      if(when_ArraySlice_l159_89) begin
        debug_1_11 = 1'b1;
      end else begin
        debug_1_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_89) begin
        debug_1_11 = 1'b1;
      end else begin
        debug_1_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_11 = 1'b0;
    if(when_ArraySlice_l158_90) begin
      if(when_ArraySlice_l159_90) begin
        debug_2_11 = 1'b1;
      end else begin
        debug_2_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_90) begin
        debug_2_11 = 1'b1;
      end else begin
        debug_2_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_11 = 1'b0;
    if(when_ArraySlice_l158_91) begin
      if(when_ArraySlice_l159_91) begin
        debug_3_11 = 1'b1;
      end else begin
        debug_3_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_91) begin
        debug_3_11 = 1'b1;
      end else begin
        debug_3_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_11 = 1'b0;
    if(when_ArraySlice_l158_92) begin
      if(when_ArraySlice_l159_92) begin
        debug_4_11 = 1'b1;
      end else begin
        debug_4_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_92) begin
        debug_4_11 = 1'b1;
      end else begin
        debug_4_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_11 = 1'b0;
    if(when_ArraySlice_l158_93) begin
      if(when_ArraySlice_l159_93) begin
        debug_5_11 = 1'b1;
      end else begin
        debug_5_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_93) begin
        debug_5_11 = 1'b1;
      end else begin
        debug_5_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_11 = 1'b0;
    if(when_ArraySlice_l158_94) begin
      if(when_ArraySlice_l159_94) begin
        debug_6_11 = 1'b1;
      end else begin
        debug_6_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_94) begin
        debug_6_11 = 1'b1;
      end else begin
        debug_6_11 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_11 = 1'b0;
    if(when_ArraySlice_l158_95) begin
      if(when_ArraySlice_l159_95) begin
        debug_7_11 = 1'b1;
      end else begin
        debug_7_11 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_95) begin
        debug_7_11 = 1'b1;
      end else begin
        debug_7_11 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_88 = (_zz_when_ArraySlice_l158_88 <= _zz_when_ArraySlice_l158_88_3);
  assign when_ArraySlice_l159_88 = (_zz_when_ArraySlice_l159_88 <= _zz_when_ArraySlice_l159_88_1);
  assign _zz_realValue_0_88 = (_zz__zz_realValue_0_88 % _zz__zz_realValue_0_88_1);
  assign when_ArraySlice_l110_88 = (_zz_realValue_0_88 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_88) begin
      realValue_0_88 = (_zz_realValue_0_88_1 - _zz_realValue_0_88);
    end else begin
      realValue_0_88 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_88 = (_zz_when_ArraySlice_l166_88 <= _zz_when_ArraySlice_l166_88_1);
  assign when_ArraySlice_l158_89 = (_zz_when_ArraySlice_l158_89 <= _zz_when_ArraySlice_l158_89_3);
  assign when_ArraySlice_l159_89 = (_zz_when_ArraySlice_l159_89 <= _zz_when_ArraySlice_l159_89_2);
  assign _zz_realValue_0_89 = (_zz__zz_realValue_0_89 % _zz__zz_realValue_0_89_1);
  assign when_ArraySlice_l110_89 = (_zz_realValue_0_89 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_89) begin
      realValue_0_89 = (_zz_realValue_0_89_1 - _zz_realValue_0_89);
    end else begin
      realValue_0_89 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_89 = (_zz_when_ArraySlice_l166_89 <= _zz_when_ArraySlice_l166_89_2);
  assign when_ArraySlice_l158_90 = (_zz_when_ArraySlice_l158_90 <= _zz_when_ArraySlice_l158_90_3);
  assign when_ArraySlice_l159_90 = (_zz_when_ArraySlice_l159_90 <= _zz_when_ArraySlice_l159_90_2);
  assign _zz_realValue_0_90 = (_zz__zz_realValue_0_90 % _zz__zz_realValue_0_90_1);
  assign when_ArraySlice_l110_90 = (_zz_realValue_0_90 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_90) begin
      realValue_0_90 = (_zz_realValue_0_90_1 - _zz_realValue_0_90);
    end else begin
      realValue_0_90 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_90 = (_zz_when_ArraySlice_l166_90 <= _zz_when_ArraySlice_l166_90_2);
  assign when_ArraySlice_l158_91 = (_zz_when_ArraySlice_l158_91 <= _zz_when_ArraySlice_l158_91_3);
  assign when_ArraySlice_l159_91 = (_zz_when_ArraySlice_l159_91 <= _zz_when_ArraySlice_l159_91_2);
  assign _zz_realValue_0_91 = (_zz__zz_realValue_0_91 % _zz__zz_realValue_0_91_1);
  assign when_ArraySlice_l110_91 = (_zz_realValue_0_91 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_91) begin
      realValue_0_91 = (_zz_realValue_0_91_1 - _zz_realValue_0_91);
    end else begin
      realValue_0_91 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_91 = (_zz_when_ArraySlice_l166_91 <= _zz_when_ArraySlice_l166_91_2);
  assign when_ArraySlice_l158_92 = (_zz_when_ArraySlice_l158_92 <= _zz_when_ArraySlice_l158_92_3);
  assign when_ArraySlice_l159_92 = (_zz_when_ArraySlice_l159_92 <= _zz_when_ArraySlice_l159_92_2);
  assign _zz_realValue_0_92 = (_zz__zz_realValue_0_92 % _zz__zz_realValue_0_92_1);
  assign when_ArraySlice_l110_92 = (_zz_realValue_0_92 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_92) begin
      realValue_0_92 = (_zz_realValue_0_92_1 - _zz_realValue_0_92);
    end else begin
      realValue_0_92 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_92 = (_zz_when_ArraySlice_l166_92 <= _zz_when_ArraySlice_l166_92_2);
  assign when_ArraySlice_l158_93 = (_zz_when_ArraySlice_l158_93 <= _zz_when_ArraySlice_l158_93_3);
  assign when_ArraySlice_l159_93 = (_zz_when_ArraySlice_l159_93 <= _zz_when_ArraySlice_l159_93_2);
  assign _zz_realValue_0_93 = (_zz__zz_realValue_0_93 % _zz__zz_realValue_0_93_1);
  assign when_ArraySlice_l110_93 = (_zz_realValue_0_93 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_93) begin
      realValue_0_93 = (_zz_realValue_0_93_1 - _zz_realValue_0_93);
    end else begin
      realValue_0_93 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_93 = (_zz_when_ArraySlice_l166_93 <= _zz_when_ArraySlice_l166_93_2);
  assign when_ArraySlice_l158_94 = (_zz_when_ArraySlice_l158_94 <= _zz_when_ArraySlice_l158_94_3);
  assign when_ArraySlice_l159_94 = (_zz_when_ArraySlice_l159_94 <= _zz_when_ArraySlice_l159_94_2);
  assign _zz_realValue_0_94 = (_zz__zz_realValue_0_94 % _zz__zz_realValue_0_94_1);
  assign when_ArraySlice_l110_94 = (_zz_realValue_0_94 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_94) begin
      realValue_0_94 = (_zz_realValue_0_94_1 - _zz_realValue_0_94);
    end else begin
      realValue_0_94 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_94 = (_zz_when_ArraySlice_l166_94 <= _zz_when_ArraySlice_l166_94_2);
  assign when_ArraySlice_l158_95 = (_zz_when_ArraySlice_l158_95 <= _zz_when_ArraySlice_l158_95_3);
  assign when_ArraySlice_l159_95 = (_zz_when_ArraySlice_l159_95 <= _zz_when_ArraySlice_l159_95_2);
  assign _zz_realValue_0_95 = (_zz__zz_realValue_0_95 % _zz__zz_realValue_0_95_1);
  assign when_ArraySlice_l110_95 = (_zz_realValue_0_95 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_95) begin
      realValue_0_95 = (_zz_realValue_0_95_1 - _zz_realValue_0_95);
    end else begin
      realValue_0_95 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_95 = (_zz_when_ArraySlice_l166_95 <= _zz_when_ArraySlice_l166_95_2);
  assign when_ArraySlice_l425_3 = (! ((((((_zz_when_ArraySlice_l425_3_1 && _zz_when_ArraySlice_l425_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l425_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_3_4 && _zz_when_ArraySlice_l425_3_5) && (debug_4_11 == _zz_when_ArraySlice_l425_3_6)) && (debug_5_11 == 1'b1)) && (debug_6_11 == 1'b1)) && (debug_7_11 == 1'b1))));
  assign when_ArraySlice_l428_3 = (_zz_when_ArraySlice_l428_3_1 <= _zz_when_ArraySlice_l428_3_2);
  assign when_ArraySlice_l431_3 = (_zz_when_ArraySlice_l431_3_1 <= _zz_when_ArraySlice_l431_3_2);
  assign outputStreamArrayData_3_fire_3 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l438_3 = ((_zz_when_ArraySlice_l438_3 == 13'h0) && outputStreamArrayData_3_fire_3);
  assign outputStreamArrayData_3_fire_4 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l449_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l449_3) && outputStreamArrayData_3_fire_4);
  assign _zz_realValue1_0_11 = (_zz__zz_realValue1_0_11 % _zz__zz_realValue1_0_11_1);
  assign when_ArraySlice_l95_11 = (_zz_realValue1_0_11 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_11) begin
      realValue1_0_11 = (_zz_realValue1_0_11_1 - _zz_realValue1_0_11);
    end else begin
      realValue1_0_11 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_3 = (_zz_when_ArraySlice_l450_3 < _zz_when_ArraySlice_l450_3_2);
  always @(*) begin
    debug_0_12 = 1'b0;
    if(when_ArraySlice_l158_96) begin
      if(when_ArraySlice_l159_96) begin
        debug_0_12 = 1'b1;
      end else begin
        debug_0_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_96) begin
        debug_0_12 = 1'b1;
      end else begin
        debug_0_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_12 = 1'b0;
    if(when_ArraySlice_l158_97) begin
      if(when_ArraySlice_l159_97) begin
        debug_1_12 = 1'b1;
      end else begin
        debug_1_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_97) begin
        debug_1_12 = 1'b1;
      end else begin
        debug_1_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_12 = 1'b0;
    if(when_ArraySlice_l158_98) begin
      if(when_ArraySlice_l159_98) begin
        debug_2_12 = 1'b1;
      end else begin
        debug_2_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_98) begin
        debug_2_12 = 1'b1;
      end else begin
        debug_2_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_12 = 1'b0;
    if(when_ArraySlice_l158_99) begin
      if(when_ArraySlice_l159_99) begin
        debug_3_12 = 1'b1;
      end else begin
        debug_3_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_99) begin
        debug_3_12 = 1'b1;
      end else begin
        debug_3_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_12 = 1'b0;
    if(when_ArraySlice_l158_100) begin
      if(when_ArraySlice_l159_100) begin
        debug_4_12 = 1'b1;
      end else begin
        debug_4_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_100) begin
        debug_4_12 = 1'b1;
      end else begin
        debug_4_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_12 = 1'b0;
    if(when_ArraySlice_l158_101) begin
      if(when_ArraySlice_l159_101) begin
        debug_5_12 = 1'b1;
      end else begin
        debug_5_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_101) begin
        debug_5_12 = 1'b1;
      end else begin
        debug_5_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_12 = 1'b0;
    if(when_ArraySlice_l158_102) begin
      if(when_ArraySlice_l159_102) begin
        debug_6_12 = 1'b1;
      end else begin
        debug_6_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_102) begin
        debug_6_12 = 1'b1;
      end else begin
        debug_6_12 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_12 = 1'b0;
    if(when_ArraySlice_l158_103) begin
      if(when_ArraySlice_l159_103) begin
        debug_7_12 = 1'b1;
      end else begin
        debug_7_12 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_103) begin
        debug_7_12 = 1'b1;
      end else begin
        debug_7_12 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_96 = (_zz_when_ArraySlice_l158_96 <= _zz_when_ArraySlice_l158_96_3);
  assign when_ArraySlice_l159_96 = (_zz_when_ArraySlice_l159_96 <= _zz_when_ArraySlice_l159_96_1);
  assign _zz_realValue_0_96 = (_zz__zz_realValue_0_96 % _zz__zz_realValue_0_96_1);
  assign when_ArraySlice_l110_96 = (_zz_realValue_0_96 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_96) begin
      realValue_0_96 = (_zz_realValue_0_96_1 - _zz_realValue_0_96);
    end else begin
      realValue_0_96 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_96 = (_zz_when_ArraySlice_l166_96 <= _zz_when_ArraySlice_l166_96_1);
  assign when_ArraySlice_l158_97 = (_zz_when_ArraySlice_l158_97 <= _zz_when_ArraySlice_l158_97_3);
  assign when_ArraySlice_l159_97 = (_zz_when_ArraySlice_l159_97 <= _zz_when_ArraySlice_l159_97_2);
  assign _zz_realValue_0_97 = (_zz__zz_realValue_0_97 % _zz__zz_realValue_0_97_1);
  assign when_ArraySlice_l110_97 = (_zz_realValue_0_97 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_97) begin
      realValue_0_97 = (_zz_realValue_0_97_1 - _zz_realValue_0_97);
    end else begin
      realValue_0_97 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_97 = (_zz_when_ArraySlice_l166_97 <= _zz_when_ArraySlice_l166_97_2);
  assign when_ArraySlice_l158_98 = (_zz_when_ArraySlice_l158_98 <= _zz_when_ArraySlice_l158_98_3);
  assign when_ArraySlice_l159_98 = (_zz_when_ArraySlice_l159_98 <= _zz_when_ArraySlice_l159_98_2);
  assign _zz_realValue_0_98 = (_zz__zz_realValue_0_98 % _zz__zz_realValue_0_98_1);
  assign when_ArraySlice_l110_98 = (_zz_realValue_0_98 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_98) begin
      realValue_0_98 = (_zz_realValue_0_98_1 - _zz_realValue_0_98);
    end else begin
      realValue_0_98 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_98 = (_zz_when_ArraySlice_l166_98 <= _zz_when_ArraySlice_l166_98_2);
  assign when_ArraySlice_l158_99 = (_zz_when_ArraySlice_l158_99 <= _zz_when_ArraySlice_l158_99_3);
  assign when_ArraySlice_l159_99 = (_zz_when_ArraySlice_l159_99 <= _zz_when_ArraySlice_l159_99_2);
  assign _zz_realValue_0_99 = (_zz__zz_realValue_0_99 % _zz__zz_realValue_0_99_1);
  assign when_ArraySlice_l110_99 = (_zz_realValue_0_99 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_99) begin
      realValue_0_99 = (_zz_realValue_0_99_1 - _zz_realValue_0_99);
    end else begin
      realValue_0_99 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_99 = (_zz_when_ArraySlice_l166_99 <= _zz_when_ArraySlice_l166_99_2);
  assign when_ArraySlice_l158_100 = (_zz_when_ArraySlice_l158_100 <= _zz_when_ArraySlice_l158_100_3);
  assign when_ArraySlice_l159_100 = (_zz_when_ArraySlice_l159_100 <= _zz_when_ArraySlice_l159_100_2);
  assign _zz_realValue_0_100 = (_zz__zz_realValue_0_100 % _zz__zz_realValue_0_100_1);
  assign when_ArraySlice_l110_100 = (_zz_realValue_0_100 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_100) begin
      realValue_0_100 = (_zz_realValue_0_100_1 - _zz_realValue_0_100);
    end else begin
      realValue_0_100 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_100 = (_zz_when_ArraySlice_l166_100 <= _zz_when_ArraySlice_l166_100_2);
  assign when_ArraySlice_l158_101 = (_zz_when_ArraySlice_l158_101 <= _zz_when_ArraySlice_l158_101_3);
  assign when_ArraySlice_l159_101 = (_zz_when_ArraySlice_l159_101 <= _zz_when_ArraySlice_l159_101_2);
  assign _zz_realValue_0_101 = (_zz__zz_realValue_0_101 % _zz__zz_realValue_0_101_1);
  assign when_ArraySlice_l110_101 = (_zz_realValue_0_101 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_101) begin
      realValue_0_101 = (_zz_realValue_0_101_1 - _zz_realValue_0_101);
    end else begin
      realValue_0_101 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_101 = (_zz_when_ArraySlice_l166_101 <= _zz_when_ArraySlice_l166_101_2);
  assign when_ArraySlice_l158_102 = (_zz_when_ArraySlice_l158_102 <= _zz_when_ArraySlice_l158_102_3);
  assign when_ArraySlice_l159_102 = (_zz_when_ArraySlice_l159_102 <= _zz_when_ArraySlice_l159_102_2);
  assign _zz_realValue_0_102 = (_zz__zz_realValue_0_102 % _zz__zz_realValue_0_102_1);
  assign when_ArraySlice_l110_102 = (_zz_realValue_0_102 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_102) begin
      realValue_0_102 = (_zz_realValue_0_102_1 - _zz_realValue_0_102);
    end else begin
      realValue_0_102 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_102 = (_zz_when_ArraySlice_l166_102 <= _zz_when_ArraySlice_l166_102_2);
  assign when_ArraySlice_l158_103 = (_zz_when_ArraySlice_l158_103 <= _zz_when_ArraySlice_l158_103_3);
  assign when_ArraySlice_l159_103 = (_zz_when_ArraySlice_l159_103 <= _zz_when_ArraySlice_l159_103_2);
  assign _zz_realValue_0_103 = (_zz__zz_realValue_0_103 % _zz__zz_realValue_0_103_1);
  assign when_ArraySlice_l110_103 = (_zz_realValue_0_103 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_103) begin
      realValue_0_103 = (_zz_realValue_0_103_1 - _zz_realValue_0_103);
    end else begin
      realValue_0_103 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_103 = (_zz_when_ArraySlice_l166_103 <= _zz_when_ArraySlice_l166_103_2);
  assign when_ArraySlice_l457_3 = (! ((((((_zz_when_ArraySlice_l457_3_1 && _zz_when_ArraySlice_l457_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l457_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_3_4 && _zz_when_ArraySlice_l457_3_5) && (debug_4_12 == _zz_when_ArraySlice_l457_3_6)) && (debug_5_12 == 1'b1)) && (debug_6_12 == 1'b1)) && (debug_7_12 == 1'b1))));
  assign outputStreamArrayData_3_fire_5 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l461_3 = ((_zz_when_ArraySlice_l461_3 == 13'h0) && outputStreamArrayData_3_fire_5);
  assign when_ArraySlice_l447_3 = (allowPadding_3 && (_zz_when_ArraySlice_l447_3_1 <= _zz_when_ArraySlice_l447_3_2));
  assign outputStreamArrayData_3_fire_6 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l468_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l468_3);
  assign when_ArraySlice_l376_4 = (_zz_when_ArraySlice_l376_4 < _zz_when_ArraySlice_l376_4_3);
  assign when_ArraySlice_l377_4 = ((! holdReadOp_4) && (_zz_when_ArraySlice_l377_4_1 != 7'h0));
  assign _zz_outputStreamArrayData_4_valid = (selectReadFifo_4 + _zz__zz_outputStreamArrayData_4_valid);
  assign _zz_7 = ({127'd0,1'b1} <<< _zz__zz_7);
  assign _zz_io_pop_ready_4 = outputStreamArrayData_4_ready;
  assign when_ArraySlice_l382_4 = (! holdReadOp_4);
  assign outputStreamArrayData_4_fire = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l383_4 = ((7'h01 < _zz_when_ArraySlice_l383_4_1) && outputStreamArrayData_4_fire);
  assign when_ArraySlice_l384_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l384_4);
  assign when_ArraySlice_l387_4 = (_zz_when_ArraySlice_l387_4 == 13'h0);
  assign outputStreamArrayData_4_fire_1 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l392_4 = ((_zz_when_ArraySlice_l392_4_1 == 7'h01) && outputStreamArrayData_4_fire_1);
  assign when_ArraySlice_l393_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l393_4);
  assign _zz_realValue1_0_12 = (_zz__zz_realValue1_0_12 % _zz__zz_realValue1_0_12_1);
  assign when_ArraySlice_l95_12 = (_zz_realValue1_0_12 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_12) begin
      realValue1_0_12 = (_zz_realValue1_0_12_1 - _zz_realValue1_0_12);
    end else begin
      realValue1_0_12 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_4 = (_zz_when_ArraySlice_l395_4 < _zz_when_ArraySlice_l395_4_2);
  always @(*) begin
    debug_0_13 = 1'b0;
    if(when_ArraySlice_l158_104) begin
      if(when_ArraySlice_l159_104) begin
        debug_0_13 = 1'b1;
      end else begin
        debug_0_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_104) begin
        debug_0_13 = 1'b1;
      end else begin
        debug_0_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_13 = 1'b0;
    if(when_ArraySlice_l158_105) begin
      if(when_ArraySlice_l159_105) begin
        debug_1_13 = 1'b1;
      end else begin
        debug_1_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_105) begin
        debug_1_13 = 1'b1;
      end else begin
        debug_1_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_13 = 1'b0;
    if(when_ArraySlice_l158_106) begin
      if(when_ArraySlice_l159_106) begin
        debug_2_13 = 1'b1;
      end else begin
        debug_2_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_106) begin
        debug_2_13 = 1'b1;
      end else begin
        debug_2_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_13 = 1'b0;
    if(when_ArraySlice_l158_107) begin
      if(when_ArraySlice_l159_107) begin
        debug_3_13 = 1'b1;
      end else begin
        debug_3_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_107) begin
        debug_3_13 = 1'b1;
      end else begin
        debug_3_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_13 = 1'b0;
    if(when_ArraySlice_l158_108) begin
      if(when_ArraySlice_l159_108) begin
        debug_4_13 = 1'b1;
      end else begin
        debug_4_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_108) begin
        debug_4_13 = 1'b1;
      end else begin
        debug_4_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_13 = 1'b0;
    if(when_ArraySlice_l158_109) begin
      if(when_ArraySlice_l159_109) begin
        debug_5_13 = 1'b1;
      end else begin
        debug_5_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_109) begin
        debug_5_13 = 1'b1;
      end else begin
        debug_5_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_13 = 1'b0;
    if(when_ArraySlice_l158_110) begin
      if(when_ArraySlice_l159_110) begin
        debug_6_13 = 1'b1;
      end else begin
        debug_6_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_110) begin
        debug_6_13 = 1'b1;
      end else begin
        debug_6_13 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_13 = 1'b0;
    if(when_ArraySlice_l158_111) begin
      if(when_ArraySlice_l159_111) begin
        debug_7_13 = 1'b1;
      end else begin
        debug_7_13 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_111) begin
        debug_7_13 = 1'b1;
      end else begin
        debug_7_13 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_104 = (_zz_when_ArraySlice_l158_104 <= _zz_when_ArraySlice_l158_104_3);
  assign when_ArraySlice_l159_104 = (_zz_when_ArraySlice_l159_104 <= _zz_when_ArraySlice_l159_104_1);
  assign _zz_realValue_0_104 = (_zz__zz_realValue_0_104 % _zz__zz_realValue_0_104_1);
  assign when_ArraySlice_l110_104 = (_zz_realValue_0_104 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_104) begin
      realValue_0_104 = (_zz_realValue_0_104_1 - _zz_realValue_0_104);
    end else begin
      realValue_0_104 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_104 = (_zz_when_ArraySlice_l166_104 <= _zz_when_ArraySlice_l166_104_1);
  assign when_ArraySlice_l158_105 = (_zz_when_ArraySlice_l158_105 <= _zz_when_ArraySlice_l158_105_3);
  assign when_ArraySlice_l159_105 = (_zz_when_ArraySlice_l159_105 <= _zz_when_ArraySlice_l159_105_2);
  assign _zz_realValue_0_105 = (_zz__zz_realValue_0_105 % _zz__zz_realValue_0_105_1);
  assign when_ArraySlice_l110_105 = (_zz_realValue_0_105 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_105) begin
      realValue_0_105 = (_zz_realValue_0_105_1 - _zz_realValue_0_105);
    end else begin
      realValue_0_105 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_105 = (_zz_when_ArraySlice_l166_105 <= _zz_when_ArraySlice_l166_105_2);
  assign when_ArraySlice_l158_106 = (_zz_when_ArraySlice_l158_106 <= _zz_when_ArraySlice_l158_106_3);
  assign when_ArraySlice_l159_106 = (_zz_when_ArraySlice_l159_106 <= _zz_when_ArraySlice_l159_106_2);
  assign _zz_realValue_0_106 = (_zz__zz_realValue_0_106 % _zz__zz_realValue_0_106_1);
  assign when_ArraySlice_l110_106 = (_zz_realValue_0_106 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_106) begin
      realValue_0_106 = (_zz_realValue_0_106_1 - _zz_realValue_0_106);
    end else begin
      realValue_0_106 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_106 = (_zz_when_ArraySlice_l166_106 <= _zz_when_ArraySlice_l166_106_2);
  assign when_ArraySlice_l158_107 = (_zz_when_ArraySlice_l158_107 <= _zz_when_ArraySlice_l158_107_3);
  assign when_ArraySlice_l159_107 = (_zz_when_ArraySlice_l159_107 <= _zz_when_ArraySlice_l159_107_2);
  assign _zz_realValue_0_107 = (_zz__zz_realValue_0_107 % _zz__zz_realValue_0_107_1);
  assign when_ArraySlice_l110_107 = (_zz_realValue_0_107 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_107) begin
      realValue_0_107 = (_zz_realValue_0_107_1 - _zz_realValue_0_107);
    end else begin
      realValue_0_107 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_107 = (_zz_when_ArraySlice_l166_107 <= _zz_when_ArraySlice_l166_107_2);
  assign when_ArraySlice_l158_108 = (_zz_when_ArraySlice_l158_108 <= _zz_when_ArraySlice_l158_108_3);
  assign when_ArraySlice_l159_108 = (_zz_when_ArraySlice_l159_108 <= _zz_when_ArraySlice_l159_108_2);
  assign _zz_realValue_0_108 = (_zz__zz_realValue_0_108 % _zz__zz_realValue_0_108_1);
  assign when_ArraySlice_l110_108 = (_zz_realValue_0_108 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_108) begin
      realValue_0_108 = (_zz_realValue_0_108_1 - _zz_realValue_0_108);
    end else begin
      realValue_0_108 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_108 = (_zz_when_ArraySlice_l166_108 <= _zz_when_ArraySlice_l166_108_2);
  assign when_ArraySlice_l158_109 = (_zz_when_ArraySlice_l158_109 <= _zz_when_ArraySlice_l158_109_3);
  assign when_ArraySlice_l159_109 = (_zz_when_ArraySlice_l159_109 <= _zz_when_ArraySlice_l159_109_2);
  assign _zz_realValue_0_109 = (_zz__zz_realValue_0_109 % _zz__zz_realValue_0_109_1);
  assign when_ArraySlice_l110_109 = (_zz_realValue_0_109 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_109) begin
      realValue_0_109 = (_zz_realValue_0_109_1 - _zz_realValue_0_109);
    end else begin
      realValue_0_109 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_109 = (_zz_when_ArraySlice_l166_109 <= _zz_when_ArraySlice_l166_109_2);
  assign when_ArraySlice_l158_110 = (_zz_when_ArraySlice_l158_110 <= _zz_when_ArraySlice_l158_110_3);
  assign when_ArraySlice_l159_110 = (_zz_when_ArraySlice_l159_110 <= _zz_when_ArraySlice_l159_110_2);
  assign _zz_realValue_0_110 = (_zz__zz_realValue_0_110 % _zz__zz_realValue_0_110_1);
  assign when_ArraySlice_l110_110 = (_zz_realValue_0_110 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_110) begin
      realValue_0_110 = (_zz_realValue_0_110_1 - _zz_realValue_0_110);
    end else begin
      realValue_0_110 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_110 = (_zz_when_ArraySlice_l166_110 <= _zz_when_ArraySlice_l166_110_2);
  assign when_ArraySlice_l158_111 = (_zz_when_ArraySlice_l158_111 <= _zz_when_ArraySlice_l158_111_3);
  assign when_ArraySlice_l159_111 = (_zz_when_ArraySlice_l159_111 <= _zz_when_ArraySlice_l159_111_2);
  assign _zz_realValue_0_111 = (_zz__zz_realValue_0_111 % _zz__zz_realValue_0_111_1);
  assign when_ArraySlice_l110_111 = (_zz_realValue_0_111 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_111) begin
      realValue_0_111 = (_zz_realValue_0_111_1 - _zz_realValue_0_111);
    end else begin
      realValue_0_111 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_111 = (_zz_when_ArraySlice_l166_111 <= _zz_when_ArraySlice_l166_111_2);
  assign when_ArraySlice_l400_4 = (! ((((((_zz_when_ArraySlice_l400_4_1 && _zz_when_ArraySlice_l400_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_4_4 && _zz_when_ArraySlice_l400_4_5) && (debug_4_13 == _zz_when_ArraySlice_l400_4_6)) && (debug_5_13 == 1'b1)) && (debug_6_13 == 1'b1)) && (debug_7_13 == 1'b1))));
  assign when_ArraySlice_l403_4 = (_zz_when_ArraySlice_l403_4_1 <= _zz_when_ArraySlice_l403_4_2);
  assign when_ArraySlice_l406_4 = (_zz_when_ArraySlice_l406_4_1 <= _zz_when_ArraySlice_l406_4_2);
  assign when_ArraySlice_l413_4 = (_zz_when_ArraySlice_l413_4 == 13'h0);
  assign when_ArraySlice_l417_4 = (_zz_when_ArraySlice_l417_4_1 == 7'h0);
  assign outputStreamArrayData_4_fire_2 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l418_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l418_4_1) && outputStreamArrayData_4_fire_2);
  assign _zz_realValue1_0_13 = (_zz__zz_realValue1_0_13 % _zz__zz_realValue1_0_13_1);
  assign when_ArraySlice_l95_13 = (_zz_realValue1_0_13 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_13) begin
      realValue1_0_13 = (_zz_realValue1_0_13_1 - _zz_realValue1_0_13);
    end else begin
      realValue1_0_13 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_4 = (_zz_when_ArraySlice_l420_4 < _zz_when_ArraySlice_l420_4_2);
  always @(*) begin
    debug_0_14 = 1'b0;
    if(when_ArraySlice_l158_112) begin
      if(when_ArraySlice_l159_112) begin
        debug_0_14 = 1'b1;
      end else begin
        debug_0_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_112) begin
        debug_0_14 = 1'b1;
      end else begin
        debug_0_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_14 = 1'b0;
    if(when_ArraySlice_l158_113) begin
      if(when_ArraySlice_l159_113) begin
        debug_1_14 = 1'b1;
      end else begin
        debug_1_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_113) begin
        debug_1_14 = 1'b1;
      end else begin
        debug_1_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_14 = 1'b0;
    if(when_ArraySlice_l158_114) begin
      if(when_ArraySlice_l159_114) begin
        debug_2_14 = 1'b1;
      end else begin
        debug_2_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_114) begin
        debug_2_14 = 1'b1;
      end else begin
        debug_2_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_14 = 1'b0;
    if(when_ArraySlice_l158_115) begin
      if(when_ArraySlice_l159_115) begin
        debug_3_14 = 1'b1;
      end else begin
        debug_3_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_115) begin
        debug_3_14 = 1'b1;
      end else begin
        debug_3_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_14 = 1'b0;
    if(when_ArraySlice_l158_116) begin
      if(when_ArraySlice_l159_116) begin
        debug_4_14 = 1'b1;
      end else begin
        debug_4_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_116) begin
        debug_4_14 = 1'b1;
      end else begin
        debug_4_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_14 = 1'b0;
    if(when_ArraySlice_l158_117) begin
      if(when_ArraySlice_l159_117) begin
        debug_5_14 = 1'b1;
      end else begin
        debug_5_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_117) begin
        debug_5_14 = 1'b1;
      end else begin
        debug_5_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_14 = 1'b0;
    if(when_ArraySlice_l158_118) begin
      if(when_ArraySlice_l159_118) begin
        debug_6_14 = 1'b1;
      end else begin
        debug_6_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_118) begin
        debug_6_14 = 1'b1;
      end else begin
        debug_6_14 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_14 = 1'b0;
    if(when_ArraySlice_l158_119) begin
      if(when_ArraySlice_l159_119) begin
        debug_7_14 = 1'b1;
      end else begin
        debug_7_14 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_119) begin
        debug_7_14 = 1'b1;
      end else begin
        debug_7_14 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_112 = (_zz_when_ArraySlice_l158_112 <= _zz_when_ArraySlice_l158_112_3);
  assign when_ArraySlice_l159_112 = (_zz_when_ArraySlice_l159_112 <= _zz_when_ArraySlice_l159_112_1);
  assign _zz_realValue_0_112 = (_zz__zz_realValue_0_112 % _zz__zz_realValue_0_112_1);
  assign when_ArraySlice_l110_112 = (_zz_realValue_0_112 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_112) begin
      realValue_0_112 = (_zz_realValue_0_112_1 - _zz_realValue_0_112);
    end else begin
      realValue_0_112 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_112 = (_zz_when_ArraySlice_l166_112 <= _zz_when_ArraySlice_l166_112_1);
  assign when_ArraySlice_l158_113 = (_zz_when_ArraySlice_l158_113 <= _zz_when_ArraySlice_l158_113_3);
  assign when_ArraySlice_l159_113 = (_zz_when_ArraySlice_l159_113 <= _zz_when_ArraySlice_l159_113_2);
  assign _zz_realValue_0_113 = (_zz__zz_realValue_0_113 % _zz__zz_realValue_0_113_1);
  assign when_ArraySlice_l110_113 = (_zz_realValue_0_113 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_113) begin
      realValue_0_113 = (_zz_realValue_0_113_1 - _zz_realValue_0_113);
    end else begin
      realValue_0_113 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_113 = (_zz_when_ArraySlice_l166_113 <= _zz_when_ArraySlice_l166_113_2);
  assign when_ArraySlice_l158_114 = (_zz_when_ArraySlice_l158_114 <= _zz_when_ArraySlice_l158_114_3);
  assign when_ArraySlice_l159_114 = (_zz_when_ArraySlice_l159_114 <= _zz_when_ArraySlice_l159_114_2);
  assign _zz_realValue_0_114 = (_zz__zz_realValue_0_114 % _zz__zz_realValue_0_114_1);
  assign when_ArraySlice_l110_114 = (_zz_realValue_0_114 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_114) begin
      realValue_0_114 = (_zz_realValue_0_114_1 - _zz_realValue_0_114);
    end else begin
      realValue_0_114 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_114 = (_zz_when_ArraySlice_l166_114 <= _zz_when_ArraySlice_l166_114_2);
  assign when_ArraySlice_l158_115 = (_zz_when_ArraySlice_l158_115 <= _zz_when_ArraySlice_l158_115_3);
  assign when_ArraySlice_l159_115 = (_zz_when_ArraySlice_l159_115 <= _zz_when_ArraySlice_l159_115_2);
  assign _zz_realValue_0_115 = (_zz__zz_realValue_0_115 % _zz__zz_realValue_0_115_1);
  assign when_ArraySlice_l110_115 = (_zz_realValue_0_115 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_115) begin
      realValue_0_115 = (_zz_realValue_0_115_1 - _zz_realValue_0_115);
    end else begin
      realValue_0_115 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_115 = (_zz_when_ArraySlice_l166_115 <= _zz_when_ArraySlice_l166_115_2);
  assign when_ArraySlice_l158_116 = (_zz_when_ArraySlice_l158_116 <= _zz_when_ArraySlice_l158_116_3);
  assign when_ArraySlice_l159_116 = (_zz_when_ArraySlice_l159_116 <= _zz_when_ArraySlice_l159_116_2);
  assign _zz_realValue_0_116 = (_zz__zz_realValue_0_116 % _zz__zz_realValue_0_116_1);
  assign when_ArraySlice_l110_116 = (_zz_realValue_0_116 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_116) begin
      realValue_0_116 = (_zz_realValue_0_116_1 - _zz_realValue_0_116);
    end else begin
      realValue_0_116 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_116 = (_zz_when_ArraySlice_l166_116 <= _zz_when_ArraySlice_l166_116_2);
  assign when_ArraySlice_l158_117 = (_zz_when_ArraySlice_l158_117 <= _zz_when_ArraySlice_l158_117_3);
  assign when_ArraySlice_l159_117 = (_zz_when_ArraySlice_l159_117 <= _zz_when_ArraySlice_l159_117_2);
  assign _zz_realValue_0_117 = (_zz__zz_realValue_0_117 % _zz__zz_realValue_0_117_1);
  assign when_ArraySlice_l110_117 = (_zz_realValue_0_117 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_117) begin
      realValue_0_117 = (_zz_realValue_0_117_1 - _zz_realValue_0_117);
    end else begin
      realValue_0_117 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_117 = (_zz_when_ArraySlice_l166_117 <= _zz_when_ArraySlice_l166_117_2);
  assign when_ArraySlice_l158_118 = (_zz_when_ArraySlice_l158_118 <= _zz_when_ArraySlice_l158_118_3);
  assign when_ArraySlice_l159_118 = (_zz_when_ArraySlice_l159_118 <= _zz_when_ArraySlice_l159_118_2);
  assign _zz_realValue_0_118 = (_zz__zz_realValue_0_118 % _zz__zz_realValue_0_118_1);
  assign when_ArraySlice_l110_118 = (_zz_realValue_0_118 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_118) begin
      realValue_0_118 = (_zz_realValue_0_118_1 - _zz_realValue_0_118);
    end else begin
      realValue_0_118 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_118 = (_zz_when_ArraySlice_l166_118 <= _zz_when_ArraySlice_l166_118_2);
  assign when_ArraySlice_l158_119 = (_zz_when_ArraySlice_l158_119 <= _zz_when_ArraySlice_l158_119_3);
  assign when_ArraySlice_l159_119 = (_zz_when_ArraySlice_l159_119 <= _zz_when_ArraySlice_l159_119_2);
  assign _zz_realValue_0_119 = (_zz__zz_realValue_0_119 % _zz__zz_realValue_0_119_1);
  assign when_ArraySlice_l110_119 = (_zz_realValue_0_119 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_119) begin
      realValue_0_119 = (_zz_realValue_0_119_1 - _zz_realValue_0_119);
    end else begin
      realValue_0_119 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_119 = (_zz_when_ArraySlice_l166_119 <= _zz_when_ArraySlice_l166_119_2);
  assign when_ArraySlice_l425_4 = (! ((((((_zz_when_ArraySlice_l425_4_1 && _zz_when_ArraySlice_l425_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l425_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_4_4 && _zz_when_ArraySlice_l425_4_5) && (debug_4_14 == _zz_when_ArraySlice_l425_4_6)) && (debug_5_14 == 1'b1)) && (debug_6_14 == 1'b1)) && (debug_7_14 == 1'b1))));
  assign when_ArraySlice_l428_4 = (_zz_when_ArraySlice_l428_4_1 <= _zz_when_ArraySlice_l428_4_2);
  assign when_ArraySlice_l431_4 = (_zz_when_ArraySlice_l431_4_1 <= _zz_when_ArraySlice_l431_4_2);
  assign outputStreamArrayData_4_fire_3 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l438_4 = ((_zz_when_ArraySlice_l438_4 == 13'h0) && outputStreamArrayData_4_fire_3);
  assign outputStreamArrayData_4_fire_4 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l449_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l449_4) && outputStreamArrayData_4_fire_4);
  assign _zz_realValue1_0_14 = (_zz__zz_realValue1_0_14 % _zz__zz_realValue1_0_14_1);
  assign when_ArraySlice_l95_14 = (_zz_realValue1_0_14 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_14) begin
      realValue1_0_14 = (_zz_realValue1_0_14_1 - _zz_realValue1_0_14);
    end else begin
      realValue1_0_14 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_4 = (_zz_when_ArraySlice_l450_4 < _zz_when_ArraySlice_l450_4_2);
  always @(*) begin
    debug_0_15 = 1'b0;
    if(when_ArraySlice_l158_120) begin
      if(when_ArraySlice_l159_120) begin
        debug_0_15 = 1'b1;
      end else begin
        debug_0_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_120) begin
        debug_0_15 = 1'b1;
      end else begin
        debug_0_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_15 = 1'b0;
    if(when_ArraySlice_l158_121) begin
      if(when_ArraySlice_l159_121) begin
        debug_1_15 = 1'b1;
      end else begin
        debug_1_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_121) begin
        debug_1_15 = 1'b1;
      end else begin
        debug_1_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_15 = 1'b0;
    if(when_ArraySlice_l158_122) begin
      if(when_ArraySlice_l159_122) begin
        debug_2_15 = 1'b1;
      end else begin
        debug_2_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_122) begin
        debug_2_15 = 1'b1;
      end else begin
        debug_2_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_15 = 1'b0;
    if(when_ArraySlice_l158_123) begin
      if(when_ArraySlice_l159_123) begin
        debug_3_15 = 1'b1;
      end else begin
        debug_3_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_123) begin
        debug_3_15 = 1'b1;
      end else begin
        debug_3_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_15 = 1'b0;
    if(when_ArraySlice_l158_124) begin
      if(when_ArraySlice_l159_124) begin
        debug_4_15 = 1'b1;
      end else begin
        debug_4_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_124) begin
        debug_4_15 = 1'b1;
      end else begin
        debug_4_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_15 = 1'b0;
    if(when_ArraySlice_l158_125) begin
      if(when_ArraySlice_l159_125) begin
        debug_5_15 = 1'b1;
      end else begin
        debug_5_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_125) begin
        debug_5_15 = 1'b1;
      end else begin
        debug_5_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_15 = 1'b0;
    if(when_ArraySlice_l158_126) begin
      if(when_ArraySlice_l159_126) begin
        debug_6_15 = 1'b1;
      end else begin
        debug_6_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_126) begin
        debug_6_15 = 1'b1;
      end else begin
        debug_6_15 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_15 = 1'b0;
    if(when_ArraySlice_l158_127) begin
      if(when_ArraySlice_l159_127) begin
        debug_7_15 = 1'b1;
      end else begin
        debug_7_15 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_127) begin
        debug_7_15 = 1'b1;
      end else begin
        debug_7_15 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_120 = (_zz_when_ArraySlice_l158_120 <= _zz_when_ArraySlice_l158_120_3);
  assign when_ArraySlice_l159_120 = (_zz_when_ArraySlice_l159_120 <= _zz_when_ArraySlice_l159_120_1);
  assign _zz_realValue_0_120 = (_zz__zz_realValue_0_120 % _zz__zz_realValue_0_120_1);
  assign when_ArraySlice_l110_120 = (_zz_realValue_0_120 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_120) begin
      realValue_0_120 = (_zz_realValue_0_120_1 - _zz_realValue_0_120);
    end else begin
      realValue_0_120 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_120 = (_zz_when_ArraySlice_l166_120 <= _zz_when_ArraySlice_l166_120_1);
  assign when_ArraySlice_l158_121 = (_zz_when_ArraySlice_l158_121 <= _zz_when_ArraySlice_l158_121_3);
  assign when_ArraySlice_l159_121 = (_zz_when_ArraySlice_l159_121 <= _zz_when_ArraySlice_l159_121_2);
  assign _zz_realValue_0_121 = (_zz__zz_realValue_0_121 % _zz__zz_realValue_0_121_1);
  assign when_ArraySlice_l110_121 = (_zz_realValue_0_121 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_121) begin
      realValue_0_121 = (_zz_realValue_0_121_1 - _zz_realValue_0_121);
    end else begin
      realValue_0_121 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_121 = (_zz_when_ArraySlice_l166_121 <= _zz_when_ArraySlice_l166_121_2);
  assign when_ArraySlice_l158_122 = (_zz_when_ArraySlice_l158_122 <= _zz_when_ArraySlice_l158_122_3);
  assign when_ArraySlice_l159_122 = (_zz_when_ArraySlice_l159_122 <= _zz_when_ArraySlice_l159_122_2);
  assign _zz_realValue_0_122 = (_zz__zz_realValue_0_122 % _zz__zz_realValue_0_122_1);
  assign when_ArraySlice_l110_122 = (_zz_realValue_0_122 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_122) begin
      realValue_0_122 = (_zz_realValue_0_122_1 - _zz_realValue_0_122);
    end else begin
      realValue_0_122 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_122 = (_zz_when_ArraySlice_l166_122 <= _zz_when_ArraySlice_l166_122_2);
  assign when_ArraySlice_l158_123 = (_zz_when_ArraySlice_l158_123 <= _zz_when_ArraySlice_l158_123_3);
  assign when_ArraySlice_l159_123 = (_zz_when_ArraySlice_l159_123 <= _zz_when_ArraySlice_l159_123_2);
  assign _zz_realValue_0_123 = (_zz__zz_realValue_0_123 % _zz__zz_realValue_0_123_1);
  assign when_ArraySlice_l110_123 = (_zz_realValue_0_123 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_123) begin
      realValue_0_123 = (_zz_realValue_0_123_1 - _zz_realValue_0_123);
    end else begin
      realValue_0_123 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_123 = (_zz_when_ArraySlice_l166_123 <= _zz_when_ArraySlice_l166_123_2);
  assign when_ArraySlice_l158_124 = (_zz_when_ArraySlice_l158_124 <= _zz_when_ArraySlice_l158_124_3);
  assign when_ArraySlice_l159_124 = (_zz_when_ArraySlice_l159_124 <= _zz_when_ArraySlice_l159_124_2);
  assign _zz_realValue_0_124 = (_zz__zz_realValue_0_124 % _zz__zz_realValue_0_124_1);
  assign when_ArraySlice_l110_124 = (_zz_realValue_0_124 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_124) begin
      realValue_0_124 = (_zz_realValue_0_124_1 - _zz_realValue_0_124);
    end else begin
      realValue_0_124 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_124 = (_zz_when_ArraySlice_l166_124 <= _zz_when_ArraySlice_l166_124_2);
  assign when_ArraySlice_l158_125 = (_zz_when_ArraySlice_l158_125 <= _zz_when_ArraySlice_l158_125_3);
  assign when_ArraySlice_l159_125 = (_zz_when_ArraySlice_l159_125 <= _zz_when_ArraySlice_l159_125_2);
  assign _zz_realValue_0_125 = (_zz__zz_realValue_0_125 % _zz__zz_realValue_0_125_1);
  assign when_ArraySlice_l110_125 = (_zz_realValue_0_125 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_125) begin
      realValue_0_125 = (_zz_realValue_0_125_1 - _zz_realValue_0_125);
    end else begin
      realValue_0_125 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_125 = (_zz_when_ArraySlice_l166_125 <= _zz_when_ArraySlice_l166_125_2);
  assign when_ArraySlice_l158_126 = (_zz_when_ArraySlice_l158_126 <= _zz_when_ArraySlice_l158_126_3);
  assign when_ArraySlice_l159_126 = (_zz_when_ArraySlice_l159_126 <= _zz_when_ArraySlice_l159_126_2);
  assign _zz_realValue_0_126 = (_zz__zz_realValue_0_126 % _zz__zz_realValue_0_126_1);
  assign when_ArraySlice_l110_126 = (_zz_realValue_0_126 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_126) begin
      realValue_0_126 = (_zz_realValue_0_126_1 - _zz_realValue_0_126);
    end else begin
      realValue_0_126 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_126 = (_zz_when_ArraySlice_l166_126 <= _zz_when_ArraySlice_l166_126_2);
  assign when_ArraySlice_l158_127 = (_zz_when_ArraySlice_l158_127 <= _zz_when_ArraySlice_l158_127_3);
  assign when_ArraySlice_l159_127 = (_zz_when_ArraySlice_l159_127 <= _zz_when_ArraySlice_l159_127_2);
  assign _zz_realValue_0_127 = (_zz__zz_realValue_0_127 % _zz__zz_realValue_0_127_1);
  assign when_ArraySlice_l110_127 = (_zz_realValue_0_127 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_127) begin
      realValue_0_127 = (_zz_realValue_0_127_1 - _zz_realValue_0_127);
    end else begin
      realValue_0_127 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_127 = (_zz_when_ArraySlice_l166_127 <= _zz_when_ArraySlice_l166_127_2);
  assign when_ArraySlice_l457_4 = (! ((((((_zz_when_ArraySlice_l457_4_1 && _zz_when_ArraySlice_l457_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l457_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_4_4 && _zz_when_ArraySlice_l457_4_5) && (debug_4_15 == _zz_when_ArraySlice_l457_4_6)) && (debug_5_15 == 1'b1)) && (debug_6_15 == 1'b1)) && (debug_7_15 == 1'b1))));
  assign outputStreamArrayData_4_fire_5 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l461_4 = ((_zz_when_ArraySlice_l461_4 == 13'h0) && outputStreamArrayData_4_fire_5);
  assign when_ArraySlice_l447_4 = (allowPadding_4 && (_zz_when_ArraySlice_l447_4 <= _zz_when_ArraySlice_l447_4_1));
  assign outputStreamArrayData_4_fire_6 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l468_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l468_4);
  assign when_ArraySlice_l376_5 = (_zz_when_ArraySlice_l376_5 < _zz_when_ArraySlice_l376_5_3);
  assign when_ArraySlice_l377_5 = ((! holdReadOp_5) && (_zz_when_ArraySlice_l377_5 != 7'h0));
  assign _zz_outputStreamArrayData_5_valid = (selectReadFifo_5 + _zz__zz_outputStreamArrayData_5_valid);
  assign _zz_8 = ({127'd0,1'b1} <<< _zz__zz_8);
  assign _zz_io_pop_ready_5 = outputStreamArrayData_5_ready;
  assign when_ArraySlice_l382_5 = (! holdReadOp_5);
  assign outputStreamArrayData_5_fire = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l383_5 = ((7'h01 < _zz_when_ArraySlice_l383_5) && outputStreamArrayData_5_fire);
  assign when_ArraySlice_l384_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l384_5);
  assign when_ArraySlice_l387_5 = (_zz_when_ArraySlice_l387_5 == 13'h0);
  assign outputStreamArrayData_5_fire_1 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l392_5 = ((_zz_when_ArraySlice_l392_5 == 7'h01) && outputStreamArrayData_5_fire_1);
  assign when_ArraySlice_l393_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l393_5);
  assign _zz_realValue1_0_15 = (_zz__zz_realValue1_0_15 % _zz__zz_realValue1_0_15_1);
  assign when_ArraySlice_l95_15 = (_zz_realValue1_0_15 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_15) begin
      realValue1_0_15 = (_zz_realValue1_0_15_1 - _zz_realValue1_0_15);
    end else begin
      realValue1_0_15 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_5 = (_zz_when_ArraySlice_l395_5 < _zz_when_ArraySlice_l395_5_2);
  always @(*) begin
    debug_0_16 = 1'b0;
    if(when_ArraySlice_l158_128) begin
      if(when_ArraySlice_l159_128) begin
        debug_0_16 = 1'b1;
      end else begin
        debug_0_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_128) begin
        debug_0_16 = 1'b1;
      end else begin
        debug_0_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_16 = 1'b0;
    if(when_ArraySlice_l158_129) begin
      if(when_ArraySlice_l159_129) begin
        debug_1_16 = 1'b1;
      end else begin
        debug_1_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_129) begin
        debug_1_16 = 1'b1;
      end else begin
        debug_1_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_16 = 1'b0;
    if(when_ArraySlice_l158_130) begin
      if(when_ArraySlice_l159_130) begin
        debug_2_16 = 1'b1;
      end else begin
        debug_2_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_130) begin
        debug_2_16 = 1'b1;
      end else begin
        debug_2_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_16 = 1'b0;
    if(when_ArraySlice_l158_131) begin
      if(when_ArraySlice_l159_131) begin
        debug_3_16 = 1'b1;
      end else begin
        debug_3_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_131) begin
        debug_3_16 = 1'b1;
      end else begin
        debug_3_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_16 = 1'b0;
    if(when_ArraySlice_l158_132) begin
      if(when_ArraySlice_l159_132) begin
        debug_4_16 = 1'b1;
      end else begin
        debug_4_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_132) begin
        debug_4_16 = 1'b1;
      end else begin
        debug_4_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_16 = 1'b0;
    if(when_ArraySlice_l158_133) begin
      if(when_ArraySlice_l159_133) begin
        debug_5_16 = 1'b1;
      end else begin
        debug_5_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_133) begin
        debug_5_16 = 1'b1;
      end else begin
        debug_5_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_16 = 1'b0;
    if(when_ArraySlice_l158_134) begin
      if(when_ArraySlice_l159_134) begin
        debug_6_16 = 1'b1;
      end else begin
        debug_6_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_134) begin
        debug_6_16 = 1'b1;
      end else begin
        debug_6_16 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_16 = 1'b0;
    if(when_ArraySlice_l158_135) begin
      if(when_ArraySlice_l159_135) begin
        debug_7_16 = 1'b1;
      end else begin
        debug_7_16 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_135) begin
        debug_7_16 = 1'b1;
      end else begin
        debug_7_16 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_128 = (_zz_when_ArraySlice_l158_128 <= _zz_when_ArraySlice_l158_128_3);
  assign when_ArraySlice_l159_128 = (_zz_when_ArraySlice_l159_128 <= _zz_when_ArraySlice_l159_128_1);
  assign _zz_realValue_0_128 = (_zz__zz_realValue_0_128 % _zz__zz_realValue_0_128_1);
  assign when_ArraySlice_l110_128 = (_zz_realValue_0_128 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_128) begin
      realValue_0_128 = (_zz_realValue_0_128_1 - _zz_realValue_0_128);
    end else begin
      realValue_0_128 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_128 = (_zz_when_ArraySlice_l166_128 <= _zz_when_ArraySlice_l166_128_1);
  assign when_ArraySlice_l158_129 = (_zz_when_ArraySlice_l158_129 <= _zz_when_ArraySlice_l158_129_3);
  assign when_ArraySlice_l159_129 = (_zz_when_ArraySlice_l159_129 <= _zz_when_ArraySlice_l159_129_2);
  assign _zz_realValue_0_129 = (_zz__zz_realValue_0_129 % _zz__zz_realValue_0_129_1);
  assign when_ArraySlice_l110_129 = (_zz_realValue_0_129 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_129) begin
      realValue_0_129 = (_zz_realValue_0_129_1 - _zz_realValue_0_129);
    end else begin
      realValue_0_129 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_129 = (_zz_when_ArraySlice_l166_129 <= _zz_when_ArraySlice_l166_129_2);
  assign when_ArraySlice_l158_130 = (_zz_when_ArraySlice_l158_130 <= _zz_when_ArraySlice_l158_130_3);
  assign when_ArraySlice_l159_130 = (_zz_when_ArraySlice_l159_130 <= _zz_when_ArraySlice_l159_130_2);
  assign _zz_realValue_0_130 = (_zz__zz_realValue_0_130 % _zz__zz_realValue_0_130_1);
  assign when_ArraySlice_l110_130 = (_zz_realValue_0_130 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_130) begin
      realValue_0_130 = (_zz_realValue_0_130_1 - _zz_realValue_0_130);
    end else begin
      realValue_0_130 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_130 = (_zz_when_ArraySlice_l166_130 <= _zz_when_ArraySlice_l166_130_2);
  assign when_ArraySlice_l158_131 = (_zz_when_ArraySlice_l158_131 <= _zz_when_ArraySlice_l158_131_3);
  assign when_ArraySlice_l159_131 = (_zz_when_ArraySlice_l159_131 <= _zz_when_ArraySlice_l159_131_2);
  assign _zz_realValue_0_131 = (_zz__zz_realValue_0_131 % _zz__zz_realValue_0_131_1);
  assign when_ArraySlice_l110_131 = (_zz_realValue_0_131 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_131) begin
      realValue_0_131 = (_zz_realValue_0_131_1 - _zz_realValue_0_131);
    end else begin
      realValue_0_131 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_131 = (_zz_when_ArraySlice_l166_131 <= _zz_when_ArraySlice_l166_131_2);
  assign when_ArraySlice_l158_132 = (_zz_when_ArraySlice_l158_132 <= _zz_when_ArraySlice_l158_132_3);
  assign when_ArraySlice_l159_132 = (_zz_when_ArraySlice_l159_132 <= _zz_when_ArraySlice_l159_132_2);
  assign _zz_realValue_0_132 = (_zz__zz_realValue_0_132 % _zz__zz_realValue_0_132_1);
  assign when_ArraySlice_l110_132 = (_zz_realValue_0_132 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_132) begin
      realValue_0_132 = (_zz_realValue_0_132_1 - _zz_realValue_0_132);
    end else begin
      realValue_0_132 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_132 = (_zz_when_ArraySlice_l166_132 <= _zz_when_ArraySlice_l166_132_2);
  assign when_ArraySlice_l158_133 = (_zz_when_ArraySlice_l158_133 <= _zz_when_ArraySlice_l158_133_3);
  assign when_ArraySlice_l159_133 = (_zz_when_ArraySlice_l159_133 <= _zz_when_ArraySlice_l159_133_2);
  assign _zz_realValue_0_133 = (_zz__zz_realValue_0_133 % _zz__zz_realValue_0_133_1);
  assign when_ArraySlice_l110_133 = (_zz_realValue_0_133 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_133) begin
      realValue_0_133 = (_zz_realValue_0_133_1 - _zz_realValue_0_133);
    end else begin
      realValue_0_133 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_133 = (_zz_when_ArraySlice_l166_133 <= _zz_when_ArraySlice_l166_133_2);
  assign when_ArraySlice_l158_134 = (_zz_when_ArraySlice_l158_134 <= _zz_when_ArraySlice_l158_134_3);
  assign when_ArraySlice_l159_134 = (_zz_when_ArraySlice_l159_134 <= _zz_when_ArraySlice_l159_134_2);
  assign _zz_realValue_0_134 = (_zz__zz_realValue_0_134 % _zz__zz_realValue_0_134_1);
  assign when_ArraySlice_l110_134 = (_zz_realValue_0_134 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_134) begin
      realValue_0_134 = (_zz_realValue_0_134_1 - _zz_realValue_0_134);
    end else begin
      realValue_0_134 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_134 = (_zz_when_ArraySlice_l166_134 <= _zz_when_ArraySlice_l166_134_2);
  assign when_ArraySlice_l158_135 = (_zz_when_ArraySlice_l158_135 <= _zz_when_ArraySlice_l158_135_3);
  assign when_ArraySlice_l159_135 = (_zz_when_ArraySlice_l159_135 <= _zz_when_ArraySlice_l159_135_2);
  assign _zz_realValue_0_135 = (_zz__zz_realValue_0_135 % _zz__zz_realValue_0_135_1);
  assign when_ArraySlice_l110_135 = (_zz_realValue_0_135 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_135) begin
      realValue_0_135 = (_zz_realValue_0_135_1 - _zz_realValue_0_135);
    end else begin
      realValue_0_135 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_135 = (_zz_when_ArraySlice_l166_135 <= _zz_when_ArraySlice_l166_135_2);
  assign when_ArraySlice_l400_5 = (! ((((((_zz_when_ArraySlice_l400_5_1 && _zz_when_ArraySlice_l400_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_5_4 && _zz_when_ArraySlice_l400_5_5) && (debug_4_16 == _zz_when_ArraySlice_l400_5_6)) && (debug_5_16 == 1'b1)) && (debug_6_16 == 1'b1)) && (debug_7_16 == 1'b1))));
  assign when_ArraySlice_l403_5 = (_zz_when_ArraySlice_l403_5_1 <= _zz_when_ArraySlice_l403_5_2);
  assign when_ArraySlice_l406_5 = (_zz_when_ArraySlice_l406_5 <= _zz_when_ArraySlice_l406_5_1);
  assign when_ArraySlice_l413_5 = (_zz_when_ArraySlice_l413_5 == 13'h0);
  assign when_ArraySlice_l417_5 = (_zz_when_ArraySlice_l417_5 == 7'h0);
  assign outputStreamArrayData_5_fire_2 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l418_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l418_5) && outputStreamArrayData_5_fire_2);
  assign _zz_realValue1_0_16 = (_zz__zz_realValue1_0_16 % _zz__zz_realValue1_0_16_1);
  assign when_ArraySlice_l95_16 = (_zz_realValue1_0_16 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_16) begin
      realValue1_0_16 = (_zz_realValue1_0_16_1 - _zz_realValue1_0_16);
    end else begin
      realValue1_0_16 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_5 = (_zz_when_ArraySlice_l420_5 < _zz_when_ArraySlice_l420_5_2);
  always @(*) begin
    debug_0_17 = 1'b0;
    if(when_ArraySlice_l158_136) begin
      if(when_ArraySlice_l159_136) begin
        debug_0_17 = 1'b1;
      end else begin
        debug_0_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_136) begin
        debug_0_17 = 1'b1;
      end else begin
        debug_0_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_17 = 1'b0;
    if(when_ArraySlice_l158_137) begin
      if(when_ArraySlice_l159_137) begin
        debug_1_17 = 1'b1;
      end else begin
        debug_1_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_137) begin
        debug_1_17 = 1'b1;
      end else begin
        debug_1_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_17 = 1'b0;
    if(when_ArraySlice_l158_138) begin
      if(when_ArraySlice_l159_138) begin
        debug_2_17 = 1'b1;
      end else begin
        debug_2_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_138) begin
        debug_2_17 = 1'b1;
      end else begin
        debug_2_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_17 = 1'b0;
    if(when_ArraySlice_l158_139) begin
      if(when_ArraySlice_l159_139) begin
        debug_3_17 = 1'b1;
      end else begin
        debug_3_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_139) begin
        debug_3_17 = 1'b1;
      end else begin
        debug_3_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_17 = 1'b0;
    if(when_ArraySlice_l158_140) begin
      if(when_ArraySlice_l159_140) begin
        debug_4_17 = 1'b1;
      end else begin
        debug_4_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_140) begin
        debug_4_17 = 1'b1;
      end else begin
        debug_4_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_17 = 1'b0;
    if(when_ArraySlice_l158_141) begin
      if(when_ArraySlice_l159_141) begin
        debug_5_17 = 1'b1;
      end else begin
        debug_5_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_141) begin
        debug_5_17 = 1'b1;
      end else begin
        debug_5_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_17 = 1'b0;
    if(when_ArraySlice_l158_142) begin
      if(when_ArraySlice_l159_142) begin
        debug_6_17 = 1'b1;
      end else begin
        debug_6_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_142) begin
        debug_6_17 = 1'b1;
      end else begin
        debug_6_17 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_17 = 1'b0;
    if(when_ArraySlice_l158_143) begin
      if(when_ArraySlice_l159_143) begin
        debug_7_17 = 1'b1;
      end else begin
        debug_7_17 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_143) begin
        debug_7_17 = 1'b1;
      end else begin
        debug_7_17 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_136 = (_zz_when_ArraySlice_l158_136 <= _zz_when_ArraySlice_l158_136_3);
  assign when_ArraySlice_l159_136 = (_zz_when_ArraySlice_l159_136 <= _zz_when_ArraySlice_l159_136_1);
  assign _zz_realValue_0_136 = (_zz__zz_realValue_0_136 % _zz__zz_realValue_0_136_1);
  assign when_ArraySlice_l110_136 = (_zz_realValue_0_136 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_136) begin
      realValue_0_136 = (_zz_realValue_0_136_1 - _zz_realValue_0_136);
    end else begin
      realValue_0_136 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_136 = (_zz_when_ArraySlice_l166_136 <= _zz_when_ArraySlice_l166_136_1);
  assign when_ArraySlice_l158_137 = (_zz_when_ArraySlice_l158_137 <= _zz_when_ArraySlice_l158_137_3);
  assign when_ArraySlice_l159_137 = (_zz_when_ArraySlice_l159_137 <= _zz_when_ArraySlice_l159_137_2);
  assign _zz_realValue_0_137 = (_zz__zz_realValue_0_137 % _zz__zz_realValue_0_137_1);
  assign when_ArraySlice_l110_137 = (_zz_realValue_0_137 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_137) begin
      realValue_0_137 = (_zz_realValue_0_137_1 - _zz_realValue_0_137);
    end else begin
      realValue_0_137 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_137 = (_zz_when_ArraySlice_l166_137 <= _zz_when_ArraySlice_l166_137_2);
  assign when_ArraySlice_l158_138 = (_zz_when_ArraySlice_l158_138 <= _zz_when_ArraySlice_l158_138_3);
  assign when_ArraySlice_l159_138 = (_zz_when_ArraySlice_l159_138 <= _zz_when_ArraySlice_l159_138_2);
  assign _zz_realValue_0_138 = (_zz__zz_realValue_0_138 % _zz__zz_realValue_0_138_1);
  assign when_ArraySlice_l110_138 = (_zz_realValue_0_138 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_138) begin
      realValue_0_138 = (_zz_realValue_0_138_1 - _zz_realValue_0_138);
    end else begin
      realValue_0_138 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_138 = (_zz_when_ArraySlice_l166_138 <= _zz_when_ArraySlice_l166_138_2);
  assign when_ArraySlice_l158_139 = (_zz_when_ArraySlice_l158_139 <= _zz_when_ArraySlice_l158_139_3);
  assign when_ArraySlice_l159_139 = (_zz_when_ArraySlice_l159_139 <= _zz_when_ArraySlice_l159_139_2);
  assign _zz_realValue_0_139 = (_zz__zz_realValue_0_139 % _zz__zz_realValue_0_139_1);
  assign when_ArraySlice_l110_139 = (_zz_realValue_0_139 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_139) begin
      realValue_0_139 = (_zz_realValue_0_139_1 - _zz_realValue_0_139);
    end else begin
      realValue_0_139 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_139 = (_zz_when_ArraySlice_l166_139 <= _zz_when_ArraySlice_l166_139_2);
  assign when_ArraySlice_l158_140 = (_zz_when_ArraySlice_l158_140 <= _zz_when_ArraySlice_l158_140_3);
  assign when_ArraySlice_l159_140 = (_zz_when_ArraySlice_l159_140 <= _zz_when_ArraySlice_l159_140_2);
  assign _zz_realValue_0_140 = (_zz__zz_realValue_0_140 % _zz__zz_realValue_0_140_1);
  assign when_ArraySlice_l110_140 = (_zz_realValue_0_140 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_140) begin
      realValue_0_140 = (_zz_realValue_0_140_1 - _zz_realValue_0_140);
    end else begin
      realValue_0_140 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_140 = (_zz_when_ArraySlice_l166_140 <= _zz_when_ArraySlice_l166_140_2);
  assign when_ArraySlice_l158_141 = (_zz_when_ArraySlice_l158_141 <= _zz_when_ArraySlice_l158_141_3);
  assign when_ArraySlice_l159_141 = (_zz_when_ArraySlice_l159_141 <= _zz_when_ArraySlice_l159_141_2);
  assign _zz_realValue_0_141 = (_zz__zz_realValue_0_141 % _zz__zz_realValue_0_141_1);
  assign when_ArraySlice_l110_141 = (_zz_realValue_0_141 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_141) begin
      realValue_0_141 = (_zz_realValue_0_141_1 - _zz_realValue_0_141);
    end else begin
      realValue_0_141 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_141 = (_zz_when_ArraySlice_l166_141 <= _zz_when_ArraySlice_l166_141_2);
  assign when_ArraySlice_l158_142 = (_zz_when_ArraySlice_l158_142 <= _zz_when_ArraySlice_l158_142_3);
  assign when_ArraySlice_l159_142 = (_zz_when_ArraySlice_l159_142 <= _zz_when_ArraySlice_l159_142_2);
  assign _zz_realValue_0_142 = (_zz__zz_realValue_0_142 % _zz__zz_realValue_0_142_1);
  assign when_ArraySlice_l110_142 = (_zz_realValue_0_142 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_142) begin
      realValue_0_142 = (_zz_realValue_0_142_1 - _zz_realValue_0_142);
    end else begin
      realValue_0_142 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_142 = (_zz_when_ArraySlice_l166_142 <= _zz_when_ArraySlice_l166_142_2);
  assign when_ArraySlice_l158_143 = (_zz_when_ArraySlice_l158_143 <= _zz_when_ArraySlice_l158_143_3);
  assign when_ArraySlice_l159_143 = (_zz_when_ArraySlice_l159_143 <= _zz_when_ArraySlice_l159_143_2);
  assign _zz_realValue_0_143 = (_zz__zz_realValue_0_143 % _zz__zz_realValue_0_143_1);
  assign when_ArraySlice_l110_143 = (_zz_realValue_0_143 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_143) begin
      realValue_0_143 = (_zz_realValue_0_143_1 - _zz_realValue_0_143);
    end else begin
      realValue_0_143 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_143 = (_zz_when_ArraySlice_l166_143 <= _zz_when_ArraySlice_l166_143_2);
  assign when_ArraySlice_l425_5 = (! ((((((_zz_when_ArraySlice_l425_5_1 && _zz_when_ArraySlice_l425_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l425_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_5_4 && _zz_when_ArraySlice_l425_5_5) && (debug_4_17 == _zz_when_ArraySlice_l425_5_6)) && (debug_5_17 == 1'b1)) && (debug_6_17 == 1'b1)) && (debug_7_17 == 1'b1))));
  assign when_ArraySlice_l428_5 = (_zz_when_ArraySlice_l428_5_1 <= _zz_when_ArraySlice_l428_5_2);
  assign when_ArraySlice_l431_5 = (_zz_when_ArraySlice_l431_5 <= _zz_when_ArraySlice_l431_5_1);
  assign outputStreamArrayData_5_fire_3 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l438_5 = ((_zz_when_ArraySlice_l438_5 == 13'h0) && outputStreamArrayData_5_fire_3);
  assign outputStreamArrayData_5_fire_4 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l449_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l449_5) && outputStreamArrayData_5_fire_4);
  assign _zz_realValue1_0_17 = (_zz__zz_realValue1_0_17 % _zz__zz_realValue1_0_17_1);
  assign when_ArraySlice_l95_17 = (_zz_realValue1_0_17 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_17) begin
      realValue1_0_17 = (_zz_realValue1_0_17_1 - _zz_realValue1_0_17);
    end else begin
      realValue1_0_17 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_5 = (_zz_when_ArraySlice_l450_5 < _zz_when_ArraySlice_l450_5_2);
  always @(*) begin
    debug_0_18 = 1'b0;
    if(when_ArraySlice_l158_144) begin
      if(when_ArraySlice_l159_144) begin
        debug_0_18 = 1'b1;
      end else begin
        debug_0_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_144) begin
        debug_0_18 = 1'b1;
      end else begin
        debug_0_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_18 = 1'b0;
    if(when_ArraySlice_l158_145) begin
      if(when_ArraySlice_l159_145) begin
        debug_1_18 = 1'b1;
      end else begin
        debug_1_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_145) begin
        debug_1_18 = 1'b1;
      end else begin
        debug_1_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_18 = 1'b0;
    if(when_ArraySlice_l158_146) begin
      if(when_ArraySlice_l159_146) begin
        debug_2_18 = 1'b1;
      end else begin
        debug_2_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_146) begin
        debug_2_18 = 1'b1;
      end else begin
        debug_2_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_18 = 1'b0;
    if(when_ArraySlice_l158_147) begin
      if(when_ArraySlice_l159_147) begin
        debug_3_18 = 1'b1;
      end else begin
        debug_3_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_147) begin
        debug_3_18 = 1'b1;
      end else begin
        debug_3_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_18 = 1'b0;
    if(when_ArraySlice_l158_148) begin
      if(when_ArraySlice_l159_148) begin
        debug_4_18 = 1'b1;
      end else begin
        debug_4_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_148) begin
        debug_4_18 = 1'b1;
      end else begin
        debug_4_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_18 = 1'b0;
    if(when_ArraySlice_l158_149) begin
      if(when_ArraySlice_l159_149) begin
        debug_5_18 = 1'b1;
      end else begin
        debug_5_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_149) begin
        debug_5_18 = 1'b1;
      end else begin
        debug_5_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_18 = 1'b0;
    if(when_ArraySlice_l158_150) begin
      if(when_ArraySlice_l159_150) begin
        debug_6_18 = 1'b1;
      end else begin
        debug_6_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_150) begin
        debug_6_18 = 1'b1;
      end else begin
        debug_6_18 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_18 = 1'b0;
    if(when_ArraySlice_l158_151) begin
      if(when_ArraySlice_l159_151) begin
        debug_7_18 = 1'b1;
      end else begin
        debug_7_18 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_151) begin
        debug_7_18 = 1'b1;
      end else begin
        debug_7_18 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_144 = (_zz_when_ArraySlice_l158_144 <= _zz_when_ArraySlice_l158_144_3);
  assign when_ArraySlice_l159_144 = (_zz_when_ArraySlice_l159_144 <= _zz_when_ArraySlice_l159_144_1);
  assign _zz_realValue_0_144 = (_zz__zz_realValue_0_144 % _zz__zz_realValue_0_144_1);
  assign when_ArraySlice_l110_144 = (_zz_realValue_0_144 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_144) begin
      realValue_0_144 = (_zz_realValue_0_144_1 - _zz_realValue_0_144);
    end else begin
      realValue_0_144 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_144 = (_zz_when_ArraySlice_l166_144 <= _zz_when_ArraySlice_l166_144_1);
  assign when_ArraySlice_l158_145 = (_zz_when_ArraySlice_l158_145 <= _zz_when_ArraySlice_l158_145_3);
  assign when_ArraySlice_l159_145 = (_zz_when_ArraySlice_l159_145 <= _zz_when_ArraySlice_l159_145_2);
  assign _zz_realValue_0_145 = (_zz__zz_realValue_0_145 % _zz__zz_realValue_0_145_1);
  assign when_ArraySlice_l110_145 = (_zz_realValue_0_145 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_145) begin
      realValue_0_145 = (_zz_realValue_0_145_1 - _zz_realValue_0_145);
    end else begin
      realValue_0_145 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_145 = (_zz_when_ArraySlice_l166_145 <= _zz_when_ArraySlice_l166_145_2);
  assign when_ArraySlice_l158_146 = (_zz_when_ArraySlice_l158_146 <= _zz_when_ArraySlice_l158_146_3);
  assign when_ArraySlice_l159_146 = (_zz_when_ArraySlice_l159_146 <= _zz_when_ArraySlice_l159_146_2);
  assign _zz_realValue_0_146 = (_zz__zz_realValue_0_146 % _zz__zz_realValue_0_146_1);
  assign when_ArraySlice_l110_146 = (_zz_realValue_0_146 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_146) begin
      realValue_0_146 = (_zz_realValue_0_146_1 - _zz_realValue_0_146);
    end else begin
      realValue_0_146 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_146 = (_zz_when_ArraySlice_l166_146 <= _zz_when_ArraySlice_l166_146_2);
  assign when_ArraySlice_l158_147 = (_zz_when_ArraySlice_l158_147 <= _zz_when_ArraySlice_l158_147_3);
  assign when_ArraySlice_l159_147 = (_zz_when_ArraySlice_l159_147 <= _zz_when_ArraySlice_l159_147_2);
  assign _zz_realValue_0_147 = (_zz__zz_realValue_0_147 % _zz__zz_realValue_0_147_1);
  assign when_ArraySlice_l110_147 = (_zz_realValue_0_147 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_147) begin
      realValue_0_147 = (_zz_realValue_0_147_1 - _zz_realValue_0_147);
    end else begin
      realValue_0_147 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_147 = (_zz_when_ArraySlice_l166_147 <= _zz_when_ArraySlice_l166_147_2);
  assign when_ArraySlice_l158_148 = (_zz_when_ArraySlice_l158_148 <= _zz_when_ArraySlice_l158_148_3);
  assign when_ArraySlice_l159_148 = (_zz_when_ArraySlice_l159_148 <= _zz_when_ArraySlice_l159_148_2);
  assign _zz_realValue_0_148 = (_zz__zz_realValue_0_148 % _zz__zz_realValue_0_148_1);
  assign when_ArraySlice_l110_148 = (_zz_realValue_0_148 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_148) begin
      realValue_0_148 = (_zz_realValue_0_148_1 - _zz_realValue_0_148);
    end else begin
      realValue_0_148 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_148 = (_zz_when_ArraySlice_l166_148 <= _zz_when_ArraySlice_l166_148_2);
  assign when_ArraySlice_l158_149 = (_zz_when_ArraySlice_l158_149 <= _zz_when_ArraySlice_l158_149_3);
  assign when_ArraySlice_l159_149 = (_zz_when_ArraySlice_l159_149 <= _zz_when_ArraySlice_l159_149_2);
  assign _zz_realValue_0_149 = (_zz__zz_realValue_0_149 % _zz__zz_realValue_0_149_1);
  assign when_ArraySlice_l110_149 = (_zz_realValue_0_149 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_149) begin
      realValue_0_149 = (_zz_realValue_0_149_1 - _zz_realValue_0_149);
    end else begin
      realValue_0_149 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_149 = (_zz_when_ArraySlice_l166_149 <= _zz_when_ArraySlice_l166_149_2);
  assign when_ArraySlice_l158_150 = (_zz_when_ArraySlice_l158_150 <= _zz_when_ArraySlice_l158_150_3);
  assign when_ArraySlice_l159_150 = (_zz_when_ArraySlice_l159_150 <= _zz_when_ArraySlice_l159_150_2);
  assign _zz_realValue_0_150 = (_zz__zz_realValue_0_150 % _zz__zz_realValue_0_150_1);
  assign when_ArraySlice_l110_150 = (_zz_realValue_0_150 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_150) begin
      realValue_0_150 = (_zz_realValue_0_150_1 - _zz_realValue_0_150);
    end else begin
      realValue_0_150 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_150 = (_zz_when_ArraySlice_l166_150 <= _zz_when_ArraySlice_l166_150_2);
  assign when_ArraySlice_l158_151 = (_zz_when_ArraySlice_l158_151 <= _zz_when_ArraySlice_l158_151_3);
  assign when_ArraySlice_l159_151 = (_zz_when_ArraySlice_l159_151 <= _zz_when_ArraySlice_l159_151_2);
  assign _zz_realValue_0_151 = (_zz__zz_realValue_0_151 % _zz__zz_realValue_0_151_1);
  assign when_ArraySlice_l110_151 = (_zz_realValue_0_151 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_151) begin
      realValue_0_151 = (_zz_realValue_0_151_1 - _zz_realValue_0_151);
    end else begin
      realValue_0_151 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_151 = (_zz_when_ArraySlice_l166_151 <= _zz_when_ArraySlice_l166_151_2);
  assign when_ArraySlice_l457_5 = (! ((((((_zz_when_ArraySlice_l457_5_1 && _zz_when_ArraySlice_l457_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l457_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_5_4 && _zz_when_ArraySlice_l457_5_5) && (debug_4_18 == _zz_when_ArraySlice_l457_5_6)) && (debug_5_18 == 1'b1)) && (debug_6_18 == 1'b1)) && (debug_7_18 == 1'b1))));
  assign outputStreamArrayData_5_fire_5 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l461_5 = ((_zz_when_ArraySlice_l461_5 == 13'h0) && outputStreamArrayData_5_fire_5);
  assign when_ArraySlice_l447_5 = (allowPadding_5 && (_zz_when_ArraySlice_l447_5 <= _zz_when_ArraySlice_l447_5_1));
  assign outputStreamArrayData_5_fire_6 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l468_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l468_5);
  assign when_ArraySlice_l376_6 = (_zz_when_ArraySlice_l376_6 < _zz_when_ArraySlice_l376_6_3);
  assign when_ArraySlice_l377_6 = ((! holdReadOp_6) && (_zz_when_ArraySlice_l377_6 != 7'h0));
  assign _zz_outputStreamArrayData_6_valid = (selectReadFifo_6 + _zz__zz_outputStreamArrayData_6_valid);
  assign _zz_9 = ({127'd0,1'b1} <<< _zz__zz_9);
  assign _zz_io_pop_ready_6 = outputStreamArrayData_6_ready;
  assign when_ArraySlice_l382_6 = (! holdReadOp_6);
  assign outputStreamArrayData_6_fire = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l383_6 = ((7'h01 < _zz_when_ArraySlice_l383_6) && outputStreamArrayData_6_fire);
  assign when_ArraySlice_l384_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l384_6);
  assign when_ArraySlice_l387_6 = (_zz_when_ArraySlice_l387_6 == 13'h0);
  assign outputStreamArrayData_6_fire_1 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l392_6 = ((_zz_when_ArraySlice_l392_6 == 7'h01) && outputStreamArrayData_6_fire_1);
  assign when_ArraySlice_l393_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l393_6);
  assign _zz_realValue1_0_18 = (_zz__zz_realValue1_0_18 % _zz__zz_realValue1_0_18_1);
  assign when_ArraySlice_l95_18 = (_zz_realValue1_0_18 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_18) begin
      realValue1_0_18 = (_zz_realValue1_0_18_1 - _zz_realValue1_0_18);
    end else begin
      realValue1_0_18 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_6 = (_zz_when_ArraySlice_l395_6 < _zz_when_ArraySlice_l395_6_2);
  always @(*) begin
    debug_0_19 = 1'b0;
    if(when_ArraySlice_l158_152) begin
      if(when_ArraySlice_l159_152) begin
        debug_0_19 = 1'b1;
      end else begin
        debug_0_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_152) begin
        debug_0_19 = 1'b1;
      end else begin
        debug_0_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_19 = 1'b0;
    if(when_ArraySlice_l158_153) begin
      if(when_ArraySlice_l159_153) begin
        debug_1_19 = 1'b1;
      end else begin
        debug_1_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_153) begin
        debug_1_19 = 1'b1;
      end else begin
        debug_1_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_19 = 1'b0;
    if(when_ArraySlice_l158_154) begin
      if(when_ArraySlice_l159_154) begin
        debug_2_19 = 1'b1;
      end else begin
        debug_2_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_154) begin
        debug_2_19 = 1'b1;
      end else begin
        debug_2_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_19 = 1'b0;
    if(when_ArraySlice_l158_155) begin
      if(when_ArraySlice_l159_155) begin
        debug_3_19 = 1'b1;
      end else begin
        debug_3_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_155) begin
        debug_3_19 = 1'b1;
      end else begin
        debug_3_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_19 = 1'b0;
    if(when_ArraySlice_l158_156) begin
      if(when_ArraySlice_l159_156) begin
        debug_4_19 = 1'b1;
      end else begin
        debug_4_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_156) begin
        debug_4_19 = 1'b1;
      end else begin
        debug_4_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_19 = 1'b0;
    if(when_ArraySlice_l158_157) begin
      if(when_ArraySlice_l159_157) begin
        debug_5_19 = 1'b1;
      end else begin
        debug_5_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_157) begin
        debug_5_19 = 1'b1;
      end else begin
        debug_5_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_19 = 1'b0;
    if(when_ArraySlice_l158_158) begin
      if(when_ArraySlice_l159_158) begin
        debug_6_19 = 1'b1;
      end else begin
        debug_6_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_158) begin
        debug_6_19 = 1'b1;
      end else begin
        debug_6_19 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_19 = 1'b0;
    if(when_ArraySlice_l158_159) begin
      if(when_ArraySlice_l159_159) begin
        debug_7_19 = 1'b1;
      end else begin
        debug_7_19 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_159) begin
        debug_7_19 = 1'b1;
      end else begin
        debug_7_19 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_152 = (_zz_when_ArraySlice_l158_152 <= _zz_when_ArraySlice_l158_152_3);
  assign when_ArraySlice_l159_152 = (_zz_when_ArraySlice_l159_152 <= _zz_when_ArraySlice_l159_152_1);
  assign _zz_realValue_0_152 = (_zz__zz_realValue_0_152 % _zz__zz_realValue_0_152_1);
  assign when_ArraySlice_l110_152 = (_zz_realValue_0_152 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_152) begin
      realValue_0_152 = (_zz_realValue_0_152_1 - _zz_realValue_0_152);
    end else begin
      realValue_0_152 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_152 = (_zz_when_ArraySlice_l166_152 <= _zz_when_ArraySlice_l166_152_1);
  assign when_ArraySlice_l158_153 = (_zz_when_ArraySlice_l158_153 <= _zz_when_ArraySlice_l158_153_3);
  assign when_ArraySlice_l159_153 = (_zz_when_ArraySlice_l159_153 <= _zz_when_ArraySlice_l159_153_2);
  assign _zz_realValue_0_153 = (_zz__zz_realValue_0_153 % _zz__zz_realValue_0_153_1);
  assign when_ArraySlice_l110_153 = (_zz_realValue_0_153 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_153) begin
      realValue_0_153 = (_zz_realValue_0_153_1 - _zz_realValue_0_153);
    end else begin
      realValue_0_153 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_153 = (_zz_when_ArraySlice_l166_153 <= _zz_when_ArraySlice_l166_153_2);
  assign when_ArraySlice_l158_154 = (_zz_when_ArraySlice_l158_154 <= _zz_when_ArraySlice_l158_154_3);
  assign when_ArraySlice_l159_154 = (_zz_when_ArraySlice_l159_154 <= _zz_when_ArraySlice_l159_154_2);
  assign _zz_realValue_0_154 = (_zz__zz_realValue_0_154 % _zz__zz_realValue_0_154_1);
  assign when_ArraySlice_l110_154 = (_zz_realValue_0_154 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_154) begin
      realValue_0_154 = (_zz_realValue_0_154_1 - _zz_realValue_0_154);
    end else begin
      realValue_0_154 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_154 = (_zz_when_ArraySlice_l166_154 <= _zz_when_ArraySlice_l166_154_2);
  assign when_ArraySlice_l158_155 = (_zz_when_ArraySlice_l158_155 <= _zz_when_ArraySlice_l158_155_3);
  assign when_ArraySlice_l159_155 = (_zz_when_ArraySlice_l159_155 <= _zz_when_ArraySlice_l159_155_2);
  assign _zz_realValue_0_155 = (_zz__zz_realValue_0_155 % _zz__zz_realValue_0_155_1);
  assign when_ArraySlice_l110_155 = (_zz_realValue_0_155 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_155) begin
      realValue_0_155 = (_zz_realValue_0_155_1 - _zz_realValue_0_155);
    end else begin
      realValue_0_155 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_155 = (_zz_when_ArraySlice_l166_155 <= _zz_when_ArraySlice_l166_155_2);
  assign when_ArraySlice_l158_156 = (_zz_when_ArraySlice_l158_156 <= _zz_when_ArraySlice_l158_156_3);
  assign when_ArraySlice_l159_156 = (_zz_when_ArraySlice_l159_156 <= _zz_when_ArraySlice_l159_156_2);
  assign _zz_realValue_0_156 = (_zz__zz_realValue_0_156 % _zz__zz_realValue_0_156_1);
  assign when_ArraySlice_l110_156 = (_zz_realValue_0_156 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_156) begin
      realValue_0_156 = (_zz_realValue_0_156_1 - _zz_realValue_0_156);
    end else begin
      realValue_0_156 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_156 = (_zz_when_ArraySlice_l166_156 <= _zz_when_ArraySlice_l166_156_2);
  assign when_ArraySlice_l158_157 = (_zz_when_ArraySlice_l158_157 <= _zz_when_ArraySlice_l158_157_3);
  assign when_ArraySlice_l159_157 = (_zz_when_ArraySlice_l159_157 <= _zz_when_ArraySlice_l159_157_2);
  assign _zz_realValue_0_157 = (_zz__zz_realValue_0_157 % _zz__zz_realValue_0_157_1);
  assign when_ArraySlice_l110_157 = (_zz_realValue_0_157 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_157) begin
      realValue_0_157 = (_zz_realValue_0_157_1 - _zz_realValue_0_157);
    end else begin
      realValue_0_157 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_157 = (_zz_when_ArraySlice_l166_157 <= _zz_when_ArraySlice_l166_157_2);
  assign when_ArraySlice_l158_158 = (_zz_when_ArraySlice_l158_158 <= _zz_when_ArraySlice_l158_158_3);
  assign when_ArraySlice_l159_158 = (_zz_when_ArraySlice_l159_158 <= _zz_when_ArraySlice_l159_158_2);
  assign _zz_realValue_0_158 = (_zz__zz_realValue_0_158 % _zz__zz_realValue_0_158_1);
  assign when_ArraySlice_l110_158 = (_zz_realValue_0_158 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_158) begin
      realValue_0_158 = (_zz_realValue_0_158_1 - _zz_realValue_0_158);
    end else begin
      realValue_0_158 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_158 = (_zz_when_ArraySlice_l166_158 <= _zz_when_ArraySlice_l166_158_2);
  assign when_ArraySlice_l158_159 = (_zz_when_ArraySlice_l158_159 <= _zz_when_ArraySlice_l158_159_3);
  assign when_ArraySlice_l159_159 = (_zz_when_ArraySlice_l159_159 <= _zz_when_ArraySlice_l159_159_2);
  assign _zz_realValue_0_159 = (_zz__zz_realValue_0_159 % _zz__zz_realValue_0_159_1);
  assign when_ArraySlice_l110_159 = (_zz_realValue_0_159 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_159) begin
      realValue_0_159 = (_zz_realValue_0_159_1 - _zz_realValue_0_159);
    end else begin
      realValue_0_159 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_159 = (_zz_when_ArraySlice_l166_159 <= _zz_when_ArraySlice_l166_159_2);
  assign when_ArraySlice_l400_6 = (! ((((((_zz_when_ArraySlice_l400_6_1 && _zz_when_ArraySlice_l400_6_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_6_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_6_4 && _zz_when_ArraySlice_l400_6_5) && (debug_4_19 == _zz_when_ArraySlice_l400_6_6)) && (debug_5_19 == 1'b1)) && (debug_6_19 == 1'b1)) && (debug_7_19 == 1'b1))));
  assign when_ArraySlice_l403_6 = (_zz_when_ArraySlice_l403_6_1 <= _zz_when_ArraySlice_l403_6_2);
  assign when_ArraySlice_l406_6 = (_zz_when_ArraySlice_l406_6 <= _zz_when_ArraySlice_l406_6_1);
  assign when_ArraySlice_l413_6 = (_zz_when_ArraySlice_l413_6 == 13'h0);
  assign when_ArraySlice_l417_6 = (_zz_when_ArraySlice_l417_6 == 7'h0);
  assign outputStreamArrayData_6_fire_2 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l418_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l418_6) && outputStreamArrayData_6_fire_2);
  assign _zz_realValue1_0_19 = (_zz__zz_realValue1_0_19 % _zz__zz_realValue1_0_19_1);
  assign when_ArraySlice_l95_19 = (_zz_realValue1_0_19 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_19) begin
      realValue1_0_19 = (_zz_realValue1_0_19_1 - _zz_realValue1_0_19);
    end else begin
      realValue1_0_19 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_6 = (_zz_when_ArraySlice_l420_6 < _zz_when_ArraySlice_l420_6_2);
  always @(*) begin
    debug_0_20 = 1'b0;
    if(when_ArraySlice_l158_160) begin
      if(when_ArraySlice_l159_160) begin
        debug_0_20 = 1'b1;
      end else begin
        debug_0_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_160) begin
        debug_0_20 = 1'b1;
      end else begin
        debug_0_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_20 = 1'b0;
    if(when_ArraySlice_l158_161) begin
      if(when_ArraySlice_l159_161) begin
        debug_1_20 = 1'b1;
      end else begin
        debug_1_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_161) begin
        debug_1_20 = 1'b1;
      end else begin
        debug_1_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_20 = 1'b0;
    if(when_ArraySlice_l158_162) begin
      if(when_ArraySlice_l159_162) begin
        debug_2_20 = 1'b1;
      end else begin
        debug_2_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_162) begin
        debug_2_20 = 1'b1;
      end else begin
        debug_2_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_20 = 1'b0;
    if(when_ArraySlice_l158_163) begin
      if(when_ArraySlice_l159_163) begin
        debug_3_20 = 1'b1;
      end else begin
        debug_3_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_163) begin
        debug_3_20 = 1'b1;
      end else begin
        debug_3_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_20 = 1'b0;
    if(when_ArraySlice_l158_164) begin
      if(when_ArraySlice_l159_164) begin
        debug_4_20 = 1'b1;
      end else begin
        debug_4_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_164) begin
        debug_4_20 = 1'b1;
      end else begin
        debug_4_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_20 = 1'b0;
    if(when_ArraySlice_l158_165) begin
      if(when_ArraySlice_l159_165) begin
        debug_5_20 = 1'b1;
      end else begin
        debug_5_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_165) begin
        debug_5_20 = 1'b1;
      end else begin
        debug_5_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_20 = 1'b0;
    if(when_ArraySlice_l158_166) begin
      if(when_ArraySlice_l159_166) begin
        debug_6_20 = 1'b1;
      end else begin
        debug_6_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_166) begin
        debug_6_20 = 1'b1;
      end else begin
        debug_6_20 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_20 = 1'b0;
    if(when_ArraySlice_l158_167) begin
      if(when_ArraySlice_l159_167) begin
        debug_7_20 = 1'b1;
      end else begin
        debug_7_20 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_167) begin
        debug_7_20 = 1'b1;
      end else begin
        debug_7_20 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_160 = (_zz_when_ArraySlice_l158_160 <= _zz_when_ArraySlice_l158_160_3);
  assign when_ArraySlice_l159_160 = (_zz_when_ArraySlice_l159_160 <= _zz_when_ArraySlice_l159_160_1);
  assign _zz_realValue_0_160 = (_zz__zz_realValue_0_160 % _zz__zz_realValue_0_160_1);
  assign when_ArraySlice_l110_160 = (_zz_realValue_0_160 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_160) begin
      realValue_0_160 = (_zz_realValue_0_160_1 - _zz_realValue_0_160);
    end else begin
      realValue_0_160 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_160 = (_zz_when_ArraySlice_l166_160 <= _zz_when_ArraySlice_l166_160_1);
  assign when_ArraySlice_l158_161 = (_zz_when_ArraySlice_l158_161 <= _zz_when_ArraySlice_l158_161_3);
  assign when_ArraySlice_l159_161 = (_zz_when_ArraySlice_l159_161 <= _zz_when_ArraySlice_l159_161_2);
  assign _zz_realValue_0_161 = (_zz__zz_realValue_0_161 % _zz__zz_realValue_0_161_1);
  assign when_ArraySlice_l110_161 = (_zz_realValue_0_161 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_161) begin
      realValue_0_161 = (_zz_realValue_0_161_1 - _zz_realValue_0_161);
    end else begin
      realValue_0_161 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_161 = (_zz_when_ArraySlice_l166_161 <= _zz_when_ArraySlice_l166_161_2);
  assign when_ArraySlice_l158_162 = (_zz_when_ArraySlice_l158_162 <= _zz_when_ArraySlice_l158_162_3);
  assign when_ArraySlice_l159_162 = (_zz_when_ArraySlice_l159_162 <= _zz_when_ArraySlice_l159_162_2);
  assign _zz_realValue_0_162 = (_zz__zz_realValue_0_162 % _zz__zz_realValue_0_162_1);
  assign when_ArraySlice_l110_162 = (_zz_realValue_0_162 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_162) begin
      realValue_0_162 = (_zz_realValue_0_162_1 - _zz_realValue_0_162);
    end else begin
      realValue_0_162 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_162 = (_zz_when_ArraySlice_l166_162 <= _zz_when_ArraySlice_l166_162_2);
  assign when_ArraySlice_l158_163 = (_zz_when_ArraySlice_l158_163 <= _zz_when_ArraySlice_l158_163_3);
  assign when_ArraySlice_l159_163 = (_zz_when_ArraySlice_l159_163 <= _zz_when_ArraySlice_l159_163_2);
  assign _zz_realValue_0_163 = (_zz__zz_realValue_0_163 % _zz__zz_realValue_0_163_1);
  assign when_ArraySlice_l110_163 = (_zz_realValue_0_163 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_163) begin
      realValue_0_163 = (_zz_realValue_0_163_1 - _zz_realValue_0_163);
    end else begin
      realValue_0_163 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_163 = (_zz_when_ArraySlice_l166_163 <= _zz_when_ArraySlice_l166_163_2);
  assign when_ArraySlice_l158_164 = (_zz_when_ArraySlice_l158_164 <= _zz_when_ArraySlice_l158_164_3);
  assign when_ArraySlice_l159_164 = (_zz_when_ArraySlice_l159_164 <= _zz_when_ArraySlice_l159_164_2);
  assign _zz_realValue_0_164 = (_zz__zz_realValue_0_164 % _zz__zz_realValue_0_164_1);
  assign when_ArraySlice_l110_164 = (_zz_realValue_0_164 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_164) begin
      realValue_0_164 = (_zz_realValue_0_164_1 - _zz_realValue_0_164);
    end else begin
      realValue_0_164 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_164 = (_zz_when_ArraySlice_l166_164 <= _zz_when_ArraySlice_l166_164_2);
  assign when_ArraySlice_l158_165 = (_zz_when_ArraySlice_l158_165 <= _zz_when_ArraySlice_l158_165_3);
  assign when_ArraySlice_l159_165 = (_zz_when_ArraySlice_l159_165 <= _zz_when_ArraySlice_l159_165_2);
  assign _zz_realValue_0_165 = (_zz__zz_realValue_0_165 % _zz__zz_realValue_0_165_1);
  assign when_ArraySlice_l110_165 = (_zz_realValue_0_165 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_165) begin
      realValue_0_165 = (_zz_realValue_0_165_1 - _zz_realValue_0_165);
    end else begin
      realValue_0_165 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_165 = (_zz_when_ArraySlice_l166_165 <= _zz_when_ArraySlice_l166_165_2);
  assign when_ArraySlice_l158_166 = (_zz_when_ArraySlice_l158_166 <= _zz_when_ArraySlice_l158_166_3);
  assign when_ArraySlice_l159_166 = (_zz_when_ArraySlice_l159_166 <= _zz_when_ArraySlice_l159_166_2);
  assign _zz_realValue_0_166 = (_zz__zz_realValue_0_166 % _zz__zz_realValue_0_166_1);
  assign when_ArraySlice_l110_166 = (_zz_realValue_0_166 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_166) begin
      realValue_0_166 = (_zz_realValue_0_166_1 - _zz_realValue_0_166);
    end else begin
      realValue_0_166 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_166 = (_zz_when_ArraySlice_l166_166 <= _zz_when_ArraySlice_l166_166_2);
  assign when_ArraySlice_l158_167 = (_zz_when_ArraySlice_l158_167 <= _zz_when_ArraySlice_l158_167_3);
  assign when_ArraySlice_l159_167 = (_zz_when_ArraySlice_l159_167 <= _zz_when_ArraySlice_l159_167_2);
  assign _zz_realValue_0_167 = (_zz__zz_realValue_0_167 % _zz__zz_realValue_0_167_1);
  assign when_ArraySlice_l110_167 = (_zz_realValue_0_167 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_167) begin
      realValue_0_167 = (_zz_realValue_0_167_1 - _zz_realValue_0_167);
    end else begin
      realValue_0_167 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_167 = (_zz_when_ArraySlice_l166_167 <= _zz_when_ArraySlice_l166_167_2);
  assign when_ArraySlice_l425_6 = (! ((((((_zz_when_ArraySlice_l425_6 && _zz_when_ArraySlice_l425_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l425_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_6_3 && _zz_when_ArraySlice_l425_6_4) && (debug_4_20 == _zz_when_ArraySlice_l425_6_5)) && (debug_5_20 == 1'b1)) && (debug_6_20 == 1'b1)) && (debug_7_20 == 1'b1))));
  assign when_ArraySlice_l428_6 = (_zz_when_ArraySlice_l428_6_1 <= _zz_when_ArraySlice_l428_6_2);
  assign when_ArraySlice_l431_6 = (_zz_when_ArraySlice_l431_6 <= _zz_when_ArraySlice_l431_6_1);
  assign outputStreamArrayData_6_fire_3 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l438_6 = ((_zz_when_ArraySlice_l438_6 == 13'h0) && outputStreamArrayData_6_fire_3);
  assign outputStreamArrayData_6_fire_4 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l449_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l449_6) && outputStreamArrayData_6_fire_4);
  assign _zz_realValue1_0_20 = (_zz__zz_realValue1_0_20 % _zz__zz_realValue1_0_20_1);
  assign when_ArraySlice_l95_20 = (_zz_realValue1_0_20 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_20) begin
      realValue1_0_20 = (_zz_realValue1_0_20_1 - _zz_realValue1_0_20);
    end else begin
      realValue1_0_20 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_6 = (_zz_when_ArraySlice_l450_6 < _zz_when_ArraySlice_l450_6_2);
  always @(*) begin
    debug_0_21 = 1'b0;
    if(when_ArraySlice_l158_168) begin
      if(when_ArraySlice_l159_168) begin
        debug_0_21 = 1'b1;
      end else begin
        debug_0_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_168) begin
        debug_0_21 = 1'b1;
      end else begin
        debug_0_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_21 = 1'b0;
    if(when_ArraySlice_l158_169) begin
      if(when_ArraySlice_l159_169) begin
        debug_1_21 = 1'b1;
      end else begin
        debug_1_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_169) begin
        debug_1_21 = 1'b1;
      end else begin
        debug_1_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_21 = 1'b0;
    if(when_ArraySlice_l158_170) begin
      if(when_ArraySlice_l159_170) begin
        debug_2_21 = 1'b1;
      end else begin
        debug_2_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_170) begin
        debug_2_21 = 1'b1;
      end else begin
        debug_2_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_21 = 1'b0;
    if(when_ArraySlice_l158_171) begin
      if(when_ArraySlice_l159_171) begin
        debug_3_21 = 1'b1;
      end else begin
        debug_3_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_171) begin
        debug_3_21 = 1'b1;
      end else begin
        debug_3_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_21 = 1'b0;
    if(when_ArraySlice_l158_172) begin
      if(when_ArraySlice_l159_172) begin
        debug_4_21 = 1'b1;
      end else begin
        debug_4_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_172) begin
        debug_4_21 = 1'b1;
      end else begin
        debug_4_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_21 = 1'b0;
    if(when_ArraySlice_l158_173) begin
      if(when_ArraySlice_l159_173) begin
        debug_5_21 = 1'b1;
      end else begin
        debug_5_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_173) begin
        debug_5_21 = 1'b1;
      end else begin
        debug_5_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_21 = 1'b0;
    if(when_ArraySlice_l158_174) begin
      if(when_ArraySlice_l159_174) begin
        debug_6_21 = 1'b1;
      end else begin
        debug_6_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_174) begin
        debug_6_21 = 1'b1;
      end else begin
        debug_6_21 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_21 = 1'b0;
    if(when_ArraySlice_l158_175) begin
      if(when_ArraySlice_l159_175) begin
        debug_7_21 = 1'b1;
      end else begin
        debug_7_21 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_175) begin
        debug_7_21 = 1'b1;
      end else begin
        debug_7_21 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_168 = (_zz_when_ArraySlice_l158_168 <= _zz_when_ArraySlice_l158_168_3);
  assign when_ArraySlice_l159_168 = (_zz_when_ArraySlice_l159_168 <= _zz_when_ArraySlice_l159_168_1);
  assign _zz_realValue_0_168 = (_zz__zz_realValue_0_168 % _zz__zz_realValue_0_168_1);
  assign when_ArraySlice_l110_168 = (_zz_realValue_0_168 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_168) begin
      realValue_0_168 = (_zz_realValue_0_168_1 - _zz_realValue_0_168);
    end else begin
      realValue_0_168 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_168 = (_zz_when_ArraySlice_l166_168 <= _zz_when_ArraySlice_l166_168_1);
  assign when_ArraySlice_l158_169 = (_zz_when_ArraySlice_l158_169 <= _zz_when_ArraySlice_l158_169_3);
  assign when_ArraySlice_l159_169 = (_zz_when_ArraySlice_l159_169 <= _zz_when_ArraySlice_l159_169_2);
  assign _zz_realValue_0_169 = (_zz__zz_realValue_0_169 % _zz__zz_realValue_0_169_1);
  assign when_ArraySlice_l110_169 = (_zz_realValue_0_169 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_169) begin
      realValue_0_169 = (_zz_realValue_0_169_1 - _zz_realValue_0_169);
    end else begin
      realValue_0_169 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_169 = (_zz_when_ArraySlice_l166_169 <= _zz_when_ArraySlice_l166_169_2);
  assign when_ArraySlice_l158_170 = (_zz_when_ArraySlice_l158_170 <= _zz_when_ArraySlice_l158_170_3);
  assign when_ArraySlice_l159_170 = (_zz_when_ArraySlice_l159_170 <= _zz_when_ArraySlice_l159_170_2);
  assign _zz_realValue_0_170 = (_zz__zz_realValue_0_170 % _zz__zz_realValue_0_170_1);
  assign when_ArraySlice_l110_170 = (_zz_realValue_0_170 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_170) begin
      realValue_0_170 = (_zz_realValue_0_170_1 - _zz_realValue_0_170);
    end else begin
      realValue_0_170 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_170 = (_zz_when_ArraySlice_l166_170 <= _zz_when_ArraySlice_l166_170_2);
  assign when_ArraySlice_l158_171 = (_zz_when_ArraySlice_l158_171 <= _zz_when_ArraySlice_l158_171_3);
  assign when_ArraySlice_l159_171 = (_zz_when_ArraySlice_l159_171 <= _zz_when_ArraySlice_l159_171_2);
  assign _zz_realValue_0_171 = (_zz__zz_realValue_0_171 % _zz__zz_realValue_0_171_1);
  assign when_ArraySlice_l110_171 = (_zz_realValue_0_171 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_171) begin
      realValue_0_171 = (_zz_realValue_0_171_1 - _zz_realValue_0_171);
    end else begin
      realValue_0_171 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_171 = (_zz_when_ArraySlice_l166_171 <= _zz_when_ArraySlice_l166_171_2);
  assign when_ArraySlice_l158_172 = (_zz_when_ArraySlice_l158_172 <= _zz_when_ArraySlice_l158_172_3);
  assign when_ArraySlice_l159_172 = (_zz_when_ArraySlice_l159_172 <= _zz_when_ArraySlice_l159_172_2);
  assign _zz_realValue_0_172 = (_zz__zz_realValue_0_172 % _zz__zz_realValue_0_172_1);
  assign when_ArraySlice_l110_172 = (_zz_realValue_0_172 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_172) begin
      realValue_0_172 = (_zz_realValue_0_172_1 - _zz_realValue_0_172);
    end else begin
      realValue_0_172 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_172 = (_zz_when_ArraySlice_l166_172 <= _zz_when_ArraySlice_l166_172_2);
  assign when_ArraySlice_l158_173 = (_zz_when_ArraySlice_l158_173 <= _zz_when_ArraySlice_l158_173_3);
  assign when_ArraySlice_l159_173 = (_zz_when_ArraySlice_l159_173 <= _zz_when_ArraySlice_l159_173_2);
  assign _zz_realValue_0_173 = (_zz__zz_realValue_0_173 % _zz__zz_realValue_0_173_1);
  assign when_ArraySlice_l110_173 = (_zz_realValue_0_173 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_173) begin
      realValue_0_173 = (_zz_realValue_0_173_1 - _zz_realValue_0_173);
    end else begin
      realValue_0_173 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_173 = (_zz_when_ArraySlice_l166_173 <= _zz_when_ArraySlice_l166_173_2);
  assign when_ArraySlice_l158_174 = (_zz_when_ArraySlice_l158_174 <= _zz_when_ArraySlice_l158_174_3);
  assign when_ArraySlice_l159_174 = (_zz_when_ArraySlice_l159_174 <= _zz_when_ArraySlice_l159_174_2);
  assign _zz_realValue_0_174 = (_zz__zz_realValue_0_174 % _zz__zz_realValue_0_174_1);
  assign when_ArraySlice_l110_174 = (_zz_realValue_0_174 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_174) begin
      realValue_0_174 = (_zz_realValue_0_174_1 - _zz_realValue_0_174);
    end else begin
      realValue_0_174 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_174 = (_zz_when_ArraySlice_l166_174 <= _zz_when_ArraySlice_l166_174_2);
  assign when_ArraySlice_l158_175 = (_zz_when_ArraySlice_l158_175 <= _zz_when_ArraySlice_l158_175_3);
  assign when_ArraySlice_l159_175 = (_zz_when_ArraySlice_l159_175 <= _zz_when_ArraySlice_l159_175_2);
  assign _zz_realValue_0_175 = (_zz__zz_realValue_0_175 % _zz__zz_realValue_0_175_1);
  assign when_ArraySlice_l110_175 = (_zz_realValue_0_175 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_175) begin
      realValue_0_175 = (_zz_realValue_0_175_1 - _zz_realValue_0_175);
    end else begin
      realValue_0_175 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_175 = (_zz_when_ArraySlice_l166_175 <= _zz_when_ArraySlice_l166_175_2);
  assign when_ArraySlice_l457_6 = (! ((((((_zz_when_ArraySlice_l457_6 && _zz_when_ArraySlice_l457_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l457_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_6_3 && _zz_when_ArraySlice_l457_6_4) && (debug_4_21 == _zz_when_ArraySlice_l457_6_5)) && (debug_5_21 == 1'b1)) && (debug_6_21 == 1'b1)) && (debug_7_21 == 1'b1))));
  assign outputStreamArrayData_6_fire_5 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l461_6 = ((_zz_when_ArraySlice_l461_6 == 13'h0) && outputStreamArrayData_6_fire_5);
  assign when_ArraySlice_l447_6 = (allowPadding_6 && (_zz_when_ArraySlice_l447_6 <= _zz_when_ArraySlice_l447_6_1));
  assign outputStreamArrayData_6_fire_6 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l468_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l468_6);
  assign when_ArraySlice_l376_7 = (_zz_when_ArraySlice_l376_7 < _zz_when_ArraySlice_l376_7_3);
  assign when_ArraySlice_l377_7 = ((! holdReadOp_7) && (_zz_when_ArraySlice_l377_7 != 7'h0));
  assign _zz_outputStreamArrayData_7_valid = (selectReadFifo_7 + _zz__zz_outputStreamArrayData_7_valid);
  assign _zz_10 = ({127'd0,1'b1} <<< _zz__zz_10);
  assign _zz_io_pop_ready_7 = outputStreamArrayData_7_ready;
  assign when_ArraySlice_l382_7 = (! holdReadOp_7);
  assign outputStreamArrayData_7_fire = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l383_7 = ((7'h01 < _zz_when_ArraySlice_l383_7) && outputStreamArrayData_7_fire);
  assign when_ArraySlice_l384_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l384_7);
  assign when_ArraySlice_l387_7 = (_zz_when_ArraySlice_l387_7 == 13'h0);
  assign outputStreamArrayData_7_fire_1 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l392_7 = ((_zz_when_ArraySlice_l392_7 == 7'h01) && outputStreamArrayData_7_fire_1);
  assign when_ArraySlice_l393_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l393_7);
  assign _zz_realValue1_0_21 = (_zz__zz_realValue1_0_21 % _zz__zz_realValue1_0_21_1);
  assign when_ArraySlice_l95_21 = (_zz_realValue1_0_21 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_21) begin
      realValue1_0_21 = (_zz_realValue1_0_21_1 - _zz_realValue1_0_21);
    end else begin
      realValue1_0_21 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l395_7 = (_zz_when_ArraySlice_l395_7 < _zz_when_ArraySlice_l395_7_2);
  always @(*) begin
    debug_0_22 = 1'b0;
    if(when_ArraySlice_l158_176) begin
      if(when_ArraySlice_l159_176) begin
        debug_0_22 = 1'b1;
      end else begin
        debug_0_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_176) begin
        debug_0_22 = 1'b1;
      end else begin
        debug_0_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_22 = 1'b0;
    if(when_ArraySlice_l158_177) begin
      if(when_ArraySlice_l159_177) begin
        debug_1_22 = 1'b1;
      end else begin
        debug_1_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_177) begin
        debug_1_22 = 1'b1;
      end else begin
        debug_1_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_22 = 1'b0;
    if(when_ArraySlice_l158_178) begin
      if(when_ArraySlice_l159_178) begin
        debug_2_22 = 1'b1;
      end else begin
        debug_2_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_178) begin
        debug_2_22 = 1'b1;
      end else begin
        debug_2_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_22 = 1'b0;
    if(when_ArraySlice_l158_179) begin
      if(when_ArraySlice_l159_179) begin
        debug_3_22 = 1'b1;
      end else begin
        debug_3_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_179) begin
        debug_3_22 = 1'b1;
      end else begin
        debug_3_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_22 = 1'b0;
    if(when_ArraySlice_l158_180) begin
      if(when_ArraySlice_l159_180) begin
        debug_4_22 = 1'b1;
      end else begin
        debug_4_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_180) begin
        debug_4_22 = 1'b1;
      end else begin
        debug_4_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_22 = 1'b0;
    if(when_ArraySlice_l158_181) begin
      if(when_ArraySlice_l159_181) begin
        debug_5_22 = 1'b1;
      end else begin
        debug_5_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_181) begin
        debug_5_22 = 1'b1;
      end else begin
        debug_5_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_22 = 1'b0;
    if(when_ArraySlice_l158_182) begin
      if(when_ArraySlice_l159_182) begin
        debug_6_22 = 1'b1;
      end else begin
        debug_6_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_182) begin
        debug_6_22 = 1'b1;
      end else begin
        debug_6_22 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_22 = 1'b0;
    if(when_ArraySlice_l158_183) begin
      if(when_ArraySlice_l159_183) begin
        debug_7_22 = 1'b1;
      end else begin
        debug_7_22 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_183) begin
        debug_7_22 = 1'b1;
      end else begin
        debug_7_22 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_176 = (_zz_when_ArraySlice_l158_176 <= _zz_when_ArraySlice_l158_176_3);
  assign when_ArraySlice_l159_176 = (_zz_when_ArraySlice_l159_176 <= _zz_when_ArraySlice_l159_176_1);
  assign _zz_realValue_0_176 = (_zz__zz_realValue_0_176 % _zz__zz_realValue_0_176_1);
  assign when_ArraySlice_l110_176 = (_zz_realValue_0_176 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_176) begin
      realValue_0_176 = (_zz_realValue_0_176_1 - _zz_realValue_0_176);
    end else begin
      realValue_0_176 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_176 = (_zz_when_ArraySlice_l166_176 <= _zz_when_ArraySlice_l166_176_1);
  assign when_ArraySlice_l158_177 = (_zz_when_ArraySlice_l158_177 <= _zz_when_ArraySlice_l158_177_3);
  assign when_ArraySlice_l159_177 = (_zz_when_ArraySlice_l159_177 <= _zz_when_ArraySlice_l159_177_2);
  assign _zz_realValue_0_177 = (_zz__zz_realValue_0_177 % _zz__zz_realValue_0_177_1);
  assign when_ArraySlice_l110_177 = (_zz_realValue_0_177 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_177) begin
      realValue_0_177 = (_zz_realValue_0_177_1 - _zz_realValue_0_177);
    end else begin
      realValue_0_177 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_177 = (_zz_when_ArraySlice_l166_177 <= _zz_when_ArraySlice_l166_177_2);
  assign when_ArraySlice_l158_178 = (_zz_when_ArraySlice_l158_178 <= _zz_when_ArraySlice_l158_178_3);
  assign when_ArraySlice_l159_178 = (_zz_when_ArraySlice_l159_178 <= _zz_when_ArraySlice_l159_178_2);
  assign _zz_realValue_0_178 = (_zz__zz_realValue_0_178 % _zz__zz_realValue_0_178_1);
  assign when_ArraySlice_l110_178 = (_zz_realValue_0_178 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_178) begin
      realValue_0_178 = (_zz_realValue_0_178_1 - _zz_realValue_0_178);
    end else begin
      realValue_0_178 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_178 = (_zz_when_ArraySlice_l166_178 <= _zz_when_ArraySlice_l166_178_2);
  assign when_ArraySlice_l158_179 = (_zz_when_ArraySlice_l158_179 <= _zz_when_ArraySlice_l158_179_3);
  assign when_ArraySlice_l159_179 = (_zz_when_ArraySlice_l159_179 <= _zz_when_ArraySlice_l159_179_2);
  assign _zz_realValue_0_179 = (_zz__zz_realValue_0_179 % _zz__zz_realValue_0_179_1);
  assign when_ArraySlice_l110_179 = (_zz_realValue_0_179 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_179) begin
      realValue_0_179 = (_zz_realValue_0_179_1 - _zz_realValue_0_179);
    end else begin
      realValue_0_179 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_179 = (_zz_when_ArraySlice_l166_179 <= _zz_when_ArraySlice_l166_179_2);
  assign when_ArraySlice_l158_180 = (_zz_when_ArraySlice_l158_180 <= _zz_when_ArraySlice_l158_180_3);
  assign when_ArraySlice_l159_180 = (_zz_when_ArraySlice_l159_180 <= _zz_when_ArraySlice_l159_180_2);
  assign _zz_realValue_0_180 = (_zz__zz_realValue_0_180 % _zz__zz_realValue_0_180_1);
  assign when_ArraySlice_l110_180 = (_zz_realValue_0_180 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_180) begin
      realValue_0_180 = (_zz_realValue_0_180_1 - _zz_realValue_0_180);
    end else begin
      realValue_0_180 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_180 = (_zz_when_ArraySlice_l166_180 <= _zz_when_ArraySlice_l166_180_2);
  assign when_ArraySlice_l158_181 = (_zz_when_ArraySlice_l158_181 <= _zz_when_ArraySlice_l158_181_3);
  assign when_ArraySlice_l159_181 = (_zz_when_ArraySlice_l159_181 <= _zz_when_ArraySlice_l159_181_2);
  assign _zz_realValue_0_181 = (_zz__zz_realValue_0_181 % _zz__zz_realValue_0_181_1);
  assign when_ArraySlice_l110_181 = (_zz_realValue_0_181 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_181) begin
      realValue_0_181 = (_zz_realValue_0_181_1 - _zz_realValue_0_181);
    end else begin
      realValue_0_181 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_181 = (_zz_when_ArraySlice_l166_181 <= _zz_when_ArraySlice_l166_181_2);
  assign when_ArraySlice_l158_182 = (_zz_when_ArraySlice_l158_182 <= _zz_when_ArraySlice_l158_182_3);
  assign when_ArraySlice_l159_182 = (_zz_when_ArraySlice_l159_182 <= _zz_when_ArraySlice_l159_182_2);
  assign _zz_realValue_0_182 = (_zz__zz_realValue_0_182 % _zz__zz_realValue_0_182_1);
  assign when_ArraySlice_l110_182 = (_zz_realValue_0_182 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_182) begin
      realValue_0_182 = (_zz_realValue_0_182_1 - _zz_realValue_0_182);
    end else begin
      realValue_0_182 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_182 = (_zz_when_ArraySlice_l166_182 <= _zz_when_ArraySlice_l166_182_2);
  assign when_ArraySlice_l158_183 = (_zz_when_ArraySlice_l158_183 <= _zz_when_ArraySlice_l158_183_3);
  assign when_ArraySlice_l159_183 = (_zz_when_ArraySlice_l159_183 <= _zz_when_ArraySlice_l159_183_2);
  assign _zz_realValue_0_183 = (_zz__zz_realValue_0_183 % _zz__zz_realValue_0_183_1);
  assign when_ArraySlice_l110_183 = (_zz_realValue_0_183 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_183) begin
      realValue_0_183 = (_zz_realValue_0_183_1 - _zz_realValue_0_183);
    end else begin
      realValue_0_183 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_183 = (_zz_when_ArraySlice_l166_183 <= _zz_when_ArraySlice_l166_183_2);
  assign when_ArraySlice_l400_7 = (! ((((((_zz_when_ArraySlice_l400_7_1 && _zz_when_ArraySlice_l400_7_2) && (holdReadOp_4 == _zz_when_ArraySlice_l400_7_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l400_7_4 && _zz_when_ArraySlice_l400_7_5) && (debug_4_22 == _zz_when_ArraySlice_l400_7_6)) && (debug_5_22 == 1'b1)) && (debug_6_22 == 1'b1)) && (debug_7_22 == 1'b1))));
  assign when_ArraySlice_l403_7 = (_zz_when_ArraySlice_l403_7_1 <= _zz_when_ArraySlice_l403_7_2);
  assign when_ArraySlice_l406_7 = (_zz_when_ArraySlice_l406_7 <= _zz_when_ArraySlice_l406_7_1);
  assign when_ArraySlice_l413_7 = (_zz_when_ArraySlice_l413_7 == 13'h0);
  assign when_ArraySlice_l417_7 = (_zz_when_ArraySlice_l417_7 == 7'h0);
  assign outputStreamArrayData_7_fire_2 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l418_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l418_7) && outputStreamArrayData_7_fire_2);
  assign _zz_realValue1_0_22 = (_zz__zz_realValue1_0_22 % _zz__zz_realValue1_0_22_1);
  assign when_ArraySlice_l95_22 = (_zz_realValue1_0_22 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_22) begin
      realValue1_0_22 = (_zz_realValue1_0_22_1 - _zz_realValue1_0_22);
    end else begin
      realValue1_0_22 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l420_7 = (_zz_when_ArraySlice_l420_7 < _zz_when_ArraySlice_l420_7_2);
  always @(*) begin
    debug_0_23 = 1'b0;
    if(when_ArraySlice_l158_184) begin
      if(when_ArraySlice_l159_184) begin
        debug_0_23 = 1'b1;
      end else begin
        debug_0_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_184) begin
        debug_0_23 = 1'b1;
      end else begin
        debug_0_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_23 = 1'b0;
    if(when_ArraySlice_l158_185) begin
      if(when_ArraySlice_l159_185) begin
        debug_1_23 = 1'b1;
      end else begin
        debug_1_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_185) begin
        debug_1_23 = 1'b1;
      end else begin
        debug_1_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_23 = 1'b0;
    if(when_ArraySlice_l158_186) begin
      if(when_ArraySlice_l159_186) begin
        debug_2_23 = 1'b1;
      end else begin
        debug_2_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_186) begin
        debug_2_23 = 1'b1;
      end else begin
        debug_2_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_23 = 1'b0;
    if(when_ArraySlice_l158_187) begin
      if(when_ArraySlice_l159_187) begin
        debug_3_23 = 1'b1;
      end else begin
        debug_3_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_187) begin
        debug_3_23 = 1'b1;
      end else begin
        debug_3_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_23 = 1'b0;
    if(when_ArraySlice_l158_188) begin
      if(when_ArraySlice_l159_188) begin
        debug_4_23 = 1'b1;
      end else begin
        debug_4_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_188) begin
        debug_4_23 = 1'b1;
      end else begin
        debug_4_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_23 = 1'b0;
    if(when_ArraySlice_l158_189) begin
      if(when_ArraySlice_l159_189) begin
        debug_5_23 = 1'b1;
      end else begin
        debug_5_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_189) begin
        debug_5_23 = 1'b1;
      end else begin
        debug_5_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_23 = 1'b0;
    if(when_ArraySlice_l158_190) begin
      if(when_ArraySlice_l159_190) begin
        debug_6_23 = 1'b1;
      end else begin
        debug_6_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_190) begin
        debug_6_23 = 1'b1;
      end else begin
        debug_6_23 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_23 = 1'b0;
    if(when_ArraySlice_l158_191) begin
      if(when_ArraySlice_l159_191) begin
        debug_7_23 = 1'b1;
      end else begin
        debug_7_23 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_191) begin
        debug_7_23 = 1'b1;
      end else begin
        debug_7_23 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_184 = (_zz_when_ArraySlice_l158_184 <= _zz_when_ArraySlice_l158_184_3);
  assign when_ArraySlice_l159_184 = (_zz_when_ArraySlice_l159_184 <= _zz_when_ArraySlice_l159_184_1);
  assign _zz_realValue_0_184 = (_zz__zz_realValue_0_184 % _zz__zz_realValue_0_184_1);
  assign when_ArraySlice_l110_184 = (_zz_realValue_0_184 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_184) begin
      realValue_0_184 = (_zz_realValue_0_184_1 - _zz_realValue_0_184);
    end else begin
      realValue_0_184 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_184 = (_zz_when_ArraySlice_l166_184 <= _zz_when_ArraySlice_l166_184_1);
  assign when_ArraySlice_l158_185 = (_zz_when_ArraySlice_l158_185 <= _zz_when_ArraySlice_l158_185_3);
  assign when_ArraySlice_l159_185 = (_zz_when_ArraySlice_l159_185 <= _zz_when_ArraySlice_l159_185_2);
  assign _zz_realValue_0_185 = (_zz__zz_realValue_0_185 % _zz__zz_realValue_0_185_1);
  assign when_ArraySlice_l110_185 = (_zz_realValue_0_185 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_185) begin
      realValue_0_185 = (_zz_realValue_0_185_1 - _zz_realValue_0_185);
    end else begin
      realValue_0_185 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_185 = (_zz_when_ArraySlice_l166_185 <= _zz_when_ArraySlice_l166_185_2);
  assign when_ArraySlice_l158_186 = (_zz_when_ArraySlice_l158_186 <= _zz_when_ArraySlice_l158_186_3);
  assign when_ArraySlice_l159_186 = (_zz_when_ArraySlice_l159_186 <= _zz_when_ArraySlice_l159_186_2);
  assign _zz_realValue_0_186 = (_zz__zz_realValue_0_186 % _zz__zz_realValue_0_186_1);
  assign when_ArraySlice_l110_186 = (_zz_realValue_0_186 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_186) begin
      realValue_0_186 = (_zz_realValue_0_186_1 - _zz_realValue_0_186);
    end else begin
      realValue_0_186 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_186 = (_zz_when_ArraySlice_l166_186 <= _zz_when_ArraySlice_l166_186_2);
  assign when_ArraySlice_l158_187 = (_zz_when_ArraySlice_l158_187 <= _zz_when_ArraySlice_l158_187_3);
  assign when_ArraySlice_l159_187 = (_zz_when_ArraySlice_l159_187 <= _zz_when_ArraySlice_l159_187_2);
  assign _zz_realValue_0_187 = (_zz__zz_realValue_0_187 % _zz__zz_realValue_0_187_1);
  assign when_ArraySlice_l110_187 = (_zz_realValue_0_187 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_187) begin
      realValue_0_187 = (_zz_realValue_0_187_1 - _zz_realValue_0_187);
    end else begin
      realValue_0_187 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_187 = (_zz_when_ArraySlice_l166_187 <= _zz_when_ArraySlice_l166_187_2);
  assign when_ArraySlice_l158_188 = (_zz_when_ArraySlice_l158_188 <= _zz_when_ArraySlice_l158_188_3);
  assign when_ArraySlice_l159_188 = (_zz_when_ArraySlice_l159_188 <= _zz_when_ArraySlice_l159_188_2);
  assign _zz_realValue_0_188 = (_zz__zz_realValue_0_188 % _zz__zz_realValue_0_188_1);
  assign when_ArraySlice_l110_188 = (_zz_realValue_0_188 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_188) begin
      realValue_0_188 = (_zz_realValue_0_188_1 - _zz_realValue_0_188);
    end else begin
      realValue_0_188 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_188 = (_zz_when_ArraySlice_l166_188 <= _zz_when_ArraySlice_l166_188_2);
  assign when_ArraySlice_l158_189 = (_zz_when_ArraySlice_l158_189 <= _zz_when_ArraySlice_l158_189_3);
  assign when_ArraySlice_l159_189 = (_zz_when_ArraySlice_l159_189 <= _zz_when_ArraySlice_l159_189_2);
  assign _zz_realValue_0_189 = (_zz__zz_realValue_0_189 % _zz__zz_realValue_0_189_1);
  assign when_ArraySlice_l110_189 = (_zz_realValue_0_189 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_189) begin
      realValue_0_189 = (_zz_realValue_0_189_1 - _zz_realValue_0_189);
    end else begin
      realValue_0_189 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_189 = (_zz_when_ArraySlice_l166_189 <= _zz_when_ArraySlice_l166_189_2);
  assign when_ArraySlice_l158_190 = (_zz_when_ArraySlice_l158_190 <= _zz_when_ArraySlice_l158_190_3);
  assign when_ArraySlice_l159_190 = (_zz_when_ArraySlice_l159_190 <= _zz_when_ArraySlice_l159_190_2);
  assign _zz_realValue_0_190 = (_zz__zz_realValue_0_190 % _zz__zz_realValue_0_190_1);
  assign when_ArraySlice_l110_190 = (_zz_realValue_0_190 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_190) begin
      realValue_0_190 = (_zz_realValue_0_190_1 - _zz_realValue_0_190);
    end else begin
      realValue_0_190 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_190 = (_zz_when_ArraySlice_l166_190 <= _zz_when_ArraySlice_l166_190_2);
  assign when_ArraySlice_l158_191 = (_zz_when_ArraySlice_l158_191 <= _zz_when_ArraySlice_l158_191_3);
  assign when_ArraySlice_l159_191 = (_zz_when_ArraySlice_l159_191 <= _zz_when_ArraySlice_l159_191_2);
  assign _zz_realValue_0_191 = (_zz__zz_realValue_0_191 % _zz__zz_realValue_0_191_1);
  assign when_ArraySlice_l110_191 = (_zz_realValue_0_191 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_191) begin
      realValue_0_191 = (_zz_realValue_0_191_1 - _zz_realValue_0_191);
    end else begin
      realValue_0_191 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_191 = (_zz_when_ArraySlice_l166_191 <= _zz_when_ArraySlice_l166_191_2);
  assign when_ArraySlice_l425_7 = (! ((((((_zz_when_ArraySlice_l425_7 && _zz_when_ArraySlice_l425_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l425_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l425_7_3 && _zz_when_ArraySlice_l425_7_4) && (debug_4_23 == _zz_when_ArraySlice_l425_7_5)) && (debug_5_23 == 1'b1)) && (debug_6_23 == 1'b1)) && (debug_7_23 == 1'b1))));
  assign when_ArraySlice_l428_7 = (_zz_when_ArraySlice_l428_7_1 <= _zz_when_ArraySlice_l428_7_2);
  assign when_ArraySlice_l431_7 = (_zz_when_ArraySlice_l431_7 <= _zz_when_ArraySlice_l431_7_1);
  assign outputStreamArrayData_7_fire_3 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l438_7 = ((_zz_when_ArraySlice_l438_7 == 13'h0) && outputStreamArrayData_7_fire_3);
  assign outputStreamArrayData_7_fire_4 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l449_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l449_7) && outputStreamArrayData_7_fire_4);
  assign _zz_realValue1_0_23 = (_zz__zz_realValue1_0_23 % _zz__zz_realValue1_0_23_1);
  assign when_ArraySlice_l95_23 = (_zz_realValue1_0_23 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_23) begin
      realValue1_0_23 = (_zz_realValue1_0_23_1 - _zz_realValue1_0_23);
    end else begin
      realValue1_0_23 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l450_7 = (_zz_when_ArraySlice_l450_7 < _zz_when_ArraySlice_l450_7_2);
  always @(*) begin
    debug_0_24 = 1'b0;
    if(when_ArraySlice_l158_192) begin
      if(when_ArraySlice_l159_192) begin
        debug_0_24 = 1'b1;
      end else begin
        debug_0_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_192) begin
        debug_0_24 = 1'b1;
      end else begin
        debug_0_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_24 = 1'b0;
    if(when_ArraySlice_l158_193) begin
      if(when_ArraySlice_l159_193) begin
        debug_1_24 = 1'b1;
      end else begin
        debug_1_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_193) begin
        debug_1_24 = 1'b1;
      end else begin
        debug_1_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_24 = 1'b0;
    if(when_ArraySlice_l158_194) begin
      if(when_ArraySlice_l159_194) begin
        debug_2_24 = 1'b1;
      end else begin
        debug_2_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_194) begin
        debug_2_24 = 1'b1;
      end else begin
        debug_2_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_24 = 1'b0;
    if(when_ArraySlice_l158_195) begin
      if(when_ArraySlice_l159_195) begin
        debug_3_24 = 1'b1;
      end else begin
        debug_3_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_195) begin
        debug_3_24 = 1'b1;
      end else begin
        debug_3_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_24 = 1'b0;
    if(when_ArraySlice_l158_196) begin
      if(when_ArraySlice_l159_196) begin
        debug_4_24 = 1'b1;
      end else begin
        debug_4_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_196) begin
        debug_4_24 = 1'b1;
      end else begin
        debug_4_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_24 = 1'b0;
    if(when_ArraySlice_l158_197) begin
      if(when_ArraySlice_l159_197) begin
        debug_5_24 = 1'b1;
      end else begin
        debug_5_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_197) begin
        debug_5_24 = 1'b1;
      end else begin
        debug_5_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_24 = 1'b0;
    if(when_ArraySlice_l158_198) begin
      if(when_ArraySlice_l159_198) begin
        debug_6_24 = 1'b1;
      end else begin
        debug_6_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_198) begin
        debug_6_24 = 1'b1;
      end else begin
        debug_6_24 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_24 = 1'b0;
    if(when_ArraySlice_l158_199) begin
      if(when_ArraySlice_l159_199) begin
        debug_7_24 = 1'b1;
      end else begin
        debug_7_24 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_199) begin
        debug_7_24 = 1'b1;
      end else begin
        debug_7_24 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_192 = (_zz_when_ArraySlice_l158_192 <= _zz_when_ArraySlice_l158_192_3);
  assign when_ArraySlice_l159_192 = (_zz_when_ArraySlice_l159_192 <= _zz_when_ArraySlice_l159_192_1);
  assign _zz_realValue_0_192 = (_zz__zz_realValue_0_192 % _zz__zz_realValue_0_192_1);
  assign when_ArraySlice_l110_192 = (_zz_realValue_0_192 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_192) begin
      realValue_0_192 = (_zz_realValue_0_192_1 - _zz_realValue_0_192);
    end else begin
      realValue_0_192 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_192 = (_zz_when_ArraySlice_l166_192 <= _zz_when_ArraySlice_l166_192_1);
  assign when_ArraySlice_l158_193 = (_zz_when_ArraySlice_l158_193 <= _zz_when_ArraySlice_l158_193_3);
  assign when_ArraySlice_l159_193 = (_zz_when_ArraySlice_l159_193 <= _zz_when_ArraySlice_l159_193_2);
  assign _zz_realValue_0_193 = (_zz__zz_realValue_0_193 % _zz__zz_realValue_0_193_1);
  assign when_ArraySlice_l110_193 = (_zz_realValue_0_193 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_193) begin
      realValue_0_193 = (_zz_realValue_0_193_1 - _zz_realValue_0_193);
    end else begin
      realValue_0_193 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_193 = (_zz_when_ArraySlice_l166_193 <= _zz_when_ArraySlice_l166_193_2);
  assign when_ArraySlice_l158_194 = (_zz_when_ArraySlice_l158_194 <= _zz_when_ArraySlice_l158_194_3);
  assign when_ArraySlice_l159_194 = (_zz_when_ArraySlice_l159_194 <= _zz_when_ArraySlice_l159_194_2);
  assign _zz_realValue_0_194 = (_zz__zz_realValue_0_194 % _zz__zz_realValue_0_194_1);
  assign when_ArraySlice_l110_194 = (_zz_realValue_0_194 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_194) begin
      realValue_0_194 = (_zz_realValue_0_194_1 - _zz_realValue_0_194);
    end else begin
      realValue_0_194 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_194 = (_zz_when_ArraySlice_l166_194 <= _zz_when_ArraySlice_l166_194_2);
  assign when_ArraySlice_l158_195 = (_zz_when_ArraySlice_l158_195 <= _zz_when_ArraySlice_l158_195_3);
  assign when_ArraySlice_l159_195 = (_zz_when_ArraySlice_l159_195 <= _zz_when_ArraySlice_l159_195_2);
  assign _zz_realValue_0_195 = (_zz__zz_realValue_0_195 % _zz__zz_realValue_0_195_1);
  assign when_ArraySlice_l110_195 = (_zz_realValue_0_195 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_195) begin
      realValue_0_195 = (_zz_realValue_0_195_1 - _zz_realValue_0_195);
    end else begin
      realValue_0_195 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_195 = (_zz_when_ArraySlice_l166_195 <= _zz_when_ArraySlice_l166_195_2);
  assign when_ArraySlice_l158_196 = (_zz_when_ArraySlice_l158_196 <= _zz_when_ArraySlice_l158_196_3);
  assign when_ArraySlice_l159_196 = (_zz_when_ArraySlice_l159_196 <= _zz_when_ArraySlice_l159_196_2);
  assign _zz_realValue_0_196 = (_zz__zz_realValue_0_196 % _zz__zz_realValue_0_196_1);
  assign when_ArraySlice_l110_196 = (_zz_realValue_0_196 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_196) begin
      realValue_0_196 = (_zz_realValue_0_196_1 - _zz_realValue_0_196);
    end else begin
      realValue_0_196 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_196 = (_zz_when_ArraySlice_l166_196 <= _zz_when_ArraySlice_l166_196_2);
  assign when_ArraySlice_l158_197 = (_zz_when_ArraySlice_l158_197 <= _zz_when_ArraySlice_l158_197_3);
  assign when_ArraySlice_l159_197 = (_zz_when_ArraySlice_l159_197 <= _zz_when_ArraySlice_l159_197_2);
  assign _zz_realValue_0_197 = (_zz__zz_realValue_0_197 % _zz__zz_realValue_0_197_1);
  assign when_ArraySlice_l110_197 = (_zz_realValue_0_197 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_197) begin
      realValue_0_197 = (_zz_realValue_0_197_1 - _zz_realValue_0_197);
    end else begin
      realValue_0_197 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_197 = (_zz_when_ArraySlice_l166_197 <= _zz_when_ArraySlice_l166_197_2);
  assign when_ArraySlice_l158_198 = (_zz_when_ArraySlice_l158_198 <= _zz_when_ArraySlice_l158_198_3);
  assign when_ArraySlice_l159_198 = (_zz_when_ArraySlice_l159_198 <= _zz_when_ArraySlice_l159_198_2);
  assign _zz_realValue_0_198 = (_zz__zz_realValue_0_198 % _zz__zz_realValue_0_198_1);
  assign when_ArraySlice_l110_198 = (_zz_realValue_0_198 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_198) begin
      realValue_0_198 = (_zz_realValue_0_198_1 - _zz_realValue_0_198);
    end else begin
      realValue_0_198 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_198 = (_zz_when_ArraySlice_l166_198 <= _zz_when_ArraySlice_l166_198_2);
  assign when_ArraySlice_l158_199 = (_zz_when_ArraySlice_l158_199 <= _zz_when_ArraySlice_l158_199_3);
  assign when_ArraySlice_l159_199 = (_zz_when_ArraySlice_l159_199 <= _zz_when_ArraySlice_l159_199_2);
  assign _zz_realValue_0_199 = (_zz__zz_realValue_0_199 % _zz__zz_realValue_0_199_1);
  assign when_ArraySlice_l110_199 = (_zz_realValue_0_199 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_199) begin
      realValue_0_199 = (_zz_realValue_0_199_1 - _zz_realValue_0_199);
    end else begin
      realValue_0_199 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_199 = (_zz_when_ArraySlice_l166_199 <= _zz_when_ArraySlice_l166_199_2);
  assign when_ArraySlice_l457_7 = (! ((((((_zz_when_ArraySlice_l457_7 && _zz_when_ArraySlice_l457_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l457_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l457_7_3 && _zz_when_ArraySlice_l457_7_4) && (debug_4_24 == _zz_when_ArraySlice_l457_7_5)) && (debug_5_24 == 1'b1)) && (debug_6_24 == 1'b1)) && (debug_7_24 == 1'b1))));
  assign outputStreamArrayData_7_fire_5 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l461_7 = ((_zz_when_ArraySlice_l461_7 == 13'h0) && outputStreamArrayData_7_fire_5);
  assign when_ArraySlice_l447_7 = (allowPadding_7 && (_zz_when_ArraySlice_l447_7 <= _zz_when_ArraySlice_l447_7_1));
  assign outputStreamArrayData_7_fire_6 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l468_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l468_7);
  always @(*) begin
    debug_0_25 = 1'b0;
    if(when_ArraySlice_l158_200) begin
      if(when_ArraySlice_l159_200) begin
        debug_0_25 = 1'b1;
      end else begin
        debug_0_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_200) begin
        debug_0_25 = 1'b1;
      end else begin
        debug_0_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_25 = 1'b0;
    if(when_ArraySlice_l158_201) begin
      if(when_ArraySlice_l159_201) begin
        debug_1_25 = 1'b1;
      end else begin
        debug_1_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_201) begin
        debug_1_25 = 1'b1;
      end else begin
        debug_1_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_25 = 1'b0;
    if(when_ArraySlice_l158_202) begin
      if(when_ArraySlice_l159_202) begin
        debug_2_25 = 1'b1;
      end else begin
        debug_2_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_202) begin
        debug_2_25 = 1'b1;
      end else begin
        debug_2_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_25 = 1'b0;
    if(when_ArraySlice_l158_203) begin
      if(when_ArraySlice_l159_203) begin
        debug_3_25 = 1'b1;
      end else begin
        debug_3_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_203) begin
        debug_3_25 = 1'b1;
      end else begin
        debug_3_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_25 = 1'b0;
    if(when_ArraySlice_l158_204) begin
      if(when_ArraySlice_l159_204) begin
        debug_4_25 = 1'b1;
      end else begin
        debug_4_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_204) begin
        debug_4_25 = 1'b1;
      end else begin
        debug_4_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_25 = 1'b0;
    if(when_ArraySlice_l158_205) begin
      if(when_ArraySlice_l159_205) begin
        debug_5_25 = 1'b1;
      end else begin
        debug_5_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_205) begin
        debug_5_25 = 1'b1;
      end else begin
        debug_5_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_25 = 1'b0;
    if(when_ArraySlice_l158_206) begin
      if(when_ArraySlice_l159_206) begin
        debug_6_25 = 1'b1;
      end else begin
        debug_6_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_206) begin
        debug_6_25 = 1'b1;
      end else begin
        debug_6_25 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_25 = 1'b0;
    if(when_ArraySlice_l158_207) begin
      if(when_ArraySlice_l159_207) begin
        debug_7_25 = 1'b1;
      end else begin
        debug_7_25 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_207) begin
        debug_7_25 = 1'b1;
      end else begin
        debug_7_25 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_200 = (_zz_when_ArraySlice_l158_200 <= _zz_when_ArraySlice_l158_200_3);
  assign when_ArraySlice_l159_200 = (_zz_when_ArraySlice_l159_200 <= _zz_when_ArraySlice_l159_200_1);
  assign _zz_realValue_0_200 = (_zz__zz_realValue_0_200 % _zz__zz_realValue_0_200_1);
  assign when_ArraySlice_l110_200 = (_zz_realValue_0_200 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_200) begin
      realValue_0_200 = (_zz_realValue_0_200_1 - _zz_realValue_0_200);
    end else begin
      realValue_0_200 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_200 = (_zz_when_ArraySlice_l166_200 <= _zz_when_ArraySlice_l166_200_1);
  assign when_ArraySlice_l158_201 = (_zz_when_ArraySlice_l158_201 <= _zz_when_ArraySlice_l158_201_3);
  assign when_ArraySlice_l159_201 = (_zz_when_ArraySlice_l159_201 <= _zz_when_ArraySlice_l159_201_2);
  assign _zz_realValue_0_201 = (_zz__zz_realValue_0_201 % _zz__zz_realValue_0_201_1);
  assign when_ArraySlice_l110_201 = (_zz_realValue_0_201 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_201) begin
      realValue_0_201 = (_zz_realValue_0_201_1 - _zz_realValue_0_201);
    end else begin
      realValue_0_201 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_201 = (_zz_when_ArraySlice_l166_201 <= _zz_when_ArraySlice_l166_201_2);
  assign when_ArraySlice_l158_202 = (_zz_when_ArraySlice_l158_202 <= _zz_when_ArraySlice_l158_202_3);
  assign when_ArraySlice_l159_202 = (_zz_when_ArraySlice_l159_202 <= _zz_when_ArraySlice_l159_202_2);
  assign _zz_realValue_0_202 = (_zz__zz_realValue_0_202 % _zz__zz_realValue_0_202_1);
  assign when_ArraySlice_l110_202 = (_zz_realValue_0_202 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_202) begin
      realValue_0_202 = (_zz_realValue_0_202_1 - _zz_realValue_0_202);
    end else begin
      realValue_0_202 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_202 = (_zz_when_ArraySlice_l166_202 <= _zz_when_ArraySlice_l166_202_2);
  assign when_ArraySlice_l158_203 = (_zz_when_ArraySlice_l158_203 <= _zz_when_ArraySlice_l158_203_3);
  assign when_ArraySlice_l159_203 = (_zz_when_ArraySlice_l159_203 <= _zz_when_ArraySlice_l159_203_2);
  assign _zz_realValue_0_203 = (_zz__zz_realValue_0_203 % _zz__zz_realValue_0_203_1);
  assign when_ArraySlice_l110_203 = (_zz_realValue_0_203 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_203) begin
      realValue_0_203 = (_zz_realValue_0_203_1 - _zz_realValue_0_203);
    end else begin
      realValue_0_203 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_203 = (_zz_when_ArraySlice_l166_203 <= _zz_when_ArraySlice_l166_203_2);
  assign when_ArraySlice_l158_204 = (_zz_when_ArraySlice_l158_204 <= _zz_when_ArraySlice_l158_204_3);
  assign when_ArraySlice_l159_204 = (_zz_when_ArraySlice_l159_204 <= _zz_when_ArraySlice_l159_204_2);
  assign _zz_realValue_0_204 = (_zz__zz_realValue_0_204 % _zz__zz_realValue_0_204_1);
  assign when_ArraySlice_l110_204 = (_zz_realValue_0_204 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_204) begin
      realValue_0_204 = (_zz_realValue_0_204_1 - _zz_realValue_0_204);
    end else begin
      realValue_0_204 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_204 = (_zz_when_ArraySlice_l166_204 <= _zz_when_ArraySlice_l166_204_2);
  assign when_ArraySlice_l158_205 = (_zz_when_ArraySlice_l158_205 <= _zz_when_ArraySlice_l158_205_3);
  assign when_ArraySlice_l159_205 = (_zz_when_ArraySlice_l159_205 <= _zz_when_ArraySlice_l159_205_2);
  assign _zz_realValue_0_205 = (_zz__zz_realValue_0_205 % _zz__zz_realValue_0_205_1);
  assign when_ArraySlice_l110_205 = (_zz_realValue_0_205 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_205) begin
      realValue_0_205 = (_zz_realValue_0_205_1 - _zz_realValue_0_205);
    end else begin
      realValue_0_205 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_205 = (_zz_when_ArraySlice_l166_205 <= _zz_when_ArraySlice_l166_205_2);
  assign when_ArraySlice_l158_206 = (_zz_when_ArraySlice_l158_206 <= _zz_when_ArraySlice_l158_206_3);
  assign when_ArraySlice_l159_206 = (_zz_when_ArraySlice_l159_206 <= _zz_when_ArraySlice_l159_206_2);
  assign _zz_realValue_0_206 = (_zz__zz_realValue_0_206 % _zz__zz_realValue_0_206_1);
  assign when_ArraySlice_l110_206 = (_zz_realValue_0_206 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_206) begin
      realValue_0_206 = (_zz_realValue_0_206_1 - _zz_realValue_0_206);
    end else begin
      realValue_0_206 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_206 = (_zz_when_ArraySlice_l166_206 <= _zz_when_ArraySlice_l166_206_2);
  assign when_ArraySlice_l158_207 = (_zz_when_ArraySlice_l158_207 <= _zz_when_ArraySlice_l158_207_3);
  assign when_ArraySlice_l159_207 = (_zz_when_ArraySlice_l159_207 <= _zz_when_ArraySlice_l159_207_2);
  assign _zz_realValue_0_207 = (_zz__zz_realValue_0_207 % _zz__zz_realValue_0_207_1);
  assign when_ArraySlice_l110_207 = (_zz_realValue_0_207 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_207) begin
      realValue_0_207 = (_zz_realValue_0_207_1 - _zz_realValue_0_207);
    end else begin
      realValue_0_207 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_207 = (_zz_when_ArraySlice_l166_207 <= _zz_when_ArraySlice_l166_207_2);
  assign when_ArraySlice_l478 = ((((((_zz_when_ArraySlice_l478 && _zz_when_ArraySlice_l478_1) && (holdReadOp_4 == _zz_when_ArraySlice_l478_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l478_3 && _zz_when_ArraySlice_l478_4) && (debug_4_25 == _zz_when_ArraySlice_l478_5)) && (debug_5_25 == 1'b1)) && (debug_6_25 == 1'b1)) && (debug_7_25 == 1'b1)));
  assign when_ArraySlice_l481 = (! allowPadding_0);
  assign when_ArraySlice_l481_1 = (! allowPadding_1);
  assign when_ArraySlice_l481_2 = (! allowPadding_2);
  assign when_ArraySlice_l481_3 = (! allowPadding_3);
  assign when_ArraySlice_l481_4 = (! allowPadding_4);
  assign when_ArraySlice_l481_5 = (! allowPadding_5);
  assign when_ArraySlice_l481_6 = (! allowPadding_6);
  assign when_ArraySlice_l481_7 = (! allowPadding_7);
  assign when_ArraySlice_l233 = (_zz_when_ArraySlice_l233 < _zz_when_ArraySlice_l233_3);
  assign when_ArraySlice_l234 = ((! holdReadOp_0) && (_zz_when_ArraySlice_l234 != 7'h0));
  assign _zz_outputStreamArrayData_0_valid_1 = (selectReadFifo_0 + _zz__zz_outputStreamArrayData_0_valid_1_1);
  assign _zz_11 = ({127'd0,1'b1} <<< _zz__zz_11);
  assign _zz_io_pop_ready_8 = outputStreamArrayData_0_ready;
  assign when_ArraySlice_l239 = (! holdReadOp_0);
  assign outputStreamArrayData_0_fire_7 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l240 = ((7'h01 < _zz_when_ArraySlice_l240) && outputStreamArrayData_0_fire_7);
  assign when_ArraySlice_l241 = (handshakeTimes_0_value == _zz_when_ArraySlice_l241);
  assign when_ArraySlice_l244 = (_zz_when_ArraySlice_l244 == 13'h0);
  assign outputStreamArrayData_0_fire_8 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l249 = ((_zz_when_ArraySlice_l249 == 7'h01) && outputStreamArrayData_0_fire_8);
  assign when_ArraySlice_l250 = (handshakeTimes_0_value == _zz_when_ArraySlice_l250);
  assign _zz_realValue1_0_24 = (_zz__zz_realValue1_0_24 % _zz__zz_realValue1_0_24_1);
  assign when_ArraySlice_l95_24 = (_zz_realValue1_0_24 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_24) begin
      realValue1_0_24 = (_zz_realValue1_0_24_1 - _zz_realValue1_0_24);
    end else begin
      realValue1_0_24 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252 = (_zz_when_ArraySlice_l252 < _zz_when_ArraySlice_l252_2);
  always @(*) begin
    debug_0_26 = 1'b0;
    if(when_ArraySlice_l158_208) begin
      if(when_ArraySlice_l159_208) begin
        debug_0_26 = 1'b1;
      end else begin
        debug_0_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_208) begin
        debug_0_26 = 1'b1;
      end else begin
        debug_0_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_26 = 1'b0;
    if(when_ArraySlice_l158_209) begin
      if(when_ArraySlice_l159_209) begin
        debug_1_26 = 1'b1;
      end else begin
        debug_1_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_209) begin
        debug_1_26 = 1'b1;
      end else begin
        debug_1_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_26 = 1'b0;
    if(when_ArraySlice_l158_210) begin
      if(when_ArraySlice_l159_210) begin
        debug_2_26 = 1'b1;
      end else begin
        debug_2_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_210) begin
        debug_2_26 = 1'b1;
      end else begin
        debug_2_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_26 = 1'b0;
    if(when_ArraySlice_l158_211) begin
      if(when_ArraySlice_l159_211) begin
        debug_3_26 = 1'b1;
      end else begin
        debug_3_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_211) begin
        debug_3_26 = 1'b1;
      end else begin
        debug_3_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_26 = 1'b0;
    if(when_ArraySlice_l158_212) begin
      if(when_ArraySlice_l159_212) begin
        debug_4_26 = 1'b1;
      end else begin
        debug_4_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_212) begin
        debug_4_26 = 1'b1;
      end else begin
        debug_4_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_26 = 1'b0;
    if(when_ArraySlice_l158_213) begin
      if(when_ArraySlice_l159_213) begin
        debug_5_26 = 1'b1;
      end else begin
        debug_5_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_213) begin
        debug_5_26 = 1'b1;
      end else begin
        debug_5_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_26 = 1'b0;
    if(when_ArraySlice_l158_214) begin
      if(when_ArraySlice_l159_214) begin
        debug_6_26 = 1'b1;
      end else begin
        debug_6_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_214) begin
        debug_6_26 = 1'b1;
      end else begin
        debug_6_26 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_26 = 1'b0;
    if(when_ArraySlice_l158_215) begin
      if(when_ArraySlice_l159_215) begin
        debug_7_26 = 1'b1;
      end else begin
        debug_7_26 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_215) begin
        debug_7_26 = 1'b1;
      end else begin
        debug_7_26 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_208 = (_zz_when_ArraySlice_l158_208 <= _zz_when_ArraySlice_l158_208_3);
  assign when_ArraySlice_l159_208 = (_zz_when_ArraySlice_l159_208 <= _zz_when_ArraySlice_l159_208_1);
  assign _zz_realValue_0_208 = (_zz__zz_realValue_0_208 % _zz__zz_realValue_0_208_1);
  assign when_ArraySlice_l110_208 = (_zz_realValue_0_208 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_208) begin
      realValue_0_208 = (_zz_realValue_0_208_1 - _zz_realValue_0_208);
    end else begin
      realValue_0_208 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_208 = (_zz_when_ArraySlice_l166_208 <= _zz_when_ArraySlice_l166_208_1);
  assign when_ArraySlice_l158_209 = (_zz_when_ArraySlice_l158_209 <= _zz_when_ArraySlice_l158_209_3);
  assign when_ArraySlice_l159_209 = (_zz_when_ArraySlice_l159_209 <= _zz_when_ArraySlice_l159_209_2);
  assign _zz_realValue_0_209 = (_zz__zz_realValue_0_209 % _zz__zz_realValue_0_209_1);
  assign when_ArraySlice_l110_209 = (_zz_realValue_0_209 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_209) begin
      realValue_0_209 = (_zz_realValue_0_209_1 - _zz_realValue_0_209);
    end else begin
      realValue_0_209 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_209 = (_zz_when_ArraySlice_l166_209 <= _zz_when_ArraySlice_l166_209_2);
  assign when_ArraySlice_l158_210 = (_zz_when_ArraySlice_l158_210 <= _zz_when_ArraySlice_l158_210_3);
  assign when_ArraySlice_l159_210 = (_zz_when_ArraySlice_l159_210 <= _zz_when_ArraySlice_l159_210_2);
  assign _zz_realValue_0_210 = (_zz__zz_realValue_0_210 % _zz__zz_realValue_0_210_1);
  assign when_ArraySlice_l110_210 = (_zz_realValue_0_210 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_210) begin
      realValue_0_210 = (_zz_realValue_0_210_1 - _zz_realValue_0_210);
    end else begin
      realValue_0_210 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_210 = (_zz_when_ArraySlice_l166_210 <= _zz_when_ArraySlice_l166_210_2);
  assign when_ArraySlice_l158_211 = (_zz_when_ArraySlice_l158_211 <= _zz_when_ArraySlice_l158_211_3);
  assign when_ArraySlice_l159_211 = (_zz_when_ArraySlice_l159_211 <= _zz_when_ArraySlice_l159_211_2);
  assign _zz_realValue_0_211 = (_zz__zz_realValue_0_211 % _zz__zz_realValue_0_211_1);
  assign when_ArraySlice_l110_211 = (_zz_realValue_0_211 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_211) begin
      realValue_0_211 = (_zz_realValue_0_211_1 - _zz_realValue_0_211);
    end else begin
      realValue_0_211 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_211 = (_zz_when_ArraySlice_l166_211 <= _zz_when_ArraySlice_l166_211_2);
  assign when_ArraySlice_l158_212 = (_zz_when_ArraySlice_l158_212 <= _zz_when_ArraySlice_l158_212_3);
  assign when_ArraySlice_l159_212 = (_zz_when_ArraySlice_l159_212 <= _zz_when_ArraySlice_l159_212_2);
  assign _zz_realValue_0_212 = (_zz__zz_realValue_0_212 % _zz__zz_realValue_0_212_1);
  assign when_ArraySlice_l110_212 = (_zz_realValue_0_212 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_212) begin
      realValue_0_212 = (_zz_realValue_0_212_1 - _zz_realValue_0_212);
    end else begin
      realValue_0_212 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_212 = (_zz_when_ArraySlice_l166_212 <= _zz_when_ArraySlice_l166_212_2);
  assign when_ArraySlice_l158_213 = (_zz_when_ArraySlice_l158_213 <= _zz_when_ArraySlice_l158_213_3);
  assign when_ArraySlice_l159_213 = (_zz_when_ArraySlice_l159_213 <= _zz_when_ArraySlice_l159_213_2);
  assign _zz_realValue_0_213 = (_zz__zz_realValue_0_213 % _zz__zz_realValue_0_213_1);
  assign when_ArraySlice_l110_213 = (_zz_realValue_0_213 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_213) begin
      realValue_0_213 = (_zz_realValue_0_213_1 - _zz_realValue_0_213);
    end else begin
      realValue_0_213 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_213 = (_zz_when_ArraySlice_l166_213 <= _zz_when_ArraySlice_l166_213_2);
  assign when_ArraySlice_l158_214 = (_zz_when_ArraySlice_l158_214 <= _zz_when_ArraySlice_l158_214_3);
  assign when_ArraySlice_l159_214 = (_zz_when_ArraySlice_l159_214 <= _zz_when_ArraySlice_l159_214_2);
  assign _zz_realValue_0_214 = (_zz__zz_realValue_0_214 % _zz__zz_realValue_0_214_1);
  assign when_ArraySlice_l110_214 = (_zz_realValue_0_214 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_214) begin
      realValue_0_214 = (_zz_realValue_0_214_1 - _zz_realValue_0_214);
    end else begin
      realValue_0_214 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_214 = (_zz_when_ArraySlice_l166_214 <= _zz_when_ArraySlice_l166_214_2);
  assign when_ArraySlice_l158_215 = (_zz_when_ArraySlice_l158_215 <= _zz_when_ArraySlice_l158_215_3);
  assign when_ArraySlice_l159_215 = (_zz_when_ArraySlice_l159_215 <= _zz_when_ArraySlice_l159_215_2);
  assign _zz_realValue_0_215 = (_zz__zz_realValue_0_215 % _zz__zz_realValue_0_215_1);
  assign when_ArraySlice_l110_215 = (_zz_realValue_0_215 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_215) begin
      realValue_0_215 = (_zz_realValue_0_215_1 - _zz_realValue_0_215);
    end else begin
      realValue_0_215 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_215 = (_zz_when_ArraySlice_l166_215 <= _zz_when_ArraySlice_l166_215_2);
  assign when_ArraySlice_l257 = (! ((((((_zz_when_ArraySlice_l257 && _zz_when_ArraySlice_l257_1) && (holdReadOp_4 == _zz_when_ArraySlice_l257_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_3 && _zz_when_ArraySlice_l257_4) && (debug_4_26 == _zz_when_ArraySlice_l257_5)) && (debug_5_26 == 1'b1)) && (debug_6_26 == 1'b1)) && (debug_7_26 == 1'b1))));
  assign when_ArraySlice_l260 = (_zz_when_ArraySlice_l260 <= _zz_when_ArraySlice_l260_1);
  assign when_ArraySlice_l263 = (_zz_when_ArraySlice_l263 <= _zz_when_ArraySlice_l263_1);
  assign when_ArraySlice_l270 = (_zz_when_ArraySlice_l270 == 13'h0);
  assign when_ArraySlice_l274 = (_zz_when_ArraySlice_l274 == 7'h0);
  assign outputStreamArrayData_0_fire_9 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l275 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l275) && outputStreamArrayData_0_fire_9);
  assign _zz_realValue1_0_25 = (_zz__zz_realValue1_0_25 % _zz__zz_realValue1_0_25_1);
  assign when_ArraySlice_l95_25 = (_zz_realValue1_0_25 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_25) begin
      realValue1_0_25 = (_zz_realValue1_0_25_1 - _zz_realValue1_0_25);
    end else begin
      realValue1_0_25 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277 = (_zz_when_ArraySlice_l277 < _zz_when_ArraySlice_l277_2);
  always @(*) begin
    debug_0_27 = 1'b0;
    if(when_ArraySlice_l158_216) begin
      if(when_ArraySlice_l159_216) begin
        debug_0_27 = 1'b1;
      end else begin
        debug_0_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_216) begin
        debug_0_27 = 1'b1;
      end else begin
        debug_0_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_27 = 1'b0;
    if(when_ArraySlice_l158_217) begin
      if(when_ArraySlice_l159_217) begin
        debug_1_27 = 1'b1;
      end else begin
        debug_1_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_217) begin
        debug_1_27 = 1'b1;
      end else begin
        debug_1_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_27 = 1'b0;
    if(when_ArraySlice_l158_218) begin
      if(when_ArraySlice_l159_218) begin
        debug_2_27 = 1'b1;
      end else begin
        debug_2_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_218) begin
        debug_2_27 = 1'b1;
      end else begin
        debug_2_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_27 = 1'b0;
    if(when_ArraySlice_l158_219) begin
      if(when_ArraySlice_l159_219) begin
        debug_3_27 = 1'b1;
      end else begin
        debug_3_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_219) begin
        debug_3_27 = 1'b1;
      end else begin
        debug_3_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_27 = 1'b0;
    if(when_ArraySlice_l158_220) begin
      if(when_ArraySlice_l159_220) begin
        debug_4_27 = 1'b1;
      end else begin
        debug_4_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_220) begin
        debug_4_27 = 1'b1;
      end else begin
        debug_4_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_27 = 1'b0;
    if(when_ArraySlice_l158_221) begin
      if(when_ArraySlice_l159_221) begin
        debug_5_27 = 1'b1;
      end else begin
        debug_5_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_221) begin
        debug_5_27 = 1'b1;
      end else begin
        debug_5_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_27 = 1'b0;
    if(when_ArraySlice_l158_222) begin
      if(when_ArraySlice_l159_222) begin
        debug_6_27 = 1'b1;
      end else begin
        debug_6_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_222) begin
        debug_6_27 = 1'b1;
      end else begin
        debug_6_27 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_27 = 1'b0;
    if(when_ArraySlice_l158_223) begin
      if(when_ArraySlice_l159_223) begin
        debug_7_27 = 1'b1;
      end else begin
        debug_7_27 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_223) begin
        debug_7_27 = 1'b1;
      end else begin
        debug_7_27 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_216 = (_zz_when_ArraySlice_l158_216 <= _zz_when_ArraySlice_l158_216_3);
  assign when_ArraySlice_l159_216 = (_zz_when_ArraySlice_l159_216 <= _zz_when_ArraySlice_l159_216_1);
  assign _zz_realValue_0_216 = (_zz__zz_realValue_0_216 % _zz__zz_realValue_0_216_1);
  assign when_ArraySlice_l110_216 = (_zz_realValue_0_216 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_216) begin
      realValue_0_216 = (_zz_realValue_0_216_1 - _zz_realValue_0_216);
    end else begin
      realValue_0_216 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_216 = (_zz_when_ArraySlice_l166_216 <= _zz_when_ArraySlice_l166_216_1);
  assign when_ArraySlice_l158_217 = (_zz_when_ArraySlice_l158_217 <= _zz_when_ArraySlice_l158_217_3);
  assign when_ArraySlice_l159_217 = (_zz_when_ArraySlice_l159_217 <= _zz_when_ArraySlice_l159_217_2);
  assign _zz_realValue_0_217 = (_zz__zz_realValue_0_217 % _zz__zz_realValue_0_217_1);
  assign when_ArraySlice_l110_217 = (_zz_realValue_0_217 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_217) begin
      realValue_0_217 = (_zz_realValue_0_217_1 - _zz_realValue_0_217);
    end else begin
      realValue_0_217 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_217 = (_zz_when_ArraySlice_l166_217 <= _zz_when_ArraySlice_l166_217_2);
  assign when_ArraySlice_l158_218 = (_zz_when_ArraySlice_l158_218 <= _zz_when_ArraySlice_l158_218_3);
  assign when_ArraySlice_l159_218 = (_zz_when_ArraySlice_l159_218 <= _zz_when_ArraySlice_l159_218_2);
  assign _zz_realValue_0_218 = (_zz__zz_realValue_0_218 % _zz__zz_realValue_0_218_1);
  assign when_ArraySlice_l110_218 = (_zz_realValue_0_218 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_218) begin
      realValue_0_218 = (_zz_realValue_0_218_1 - _zz_realValue_0_218);
    end else begin
      realValue_0_218 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_218 = (_zz_when_ArraySlice_l166_218 <= _zz_when_ArraySlice_l166_218_2);
  assign when_ArraySlice_l158_219 = (_zz_when_ArraySlice_l158_219 <= _zz_when_ArraySlice_l158_219_3);
  assign when_ArraySlice_l159_219 = (_zz_when_ArraySlice_l159_219 <= _zz_when_ArraySlice_l159_219_2);
  assign _zz_realValue_0_219 = (_zz__zz_realValue_0_219 % _zz__zz_realValue_0_219_1);
  assign when_ArraySlice_l110_219 = (_zz_realValue_0_219 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_219) begin
      realValue_0_219 = (_zz_realValue_0_219_1 - _zz_realValue_0_219);
    end else begin
      realValue_0_219 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_219 = (_zz_when_ArraySlice_l166_219 <= _zz_when_ArraySlice_l166_219_2);
  assign when_ArraySlice_l158_220 = (_zz_when_ArraySlice_l158_220 <= _zz_when_ArraySlice_l158_220_3);
  assign when_ArraySlice_l159_220 = (_zz_when_ArraySlice_l159_220 <= _zz_when_ArraySlice_l159_220_2);
  assign _zz_realValue_0_220 = (_zz__zz_realValue_0_220 % _zz__zz_realValue_0_220_1);
  assign when_ArraySlice_l110_220 = (_zz_realValue_0_220 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_220) begin
      realValue_0_220 = (_zz_realValue_0_220_1 - _zz_realValue_0_220);
    end else begin
      realValue_0_220 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_220 = (_zz_when_ArraySlice_l166_220 <= _zz_when_ArraySlice_l166_220_2);
  assign when_ArraySlice_l158_221 = (_zz_when_ArraySlice_l158_221 <= _zz_when_ArraySlice_l158_221_3);
  assign when_ArraySlice_l159_221 = (_zz_when_ArraySlice_l159_221 <= _zz_when_ArraySlice_l159_221_2);
  assign _zz_realValue_0_221 = (_zz__zz_realValue_0_221 % _zz__zz_realValue_0_221_1);
  assign when_ArraySlice_l110_221 = (_zz_realValue_0_221 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_221) begin
      realValue_0_221 = (_zz_realValue_0_221_1 - _zz_realValue_0_221);
    end else begin
      realValue_0_221 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_221 = (_zz_when_ArraySlice_l166_221 <= _zz_when_ArraySlice_l166_221_2);
  assign when_ArraySlice_l158_222 = (_zz_when_ArraySlice_l158_222 <= _zz_when_ArraySlice_l158_222_3);
  assign when_ArraySlice_l159_222 = (_zz_when_ArraySlice_l159_222 <= _zz_when_ArraySlice_l159_222_2);
  assign _zz_realValue_0_222 = (_zz__zz_realValue_0_222 % _zz__zz_realValue_0_222_1);
  assign when_ArraySlice_l110_222 = (_zz_realValue_0_222 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_222) begin
      realValue_0_222 = (_zz_realValue_0_222_1 - _zz_realValue_0_222);
    end else begin
      realValue_0_222 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_222 = (_zz_when_ArraySlice_l166_222 <= _zz_when_ArraySlice_l166_222_2);
  assign when_ArraySlice_l158_223 = (_zz_when_ArraySlice_l158_223 <= _zz_when_ArraySlice_l158_223_3);
  assign when_ArraySlice_l159_223 = (_zz_when_ArraySlice_l159_223 <= _zz_when_ArraySlice_l159_223_2);
  assign _zz_realValue_0_223 = (_zz__zz_realValue_0_223 % _zz__zz_realValue_0_223_1);
  assign when_ArraySlice_l110_223 = (_zz_realValue_0_223 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_223) begin
      realValue_0_223 = (_zz_realValue_0_223_1 - _zz_realValue_0_223);
    end else begin
      realValue_0_223 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_223 = (_zz_when_ArraySlice_l166_223 <= _zz_when_ArraySlice_l166_223_2);
  assign when_ArraySlice_l282 = (! ((((((_zz_when_ArraySlice_l282 && _zz_when_ArraySlice_l282_1) && (holdReadOp_4 == _zz_when_ArraySlice_l282_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_3 && _zz_when_ArraySlice_l282_4) && (debug_4_27 == _zz_when_ArraySlice_l282_5)) && (debug_5_27 == 1'b1)) && (debug_6_27 == 1'b1)) && (debug_7_27 == 1'b1))));
  assign when_ArraySlice_l285 = (_zz_when_ArraySlice_l285 <= _zz_when_ArraySlice_l285_1);
  assign when_ArraySlice_l288 = (_zz_when_ArraySlice_l288 <= _zz_when_ArraySlice_l288_1);
  assign outputStreamArrayData_0_fire_10 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l295 = ((_zz_when_ArraySlice_l295 == 13'h0) && outputStreamArrayData_0_fire_10);
  assign outputStreamArrayData_0_fire_11 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l306 = ((handshakeTimes_0_value == _zz_when_ArraySlice_l306) && outputStreamArrayData_0_fire_11);
  assign _zz_realValue1_0_26 = (_zz__zz_realValue1_0_26 % _zz__zz_realValue1_0_26_1);
  assign when_ArraySlice_l95_26 = (_zz_realValue1_0_26 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_26) begin
      realValue1_0_26 = (_zz_realValue1_0_26_1 - _zz_realValue1_0_26);
    end else begin
      realValue1_0_26 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307 = (_zz_when_ArraySlice_l307 < _zz_when_ArraySlice_l307_2);
  always @(*) begin
    debug_0_28 = 1'b0;
    if(when_ArraySlice_l158_224) begin
      if(when_ArraySlice_l159_224) begin
        debug_0_28 = 1'b1;
      end else begin
        debug_0_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_224) begin
        debug_0_28 = 1'b1;
      end else begin
        debug_0_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_28 = 1'b0;
    if(when_ArraySlice_l158_225) begin
      if(when_ArraySlice_l159_225) begin
        debug_1_28 = 1'b1;
      end else begin
        debug_1_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_225) begin
        debug_1_28 = 1'b1;
      end else begin
        debug_1_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_28 = 1'b0;
    if(when_ArraySlice_l158_226) begin
      if(when_ArraySlice_l159_226) begin
        debug_2_28 = 1'b1;
      end else begin
        debug_2_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_226) begin
        debug_2_28 = 1'b1;
      end else begin
        debug_2_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_28 = 1'b0;
    if(when_ArraySlice_l158_227) begin
      if(when_ArraySlice_l159_227) begin
        debug_3_28 = 1'b1;
      end else begin
        debug_3_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_227) begin
        debug_3_28 = 1'b1;
      end else begin
        debug_3_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_28 = 1'b0;
    if(when_ArraySlice_l158_228) begin
      if(when_ArraySlice_l159_228) begin
        debug_4_28 = 1'b1;
      end else begin
        debug_4_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_228) begin
        debug_4_28 = 1'b1;
      end else begin
        debug_4_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_28 = 1'b0;
    if(when_ArraySlice_l158_229) begin
      if(when_ArraySlice_l159_229) begin
        debug_5_28 = 1'b1;
      end else begin
        debug_5_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_229) begin
        debug_5_28 = 1'b1;
      end else begin
        debug_5_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_28 = 1'b0;
    if(when_ArraySlice_l158_230) begin
      if(when_ArraySlice_l159_230) begin
        debug_6_28 = 1'b1;
      end else begin
        debug_6_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_230) begin
        debug_6_28 = 1'b1;
      end else begin
        debug_6_28 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_28 = 1'b0;
    if(when_ArraySlice_l158_231) begin
      if(when_ArraySlice_l159_231) begin
        debug_7_28 = 1'b1;
      end else begin
        debug_7_28 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_231) begin
        debug_7_28 = 1'b1;
      end else begin
        debug_7_28 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_224 = (_zz_when_ArraySlice_l158_224 <= _zz_when_ArraySlice_l158_224_3);
  assign when_ArraySlice_l159_224 = (_zz_when_ArraySlice_l159_224 <= _zz_when_ArraySlice_l159_224_1);
  assign _zz_realValue_0_224 = (_zz__zz_realValue_0_224 % _zz__zz_realValue_0_224_1);
  assign when_ArraySlice_l110_224 = (_zz_realValue_0_224 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_224) begin
      realValue_0_224 = (_zz_realValue_0_224_1 - _zz_realValue_0_224);
    end else begin
      realValue_0_224 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_224 = (_zz_when_ArraySlice_l166_224 <= _zz_when_ArraySlice_l166_224_1);
  assign when_ArraySlice_l158_225 = (_zz_when_ArraySlice_l158_225 <= _zz_when_ArraySlice_l158_225_3);
  assign when_ArraySlice_l159_225 = (_zz_when_ArraySlice_l159_225 <= _zz_when_ArraySlice_l159_225_2);
  assign _zz_realValue_0_225 = (_zz__zz_realValue_0_225 % _zz__zz_realValue_0_225_1);
  assign when_ArraySlice_l110_225 = (_zz_realValue_0_225 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_225) begin
      realValue_0_225 = (_zz_realValue_0_225_1 - _zz_realValue_0_225);
    end else begin
      realValue_0_225 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_225 = (_zz_when_ArraySlice_l166_225 <= _zz_when_ArraySlice_l166_225_2);
  assign when_ArraySlice_l158_226 = (_zz_when_ArraySlice_l158_226 <= _zz_when_ArraySlice_l158_226_3);
  assign when_ArraySlice_l159_226 = (_zz_when_ArraySlice_l159_226 <= _zz_when_ArraySlice_l159_226_2);
  assign _zz_realValue_0_226 = (_zz__zz_realValue_0_226 % _zz__zz_realValue_0_226_1);
  assign when_ArraySlice_l110_226 = (_zz_realValue_0_226 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_226) begin
      realValue_0_226 = (_zz_realValue_0_226_1 - _zz_realValue_0_226);
    end else begin
      realValue_0_226 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_226 = (_zz_when_ArraySlice_l166_226 <= _zz_when_ArraySlice_l166_226_2);
  assign when_ArraySlice_l158_227 = (_zz_when_ArraySlice_l158_227 <= _zz_when_ArraySlice_l158_227_3);
  assign when_ArraySlice_l159_227 = (_zz_when_ArraySlice_l159_227 <= _zz_when_ArraySlice_l159_227_2);
  assign _zz_realValue_0_227 = (_zz__zz_realValue_0_227 % _zz__zz_realValue_0_227_1);
  assign when_ArraySlice_l110_227 = (_zz_realValue_0_227 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_227) begin
      realValue_0_227 = (_zz_realValue_0_227_1 - _zz_realValue_0_227);
    end else begin
      realValue_0_227 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_227 = (_zz_when_ArraySlice_l166_227 <= _zz_when_ArraySlice_l166_227_2);
  assign when_ArraySlice_l158_228 = (_zz_when_ArraySlice_l158_228 <= _zz_when_ArraySlice_l158_228_3);
  assign when_ArraySlice_l159_228 = (_zz_when_ArraySlice_l159_228 <= _zz_when_ArraySlice_l159_228_2);
  assign _zz_realValue_0_228 = (_zz__zz_realValue_0_228 % _zz__zz_realValue_0_228_1);
  assign when_ArraySlice_l110_228 = (_zz_realValue_0_228 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_228) begin
      realValue_0_228 = (_zz_realValue_0_228_1 - _zz_realValue_0_228);
    end else begin
      realValue_0_228 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_228 = (_zz_when_ArraySlice_l166_228 <= _zz_when_ArraySlice_l166_228_2);
  assign when_ArraySlice_l158_229 = (_zz_when_ArraySlice_l158_229 <= _zz_when_ArraySlice_l158_229_3);
  assign when_ArraySlice_l159_229 = (_zz_when_ArraySlice_l159_229 <= _zz_when_ArraySlice_l159_229_2);
  assign _zz_realValue_0_229 = (_zz__zz_realValue_0_229 % _zz__zz_realValue_0_229_1);
  assign when_ArraySlice_l110_229 = (_zz_realValue_0_229 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_229) begin
      realValue_0_229 = (_zz_realValue_0_229_1 - _zz_realValue_0_229);
    end else begin
      realValue_0_229 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_229 = (_zz_when_ArraySlice_l166_229 <= _zz_when_ArraySlice_l166_229_2);
  assign when_ArraySlice_l158_230 = (_zz_when_ArraySlice_l158_230 <= _zz_when_ArraySlice_l158_230_3);
  assign when_ArraySlice_l159_230 = (_zz_when_ArraySlice_l159_230 <= _zz_when_ArraySlice_l159_230_2);
  assign _zz_realValue_0_230 = (_zz__zz_realValue_0_230 % _zz__zz_realValue_0_230_1);
  assign when_ArraySlice_l110_230 = (_zz_realValue_0_230 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_230) begin
      realValue_0_230 = (_zz_realValue_0_230_1 - _zz_realValue_0_230);
    end else begin
      realValue_0_230 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_230 = (_zz_when_ArraySlice_l166_230 <= _zz_when_ArraySlice_l166_230_2);
  assign when_ArraySlice_l158_231 = (_zz_when_ArraySlice_l158_231 <= _zz_when_ArraySlice_l158_231_3);
  assign when_ArraySlice_l159_231 = (_zz_when_ArraySlice_l159_231 <= _zz_when_ArraySlice_l159_231_2);
  assign _zz_realValue_0_231 = (_zz__zz_realValue_0_231 % _zz__zz_realValue_0_231_1);
  assign when_ArraySlice_l110_231 = (_zz_realValue_0_231 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_231) begin
      realValue_0_231 = (_zz_realValue_0_231_1 - _zz_realValue_0_231);
    end else begin
      realValue_0_231 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_231 = (_zz_when_ArraySlice_l166_231 <= _zz_when_ArraySlice_l166_231_2);
  assign when_ArraySlice_l314 = (! ((((((_zz_when_ArraySlice_l314 && _zz_when_ArraySlice_l314_1) && (holdReadOp_4 == _zz_when_ArraySlice_l314_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_3 && _zz_when_ArraySlice_l314_4) && (debug_4_28 == _zz_when_ArraySlice_l314_5)) && (debug_5_28 == 1'b1)) && (debug_6_28 == 1'b1)) && (debug_7_28 == 1'b1))));
  assign outputStreamArrayData_0_fire_12 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l318 = ((_zz_when_ArraySlice_l318 == 13'h0) && outputStreamArrayData_0_fire_12);
  assign when_ArraySlice_l304 = (allowPadding_0 && (_zz_when_ArraySlice_l304 <= _zz_when_ArraySlice_l304_1));
  assign outputStreamArrayData_0_fire_13 = (outputStreamArrayData_0_valid && outputStreamArrayData_0_ready);
  assign when_ArraySlice_l325 = (handshakeTimes_0_value == _zz_when_ArraySlice_l325);
  assign when_ArraySlice_l233_1 = (_zz_when_ArraySlice_l233_1_1 < _zz_when_ArraySlice_l233_1_4);
  assign when_ArraySlice_l234_1 = ((! holdReadOp_1) && (_zz_when_ArraySlice_l234_1_1 != 7'h0));
  assign _zz_outputStreamArrayData_1_valid_1 = (selectReadFifo_1 + _zz__zz_outputStreamArrayData_1_valid_1_1);
  assign _zz_12 = ({127'd0,1'b1} <<< _zz__zz_12);
  assign _zz_io_pop_ready_9 = outputStreamArrayData_1_ready;
  assign when_ArraySlice_l239_1 = (! holdReadOp_1);
  assign outputStreamArrayData_1_fire_7 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l240_1 = ((7'h01 < _zz_when_ArraySlice_l240_1_1) && outputStreamArrayData_1_fire_7);
  assign when_ArraySlice_l241_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l241_1_1);
  assign when_ArraySlice_l244_1 = (_zz_when_ArraySlice_l244_1_1 == 13'h0);
  assign outputStreamArrayData_1_fire_8 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l249_1 = ((_zz_when_ArraySlice_l249_1_1 == 7'h01) && outputStreamArrayData_1_fire_8);
  assign when_ArraySlice_l250_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l250_1_1);
  assign _zz_realValue1_0_27 = (_zz__zz_realValue1_0_27 % _zz__zz_realValue1_0_27_1);
  assign when_ArraySlice_l95_27 = (_zz_realValue1_0_27 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_27) begin
      realValue1_0_27 = (_zz_realValue1_0_27_1 - _zz_realValue1_0_27);
    end else begin
      realValue1_0_27 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_1 = (_zz_when_ArraySlice_l252_1_1 < _zz_when_ArraySlice_l252_1_3);
  always @(*) begin
    debug_0_29 = 1'b0;
    if(when_ArraySlice_l158_232) begin
      if(when_ArraySlice_l159_232) begin
        debug_0_29 = 1'b1;
      end else begin
        debug_0_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_232) begin
        debug_0_29 = 1'b1;
      end else begin
        debug_0_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_29 = 1'b0;
    if(when_ArraySlice_l158_233) begin
      if(when_ArraySlice_l159_233) begin
        debug_1_29 = 1'b1;
      end else begin
        debug_1_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_233) begin
        debug_1_29 = 1'b1;
      end else begin
        debug_1_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_29 = 1'b0;
    if(when_ArraySlice_l158_234) begin
      if(when_ArraySlice_l159_234) begin
        debug_2_29 = 1'b1;
      end else begin
        debug_2_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_234) begin
        debug_2_29 = 1'b1;
      end else begin
        debug_2_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_29 = 1'b0;
    if(when_ArraySlice_l158_235) begin
      if(when_ArraySlice_l159_235) begin
        debug_3_29 = 1'b1;
      end else begin
        debug_3_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_235) begin
        debug_3_29 = 1'b1;
      end else begin
        debug_3_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_29 = 1'b0;
    if(when_ArraySlice_l158_236) begin
      if(when_ArraySlice_l159_236) begin
        debug_4_29 = 1'b1;
      end else begin
        debug_4_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_236) begin
        debug_4_29 = 1'b1;
      end else begin
        debug_4_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_29 = 1'b0;
    if(when_ArraySlice_l158_237) begin
      if(when_ArraySlice_l159_237) begin
        debug_5_29 = 1'b1;
      end else begin
        debug_5_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_237) begin
        debug_5_29 = 1'b1;
      end else begin
        debug_5_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_29 = 1'b0;
    if(when_ArraySlice_l158_238) begin
      if(when_ArraySlice_l159_238) begin
        debug_6_29 = 1'b1;
      end else begin
        debug_6_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_238) begin
        debug_6_29 = 1'b1;
      end else begin
        debug_6_29 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_29 = 1'b0;
    if(when_ArraySlice_l158_239) begin
      if(when_ArraySlice_l159_239) begin
        debug_7_29 = 1'b1;
      end else begin
        debug_7_29 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_239) begin
        debug_7_29 = 1'b1;
      end else begin
        debug_7_29 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_232 = (_zz_when_ArraySlice_l158_232 <= _zz_when_ArraySlice_l158_232_3);
  assign when_ArraySlice_l159_232 = (_zz_when_ArraySlice_l159_232 <= _zz_when_ArraySlice_l159_232_1);
  assign _zz_realValue_0_232 = (_zz__zz_realValue_0_232 % _zz__zz_realValue_0_232_1);
  assign when_ArraySlice_l110_232 = (_zz_realValue_0_232 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_232) begin
      realValue_0_232 = (_zz_realValue_0_232_1 - _zz_realValue_0_232);
    end else begin
      realValue_0_232 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_232 = (_zz_when_ArraySlice_l166_232 <= _zz_when_ArraySlice_l166_232_1);
  assign when_ArraySlice_l158_233 = (_zz_when_ArraySlice_l158_233 <= _zz_when_ArraySlice_l158_233_3);
  assign when_ArraySlice_l159_233 = (_zz_when_ArraySlice_l159_233 <= _zz_when_ArraySlice_l159_233_2);
  assign _zz_realValue_0_233 = (_zz__zz_realValue_0_233 % _zz__zz_realValue_0_233_1);
  assign when_ArraySlice_l110_233 = (_zz_realValue_0_233 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_233) begin
      realValue_0_233 = (_zz_realValue_0_233_1 - _zz_realValue_0_233);
    end else begin
      realValue_0_233 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_233 = (_zz_when_ArraySlice_l166_233 <= _zz_when_ArraySlice_l166_233_2);
  assign when_ArraySlice_l158_234 = (_zz_when_ArraySlice_l158_234 <= _zz_when_ArraySlice_l158_234_3);
  assign when_ArraySlice_l159_234 = (_zz_when_ArraySlice_l159_234 <= _zz_when_ArraySlice_l159_234_2);
  assign _zz_realValue_0_234 = (_zz__zz_realValue_0_234 % _zz__zz_realValue_0_234_1);
  assign when_ArraySlice_l110_234 = (_zz_realValue_0_234 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_234) begin
      realValue_0_234 = (_zz_realValue_0_234_1 - _zz_realValue_0_234);
    end else begin
      realValue_0_234 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_234 = (_zz_when_ArraySlice_l166_234 <= _zz_when_ArraySlice_l166_234_2);
  assign when_ArraySlice_l158_235 = (_zz_when_ArraySlice_l158_235 <= _zz_when_ArraySlice_l158_235_3);
  assign when_ArraySlice_l159_235 = (_zz_when_ArraySlice_l159_235 <= _zz_when_ArraySlice_l159_235_2);
  assign _zz_realValue_0_235 = (_zz__zz_realValue_0_235 % _zz__zz_realValue_0_235_1);
  assign when_ArraySlice_l110_235 = (_zz_realValue_0_235 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_235) begin
      realValue_0_235 = (_zz_realValue_0_235_1 - _zz_realValue_0_235);
    end else begin
      realValue_0_235 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_235 = (_zz_when_ArraySlice_l166_235 <= _zz_when_ArraySlice_l166_235_2);
  assign when_ArraySlice_l158_236 = (_zz_when_ArraySlice_l158_236 <= _zz_when_ArraySlice_l158_236_3);
  assign when_ArraySlice_l159_236 = (_zz_when_ArraySlice_l159_236 <= _zz_when_ArraySlice_l159_236_2);
  assign _zz_realValue_0_236 = (_zz__zz_realValue_0_236 % _zz__zz_realValue_0_236_1);
  assign when_ArraySlice_l110_236 = (_zz_realValue_0_236 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_236) begin
      realValue_0_236 = (_zz_realValue_0_236_1 - _zz_realValue_0_236);
    end else begin
      realValue_0_236 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_236 = (_zz_when_ArraySlice_l166_236 <= _zz_when_ArraySlice_l166_236_2);
  assign when_ArraySlice_l158_237 = (_zz_when_ArraySlice_l158_237 <= _zz_when_ArraySlice_l158_237_3);
  assign when_ArraySlice_l159_237 = (_zz_when_ArraySlice_l159_237 <= _zz_when_ArraySlice_l159_237_2);
  assign _zz_realValue_0_237 = (_zz__zz_realValue_0_237 % _zz__zz_realValue_0_237_1);
  assign when_ArraySlice_l110_237 = (_zz_realValue_0_237 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_237) begin
      realValue_0_237 = (_zz_realValue_0_237_1 - _zz_realValue_0_237);
    end else begin
      realValue_0_237 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_237 = (_zz_when_ArraySlice_l166_237 <= _zz_when_ArraySlice_l166_237_2);
  assign when_ArraySlice_l158_238 = (_zz_when_ArraySlice_l158_238 <= _zz_when_ArraySlice_l158_238_3);
  assign when_ArraySlice_l159_238 = (_zz_when_ArraySlice_l159_238 <= _zz_when_ArraySlice_l159_238_2);
  assign _zz_realValue_0_238 = (_zz__zz_realValue_0_238 % _zz__zz_realValue_0_238_1);
  assign when_ArraySlice_l110_238 = (_zz_realValue_0_238 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_238) begin
      realValue_0_238 = (_zz_realValue_0_238_1 - _zz_realValue_0_238);
    end else begin
      realValue_0_238 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_238 = (_zz_when_ArraySlice_l166_238 <= _zz_when_ArraySlice_l166_238_2);
  assign when_ArraySlice_l158_239 = (_zz_when_ArraySlice_l158_239 <= _zz_when_ArraySlice_l158_239_3);
  assign when_ArraySlice_l159_239 = (_zz_when_ArraySlice_l159_239 <= _zz_when_ArraySlice_l159_239_2);
  assign _zz_realValue_0_239 = (_zz__zz_realValue_0_239 % _zz__zz_realValue_0_239_1);
  assign when_ArraySlice_l110_239 = (_zz_realValue_0_239 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_239) begin
      realValue_0_239 = (_zz_realValue_0_239_1 - _zz_realValue_0_239);
    end else begin
      realValue_0_239 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_239 = (_zz_when_ArraySlice_l166_239 <= _zz_when_ArraySlice_l166_239_2);
  assign when_ArraySlice_l257_1 = (! ((((((_zz_when_ArraySlice_l257_1_1 && _zz_when_ArraySlice_l257_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l257_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_1_4 && _zz_when_ArraySlice_l257_1_5) && (debug_4_29 == _zz_when_ArraySlice_l257_1_6)) && (debug_5_29 == 1'b1)) && (debug_6_29 == 1'b1)) && (debug_7_29 == 1'b1))));
  assign when_ArraySlice_l260_1 = (_zz_when_ArraySlice_l260_1_1 <= _zz_when_ArraySlice_l260_1_2);
  assign when_ArraySlice_l263_1 = (_zz_when_ArraySlice_l263_1_1 <= _zz_when_ArraySlice_l263_1_2);
  assign when_ArraySlice_l270_1 = (_zz_when_ArraySlice_l270_1_1 == 13'h0);
  assign when_ArraySlice_l274_1 = (_zz_when_ArraySlice_l274_1_1 == 7'h0);
  assign outputStreamArrayData_1_fire_9 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l275_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l275_1_1) && outputStreamArrayData_1_fire_9);
  assign _zz_realValue1_0_28 = (_zz__zz_realValue1_0_28 % _zz__zz_realValue1_0_28_1);
  assign when_ArraySlice_l95_28 = (_zz_realValue1_0_28 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_28) begin
      realValue1_0_28 = (_zz_realValue1_0_28_1 - _zz_realValue1_0_28);
    end else begin
      realValue1_0_28 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_1 = (_zz_when_ArraySlice_l277_1_1 < _zz_when_ArraySlice_l277_1_3);
  always @(*) begin
    debug_0_30 = 1'b0;
    if(when_ArraySlice_l158_240) begin
      if(when_ArraySlice_l159_240) begin
        debug_0_30 = 1'b1;
      end else begin
        debug_0_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_240) begin
        debug_0_30 = 1'b1;
      end else begin
        debug_0_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_30 = 1'b0;
    if(when_ArraySlice_l158_241) begin
      if(when_ArraySlice_l159_241) begin
        debug_1_30 = 1'b1;
      end else begin
        debug_1_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_241) begin
        debug_1_30 = 1'b1;
      end else begin
        debug_1_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_30 = 1'b0;
    if(when_ArraySlice_l158_242) begin
      if(when_ArraySlice_l159_242) begin
        debug_2_30 = 1'b1;
      end else begin
        debug_2_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_242) begin
        debug_2_30 = 1'b1;
      end else begin
        debug_2_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_30 = 1'b0;
    if(when_ArraySlice_l158_243) begin
      if(when_ArraySlice_l159_243) begin
        debug_3_30 = 1'b1;
      end else begin
        debug_3_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_243) begin
        debug_3_30 = 1'b1;
      end else begin
        debug_3_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_30 = 1'b0;
    if(when_ArraySlice_l158_244) begin
      if(when_ArraySlice_l159_244) begin
        debug_4_30 = 1'b1;
      end else begin
        debug_4_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_244) begin
        debug_4_30 = 1'b1;
      end else begin
        debug_4_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_30 = 1'b0;
    if(when_ArraySlice_l158_245) begin
      if(when_ArraySlice_l159_245) begin
        debug_5_30 = 1'b1;
      end else begin
        debug_5_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_245) begin
        debug_5_30 = 1'b1;
      end else begin
        debug_5_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_30 = 1'b0;
    if(when_ArraySlice_l158_246) begin
      if(when_ArraySlice_l159_246) begin
        debug_6_30 = 1'b1;
      end else begin
        debug_6_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_246) begin
        debug_6_30 = 1'b1;
      end else begin
        debug_6_30 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_30 = 1'b0;
    if(when_ArraySlice_l158_247) begin
      if(when_ArraySlice_l159_247) begin
        debug_7_30 = 1'b1;
      end else begin
        debug_7_30 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_247) begin
        debug_7_30 = 1'b1;
      end else begin
        debug_7_30 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_240 = (_zz_when_ArraySlice_l158_240 <= _zz_when_ArraySlice_l158_240_3);
  assign when_ArraySlice_l159_240 = (_zz_when_ArraySlice_l159_240 <= _zz_when_ArraySlice_l159_240_1);
  assign _zz_realValue_0_240 = (_zz__zz_realValue_0_240 % _zz__zz_realValue_0_240_1);
  assign when_ArraySlice_l110_240 = (_zz_realValue_0_240 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_240) begin
      realValue_0_240 = (_zz_realValue_0_240_1 - _zz_realValue_0_240);
    end else begin
      realValue_0_240 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_240 = (_zz_when_ArraySlice_l166_240 <= _zz_when_ArraySlice_l166_240_1);
  assign when_ArraySlice_l158_241 = (_zz_when_ArraySlice_l158_241 <= _zz_when_ArraySlice_l158_241_3);
  assign when_ArraySlice_l159_241 = (_zz_when_ArraySlice_l159_241 <= _zz_when_ArraySlice_l159_241_2);
  assign _zz_realValue_0_241 = (_zz__zz_realValue_0_241 % _zz__zz_realValue_0_241_1);
  assign when_ArraySlice_l110_241 = (_zz_realValue_0_241 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_241) begin
      realValue_0_241 = (_zz_realValue_0_241_1 - _zz_realValue_0_241);
    end else begin
      realValue_0_241 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_241 = (_zz_when_ArraySlice_l166_241 <= _zz_when_ArraySlice_l166_241_2);
  assign when_ArraySlice_l158_242 = (_zz_when_ArraySlice_l158_242 <= _zz_when_ArraySlice_l158_242_3);
  assign when_ArraySlice_l159_242 = (_zz_when_ArraySlice_l159_242 <= _zz_when_ArraySlice_l159_242_2);
  assign _zz_realValue_0_242 = (_zz__zz_realValue_0_242 % _zz__zz_realValue_0_242_1);
  assign when_ArraySlice_l110_242 = (_zz_realValue_0_242 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_242) begin
      realValue_0_242 = (_zz_realValue_0_242_1 - _zz_realValue_0_242);
    end else begin
      realValue_0_242 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_242 = (_zz_when_ArraySlice_l166_242 <= _zz_when_ArraySlice_l166_242_2);
  assign when_ArraySlice_l158_243 = (_zz_when_ArraySlice_l158_243 <= _zz_when_ArraySlice_l158_243_3);
  assign when_ArraySlice_l159_243 = (_zz_when_ArraySlice_l159_243 <= _zz_when_ArraySlice_l159_243_2);
  assign _zz_realValue_0_243 = (_zz__zz_realValue_0_243 % _zz__zz_realValue_0_243_1);
  assign when_ArraySlice_l110_243 = (_zz_realValue_0_243 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_243) begin
      realValue_0_243 = (_zz_realValue_0_243_1 - _zz_realValue_0_243);
    end else begin
      realValue_0_243 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_243 = (_zz_when_ArraySlice_l166_243 <= _zz_when_ArraySlice_l166_243_2);
  assign when_ArraySlice_l158_244 = (_zz_when_ArraySlice_l158_244 <= _zz_when_ArraySlice_l158_244_3);
  assign when_ArraySlice_l159_244 = (_zz_when_ArraySlice_l159_244 <= _zz_when_ArraySlice_l159_244_2);
  assign _zz_realValue_0_244 = (_zz__zz_realValue_0_244 % _zz__zz_realValue_0_244_1);
  assign when_ArraySlice_l110_244 = (_zz_realValue_0_244 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_244) begin
      realValue_0_244 = (_zz_realValue_0_244_1 - _zz_realValue_0_244);
    end else begin
      realValue_0_244 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_244 = (_zz_when_ArraySlice_l166_244 <= _zz_when_ArraySlice_l166_244_2);
  assign when_ArraySlice_l158_245 = (_zz_when_ArraySlice_l158_245 <= _zz_when_ArraySlice_l158_245_3);
  assign when_ArraySlice_l159_245 = (_zz_when_ArraySlice_l159_245 <= _zz_when_ArraySlice_l159_245_2);
  assign _zz_realValue_0_245 = (_zz__zz_realValue_0_245 % _zz__zz_realValue_0_245_1);
  assign when_ArraySlice_l110_245 = (_zz_realValue_0_245 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_245) begin
      realValue_0_245 = (_zz_realValue_0_245_1 - _zz_realValue_0_245);
    end else begin
      realValue_0_245 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_245 = (_zz_when_ArraySlice_l166_245 <= _zz_when_ArraySlice_l166_245_2);
  assign when_ArraySlice_l158_246 = (_zz_when_ArraySlice_l158_246 <= _zz_when_ArraySlice_l158_246_3);
  assign when_ArraySlice_l159_246 = (_zz_when_ArraySlice_l159_246 <= _zz_when_ArraySlice_l159_246_2);
  assign _zz_realValue_0_246 = (_zz__zz_realValue_0_246 % _zz__zz_realValue_0_246_1);
  assign when_ArraySlice_l110_246 = (_zz_realValue_0_246 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_246) begin
      realValue_0_246 = (_zz_realValue_0_246_1 - _zz_realValue_0_246);
    end else begin
      realValue_0_246 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_246 = (_zz_when_ArraySlice_l166_246 <= _zz_when_ArraySlice_l166_246_2);
  assign when_ArraySlice_l158_247 = (_zz_when_ArraySlice_l158_247 <= _zz_when_ArraySlice_l158_247_3);
  assign when_ArraySlice_l159_247 = (_zz_when_ArraySlice_l159_247 <= _zz_when_ArraySlice_l159_247_2);
  assign _zz_realValue_0_247 = (_zz__zz_realValue_0_247 % _zz__zz_realValue_0_247_1);
  assign when_ArraySlice_l110_247 = (_zz_realValue_0_247 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_247) begin
      realValue_0_247 = (_zz_realValue_0_247_1 - _zz_realValue_0_247);
    end else begin
      realValue_0_247 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_247 = (_zz_when_ArraySlice_l166_247 <= _zz_when_ArraySlice_l166_247_2);
  assign when_ArraySlice_l282_1 = (! ((((((_zz_when_ArraySlice_l282_1_1 && _zz_when_ArraySlice_l282_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l282_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_1_4 && _zz_when_ArraySlice_l282_1_5) && (debug_4_30 == _zz_when_ArraySlice_l282_1_6)) && (debug_5_30 == 1'b1)) && (debug_6_30 == 1'b1)) && (debug_7_30 == 1'b1))));
  assign when_ArraySlice_l285_1 = (_zz_when_ArraySlice_l285_1_1 <= _zz_when_ArraySlice_l285_1_2);
  assign when_ArraySlice_l288_1 = (_zz_when_ArraySlice_l288_1_1 <= _zz_when_ArraySlice_l288_1_2);
  assign outputStreamArrayData_1_fire_10 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l295_1 = ((_zz_when_ArraySlice_l295_1_1 == 13'h0) && outputStreamArrayData_1_fire_10);
  assign outputStreamArrayData_1_fire_11 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l306_1 = ((handshakeTimes_1_value == _zz_when_ArraySlice_l306_1_1) && outputStreamArrayData_1_fire_11);
  assign _zz_realValue1_0_29 = (_zz__zz_realValue1_0_29 % _zz__zz_realValue1_0_29_1);
  assign when_ArraySlice_l95_29 = (_zz_realValue1_0_29 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_29) begin
      realValue1_0_29 = (_zz_realValue1_0_29_1 - _zz_realValue1_0_29);
    end else begin
      realValue1_0_29 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_1 = (_zz_when_ArraySlice_l307_1_1 < _zz_when_ArraySlice_l307_1_3);
  always @(*) begin
    debug_0_31 = 1'b0;
    if(when_ArraySlice_l158_248) begin
      if(when_ArraySlice_l159_248) begin
        debug_0_31 = 1'b1;
      end else begin
        debug_0_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_248) begin
        debug_0_31 = 1'b1;
      end else begin
        debug_0_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_31 = 1'b0;
    if(when_ArraySlice_l158_249) begin
      if(when_ArraySlice_l159_249) begin
        debug_1_31 = 1'b1;
      end else begin
        debug_1_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_249) begin
        debug_1_31 = 1'b1;
      end else begin
        debug_1_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_31 = 1'b0;
    if(when_ArraySlice_l158_250) begin
      if(when_ArraySlice_l159_250) begin
        debug_2_31 = 1'b1;
      end else begin
        debug_2_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_250) begin
        debug_2_31 = 1'b1;
      end else begin
        debug_2_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_31 = 1'b0;
    if(when_ArraySlice_l158_251) begin
      if(when_ArraySlice_l159_251) begin
        debug_3_31 = 1'b1;
      end else begin
        debug_3_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_251) begin
        debug_3_31 = 1'b1;
      end else begin
        debug_3_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_31 = 1'b0;
    if(when_ArraySlice_l158_252) begin
      if(when_ArraySlice_l159_252) begin
        debug_4_31 = 1'b1;
      end else begin
        debug_4_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_252) begin
        debug_4_31 = 1'b1;
      end else begin
        debug_4_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_31 = 1'b0;
    if(when_ArraySlice_l158_253) begin
      if(when_ArraySlice_l159_253) begin
        debug_5_31 = 1'b1;
      end else begin
        debug_5_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_253) begin
        debug_5_31 = 1'b1;
      end else begin
        debug_5_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_31 = 1'b0;
    if(when_ArraySlice_l158_254) begin
      if(when_ArraySlice_l159_254) begin
        debug_6_31 = 1'b1;
      end else begin
        debug_6_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_254) begin
        debug_6_31 = 1'b1;
      end else begin
        debug_6_31 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_31 = 1'b0;
    if(when_ArraySlice_l158_255) begin
      if(when_ArraySlice_l159_255) begin
        debug_7_31 = 1'b1;
      end else begin
        debug_7_31 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_255) begin
        debug_7_31 = 1'b1;
      end else begin
        debug_7_31 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_248 = (_zz_when_ArraySlice_l158_248 <= _zz_when_ArraySlice_l158_248_3);
  assign when_ArraySlice_l159_248 = (_zz_when_ArraySlice_l159_248 <= _zz_when_ArraySlice_l159_248_1);
  assign _zz_realValue_0_248 = (_zz__zz_realValue_0_248 % _zz__zz_realValue_0_248_1);
  assign when_ArraySlice_l110_248 = (_zz_realValue_0_248 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_248) begin
      realValue_0_248 = (_zz_realValue_0_248_1 - _zz_realValue_0_248);
    end else begin
      realValue_0_248 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_248 = (_zz_when_ArraySlice_l166_248 <= _zz_when_ArraySlice_l166_248_1);
  assign when_ArraySlice_l158_249 = (_zz_when_ArraySlice_l158_249 <= _zz_when_ArraySlice_l158_249_3);
  assign when_ArraySlice_l159_249 = (_zz_when_ArraySlice_l159_249 <= _zz_when_ArraySlice_l159_249_2);
  assign _zz_realValue_0_249 = (_zz__zz_realValue_0_249 % _zz__zz_realValue_0_249_1);
  assign when_ArraySlice_l110_249 = (_zz_realValue_0_249 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_249) begin
      realValue_0_249 = (_zz_realValue_0_249_1 - _zz_realValue_0_249);
    end else begin
      realValue_0_249 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_249 = (_zz_when_ArraySlice_l166_249 <= _zz_when_ArraySlice_l166_249_2);
  assign when_ArraySlice_l158_250 = (_zz_when_ArraySlice_l158_250 <= _zz_when_ArraySlice_l158_250_3);
  assign when_ArraySlice_l159_250 = (_zz_when_ArraySlice_l159_250 <= _zz_when_ArraySlice_l159_250_2);
  assign _zz_realValue_0_250 = (_zz__zz_realValue_0_250 % _zz__zz_realValue_0_250_1);
  assign when_ArraySlice_l110_250 = (_zz_realValue_0_250 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_250) begin
      realValue_0_250 = (_zz_realValue_0_250_1 - _zz_realValue_0_250);
    end else begin
      realValue_0_250 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_250 = (_zz_when_ArraySlice_l166_250 <= _zz_when_ArraySlice_l166_250_2);
  assign when_ArraySlice_l158_251 = (_zz_when_ArraySlice_l158_251 <= _zz_when_ArraySlice_l158_251_3);
  assign when_ArraySlice_l159_251 = (_zz_when_ArraySlice_l159_251 <= _zz_when_ArraySlice_l159_251_2);
  assign _zz_realValue_0_251 = (_zz__zz_realValue_0_251 % _zz__zz_realValue_0_251_1);
  assign when_ArraySlice_l110_251 = (_zz_realValue_0_251 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_251) begin
      realValue_0_251 = (_zz_realValue_0_251_1 - _zz_realValue_0_251);
    end else begin
      realValue_0_251 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_251 = (_zz_when_ArraySlice_l166_251 <= _zz_when_ArraySlice_l166_251_2);
  assign when_ArraySlice_l158_252 = (_zz_when_ArraySlice_l158_252 <= _zz_when_ArraySlice_l158_252_3);
  assign when_ArraySlice_l159_252 = (_zz_when_ArraySlice_l159_252 <= _zz_when_ArraySlice_l159_252_2);
  assign _zz_realValue_0_252 = (_zz__zz_realValue_0_252 % _zz__zz_realValue_0_252_1);
  assign when_ArraySlice_l110_252 = (_zz_realValue_0_252 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_252) begin
      realValue_0_252 = (_zz_realValue_0_252_1 - _zz_realValue_0_252);
    end else begin
      realValue_0_252 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_252 = (_zz_when_ArraySlice_l166_252 <= _zz_when_ArraySlice_l166_252_2);
  assign when_ArraySlice_l158_253 = (_zz_when_ArraySlice_l158_253 <= _zz_when_ArraySlice_l158_253_3);
  assign when_ArraySlice_l159_253 = (_zz_when_ArraySlice_l159_253 <= _zz_when_ArraySlice_l159_253_2);
  assign _zz_realValue_0_253 = (_zz__zz_realValue_0_253 % _zz__zz_realValue_0_253_1);
  assign when_ArraySlice_l110_253 = (_zz_realValue_0_253 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_253) begin
      realValue_0_253 = (_zz_realValue_0_253_1 - _zz_realValue_0_253);
    end else begin
      realValue_0_253 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_253 = (_zz_when_ArraySlice_l166_253 <= _zz_when_ArraySlice_l166_253_2);
  assign when_ArraySlice_l158_254 = (_zz_when_ArraySlice_l158_254 <= _zz_when_ArraySlice_l158_254_3);
  assign when_ArraySlice_l159_254 = (_zz_when_ArraySlice_l159_254 <= _zz_when_ArraySlice_l159_254_2);
  assign _zz_realValue_0_254 = (_zz__zz_realValue_0_254 % _zz__zz_realValue_0_254_1);
  assign when_ArraySlice_l110_254 = (_zz_realValue_0_254 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_254) begin
      realValue_0_254 = (_zz_realValue_0_254_1 - _zz_realValue_0_254);
    end else begin
      realValue_0_254 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_254 = (_zz_when_ArraySlice_l166_254 <= _zz_when_ArraySlice_l166_254_2);
  assign when_ArraySlice_l158_255 = (_zz_when_ArraySlice_l158_255 <= _zz_when_ArraySlice_l158_255_3);
  assign when_ArraySlice_l159_255 = (_zz_when_ArraySlice_l159_255 <= _zz_when_ArraySlice_l159_255_2);
  assign _zz_realValue_0_255 = (_zz__zz_realValue_0_255 % _zz__zz_realValue_0_255_1);
  assign when_ArraySlice_l110_255 = (_zz_realValue_0_255 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_255) begin
      realValue_0_255 = (_zz_realValue_0_255_1 - _zz_realValue_0_255);
    end else begin
      realValue_0_255 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_255 = (_zz_when_ArraySlice_l166_255 <= _zz_when_ArraySlice_l166_255_2);
  assign when_ArraySlice_l314_1 = (! ((((((_zz_when_ArraySlice_l314_1_1 && _zz_when_ArraySlice_l314_1_2) && (holdReadOp_4 == _zz_when_ArraySlice_l314_1_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_1_4 && _zz_when_ArraySlice_l314_1_5) && (debug_4_31 == _zz_when_ArraySlice_l314_1_6)) && (debug_5_31 == 1'b1)) && (debug_6_31 == 1'b1)) && (debug_7_31 == 1'b1))));
  assign outputStreamArrayData_1_fire_12 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l318_1 = ((_zz_when_ArraySlice_l318_1_1 == 13'h0) && outputStreamArrayData_1_fire_12);
  assign when_ArraySlice_l304_1 = (allowPadding_1 && (_zz_when_ArraySlice_l304_1_1 <= _zz_when_ArraySlice_l304_1_2));
  assign outputStreamArrayData_1_fire_13 = (outputStreamArrayData_1_valid && outputStreamArrayData_1_ready);
  assign when_ArraySlice_l325_1 = (handshakeTimes_1_value == _zz_when_ArraySlice_l325_1_1);
  assign when_ArraySlice_l233_2 = (_zz_when_ArraySlice_l233_2_1 < _zz_when_ArraySlice_l233_2_4);
  assign when_ArraySlice_l234_2 = ((! holdReadOp_2) && (_zz_when_ArraySlice_l234_2_1 != 7'h0));
  assign _zz_outputStreamArrayData_2_valid_1 = (selectReadFifo_2 + _zz__zz_outputStreamArrayData_2_valid_1_1);
  assign _zz_13 = ({127'd0,1'b1} <<< _zz__zz_13);
  assign _zz_io_pop_ready_10 = outputStreamArrayData_2_ready;
  assign when_ArraySlice_l239_2 = (! holdReadOp_2);
  assign outputStreamArrayData_2_fire_7 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l240_2 = ((7'h01 < _zz_when_ArraySlice_l240_2_1) && outputStreamArrayData_2_fire_7);
  assign when_ArraySlice_l241_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l241_2_1);
  assign when_ArraySlice_l244_2 = (_zz_when_ArraySlice_l244_2 == 13'h0);
  assign outputStreamArrayData_2_fire_8 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l249_2 = ((_zz_when_ArraySlice_l249_2_1 == 7'h01) && outputStreamArrayData_2_fire_8);
  assign when_ArraySlice_l250_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l250_2_1);
  assign _zz_realValue1_0_30 = (_zz__zz_realValue1_0_30 % _zz__zz_realValue1_0_30_1);
  assign when_ArraySlice_l95_30 = (_zz_realValue1_0_30 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_30) begin
      realValue1_0_30 = (_zz_realValue1_0_30_1 - _zz_realValue1_0_30);
    end else begin
      realValue1_0_30 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_2 = (_zz_when_ArraySlice_l252_2_1 < _zz_when_ArraySlice_l252_2_3);
  always @(*) begin
    debug_0_32 = 1'b0;
    if(when_ArraySlice_l158_256) begin
      if(when_ArraySlice_l159_256) begin
        debug_0_32 = 1'b1;
      end else begin
        debug_0_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_256) begin
        debug_0_32 = 1'b1;
      end else begin
        debug_0_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_32 = 1'b0;
    if(when_ArraySlice_l158_257) begin
      if(when_ArraySlice_l159_257) begin
        debug_1_32 = 1'b1;
      end else begin
        debug_1_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_257) begin
        debug_1_32 = 1'b1;
      end else begin
        debug_1_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_32 = 1'b0;
    if(when_ArraySlice_l158_258) begin
      if(when_ArraySlice_l159_258) begin
        debug_2_32 = 1'b1;
      end else begin
        debug_2_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_258) begin
        debug_2_32 = 1'b1;
      end else begin
        debug_2_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_32 = 1'b0;
    if(when_ArraySlice_l158_259) begin
      if(when_ArraySlice_l159_259) begin
        debug_3_32 = 1'b1;
      end else begin
        debug_3_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_259) begin
        debug_3_32 = 1'b1;
      end else begin
        debug_3_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_32 = 1'b0;
    if(when_ArraySlice_l158_260) begin
      if(when_ArraySlice_l159_260) begin
        debug_4_32 = 1'b1;
      end else begin
        debug_4_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_260) begin
        debug_4_32 = 1'b1;
      end else begin
        debug_4_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_32 = 1'b0;
    if(when_ArraySlice_l158_261) begin
      if(when_ArraySlice_l159_261) begin
        debug_5_32 = 1'b1;
      end else begin
        debug_5_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_261) begin
        debug_5_32 = 1'b1;
      end else begin
        debug_5_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_32 = 1'b0;
    if(when_ArraySlice_l158_262) begin
      if(when_ArraySlice_l159_262) begin
        debug_6_32 = 1'b1;
      end else begin
        debug_6_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_262) begin
        debug_6_32 = 1'b1;
      end else begin
        debug_6_32 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_32 = 1'b0;
    if(when_ArraySlice_l158_263) begin
      if(when_ArraySlice_l159_263) begin
        debug_7_32 = 1'b1;
      end else begin
        debug_7_32 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_263) begin
        debug_7_32 = 1'b1;
      end else begin
        debug_7_32 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_256 = (_zz_when_ArraySlice_l158_256 <= _zz_when_ArraySlice_l158_256_3);
  assign when_ArraySlice_l159_256 = (_zz_when_ArraySlice_l159_256 <= _zz_when_ArraySlice_l159_256_1);
  assign _zz_realValue_0_256 = (_zz__zz_realValue_0_256 % _zz__zz_realValue_0_256_1);
  assign when_ArraySlice_l110_256 = (_zz_realValue_0_256 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_256) begin
      realValue_0_256 = (_zz_realValue_0_256_1 - _zz_realValue_0_256);
    end else begin
      realValue_0_256 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_256 = (_zz_when_ArraySlice_l166_256 <= _zz_when_ArraySlice_l166_256_1);
  assign when_ArraySlice_l158_257 = (_zz_when_ArraySlice_l158_257 <= _zz_when_ArraySlice_l158_257_3);
  assign when_ArraySlice_l159_257 = (_zz_when_ArraySlice_l159_257 <= _zz_when_ArraySlice_l159_257_2);
  assign _zz_realValue_0_257 = (_zz__zz_realValue_0_257 % _zz__zz_realValue_0_257_1);
  assign when_ArraySlice_l110_257 = (_zz_realValue_0_257 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_257) begin
      realValue_0_257 = (_zz_realValue_0_257_1 - _zz_realValue_0_257);
    end else begin
      realValue_0_257 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_257 = (_zz_when_ArraySlice_l166_257 <= _zz_when_ArraySlice_l166_257_2);
  assign when_ArraySlice_l158_258 = (_zz_when_ArraySlice_l158_258 <= _zz_when_ArraySlice_l158_258_3);
  assign when_ArraySlice_l159_258 = (_zz_when_ArraySlice_l159_258 <= _zz_when_ArraySlice_l159_258_2);
  assign _zz_realValue_0_258 = (_zz__zz_realValue_0_258 % _zz__zz_realValue_0_258_1);
  assign when_ArraySlice_l110_258 = (_zz_realValue_0_258 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_258) begin
      realValue_0_258 = (_zz_realValue_0_258_1 - _zz_realValue_0_258);
    end else begin
      realValue_0_258 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_258 = (_zz_when_ArraySlice_l166_258 <= _zz_when_ArraySlice_l166_258_2);
  assign when_ArraySlice_l158_259 = (_zz_when_ArraySlice_l158_259 <= _zz_when_ArraySlice_l158_259_3);
  assign when_ArraySlice_l159_259 = (_zz_when_ArraySlice_l159_259 <= _zz_when_ArraySlice_l159_259_2);
  assign _zz_realValue_0_259 = (_zz__zz_realValue_0_259 % _zz__zz_realValue_0_259_1);
  assign when_ArraySlice_l110_259 = (_zz_realValue_0_259 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_259) begin
      realValue_0_259 = (_zz_realValue_0_259_1 - _zz_realValue_0_259);
    end else begin
      realValue_0_259 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_259 = (_zz_when_ArraySlice_l166_259 <= _zz_when_ArraySlice_l166_259_2);
  assign when_ArraySlice_l158_260 = (_zz_when_ArraySlice_l158_260 <= _zz_when_ArraySlice_l158_260_3);
  assign when_ArraySlice_l159_260 = (_zz_when_ArraySlice_l159_260 <= _zz_when_ArraySlice_l159_260_2);
  assign _zz_realValue_0_260 = (_zz__zz_realValue_0_260 % _zz__zz_realValue_0_260_1);
  assign when_ArraySlice_l110_260 = (_zz_realValue_0_260 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_260) begin
      realValue_0_260 = (_zz_realValue_0_260_1 - _zz_realValue_0_260);
    end else begin
      realValue_0_260 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_260 = (_zz_when_ArraySlice_l166_260 <= _zz_when_ArraySlice_l166_260_2);
  assign when_ArraySlice_l158_261 = (_zz_when_ArraySlice_l158_261 <= _zz_when_ArraySlice_l158_261_3);
  assign when_ArraySlice_l159_261 = (_zz_when_ArraySlice_l159_261 <= _zz_when_ArraySlice_l159_261_2);
  assign _zz_realValue_0_261 = (_zz__zz_realValue_0_261 % _zz__zz_realValue_0_261_1);
  assign when_ArraySlice_l110_261 = (_zz_realValue_0_261 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_261) begin
      realValue_0_261 = (_zz_realValue_0_261_1 - _zz_realValue_0_261);
    end else begin
      realValue_0_261 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_261 = (_zz_when_ArraySlice_l166_261 <= _zz_when_ArraySlice_l166_261_2);
  assign when_ArraySlice_l158_262 = (_zz_when_ArraySlice_l158_262 <= _zz_when_ArraySlice_l158_262_3);
  assign when_ArraySlice_l159_262 = (_zz_when_ArraySlice_l159_262 <= _zz_when_ArraySlice_l159_262_2);
  assign _zz_realValue_0_262 = (_zz__zz_realValue_0_262 % _zz__zz_realValue_0_262_1);
  assign when_ArraySlice_l110_262 = (_zz_realValue_0_262 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_262) begin
      realValue_0_262 = (_zz_realValue_0_262_1 - _zz_realValue_0_262);
    end else begin
      realValue_0_262 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_262 = (_zz_when_ArraySlice_l166_262 <= _zz_when_ArraySlice_l166_262_2);
  assign when_ArraySlice_l158_263 = (_zz_when_ArraySlice_l158_263 <= _zz_when_ArraySlice_l158_263_3);
  assign when_ArraySlice_l159_263 = (_zz_when_ArraySlice_l159_263 <= _zz_when_ArraySlice_l159_263_2);
  assign _zz_realValue_0_263 = (_zz__zz_realValue_0_263 % _zz__zz_realValue_0_263_1);
  assign when_ArraySlice_l110_263 = (_zz_realValue_0_263 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_263) begin
      realValue_0_263 = (_zz_realValue_0_263_1 - _zz_realValue_0_263);
    end else begin
      realValue_0_263 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_263 = (_zz_when_ArraySlice_l166_263 <= _zz_when_ArraySlice_l166_263_2);
  assign when_ArraySlice_l257_2 = (! ((((((_zz_when_ArraySlice_l257_2_1 && _zz_when_ArraySlice_l257_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l257_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_2_4 && _zz_when_ArraySlice_l257_2_5) && (debug_4_32 == _zz_when_ArraySlice_l257_2_6)) && (debug_5_32 == 1'b1)) && (debug_6_32 == 1'b1)) && (debug_7_32 == 1'b1))));
  assign when_ArraySlice_l260_2 = (_zz_when_ArraySlice_l260_2_1 <= _zz_when_ArraySlice_l260_2_2);
  assign when_ArraySlice_l263_2 = (_zz_when_ArraySlice_l263_2_1 <= _zz_when_ArraySlice_l263_2_2);
  assign when_ArraySlice_l270_2 = (_zz_when_ArraySlice_l270_2 == 13'h0);
  assign when_ArraySlice_l274_2 = (_zz_when_ArraySlice_l274_2_1 == 7'h0);
  assign outputStreamArrayData_2_fire_9 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l275_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l275_2_1) && outputStreamArrayData_2_fire_9);
  assign _zz_realValue1_0_31 = (_zz__zz_realValue1_0_31 % _zz__zz_realValue1_0_31_1);
  assign when_ArraySlice_l95_31 = (_zz_realValue1_0_31 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_31) begin
      realValue1_0_31 = (_zz_realValue1_0_31_1 - _zz_realValue1_0_31);
    end else begin
      realValue1_0_31 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_2 = (_zz_when_ArraySlice_l277_2_1 < _zz_when_ArraySlice_l277_2_3);
  always @(*) begin
    debug_0_33 = 1'b0;
    if(when_ArraySlice_l158_264) begin
      if(when_ArraySlice_l159_264) begin
        debug_0_33 = 1'b1;
      end else begin
        debug_0_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_264) begin
        debug_0_33 = 1'b1;
      end else begin
        debug_0_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_33 = 1'b0;
    if(when_ArraySlice_l158_265) begin
      if(when_ArraySlice_l159_265) begin
        debug_1_33 = 1'b1;
      end else begin
        debug_1_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_265) begin
        debug_1_33 = 1'b1;
      end else begin
        debug_1_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_33 = 1'b0;
    if(when_ArraySlice_l158_266) begin
      if(when_ArraySlice_l159_266) begin
        debug_2_33 = 1'b1;
      end else begin
        debug_2_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_266) begin
        debug_2_33 = 1'b1;
      end else begin
        debug_2_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_33 = 1'b0;
    if(when_ArraySlice_l158_267) begin
      if(when_ArraySlice_l159_267) begin
        debug_3_33 = 1'b1;
      end else begin
        debug_3_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_267) begin
        debug_3_33 = 1'b1;
      end else begin
        debug_3_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_33 = 1'b0;
    if(when_ArraySlice_l158_268) begin
      if(when_ArraySlice_l159_268) begin
        debug_4_33 = 1'b1;
      end else begin
        debug_4_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_268) begin
        debug_4_33 = 1'b1;
      end else begin
        debug_4_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_33 = 1'b0;
    if(when_ArraySlice_l158_269) begin
      if(when_ArraySlice_l159_269) begin
        debug_5_33 = 1'b1;
      end else begin
        debug_5_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_269) begin
        debug_5_33 = 1'b1;
      end else begin
        debug_5_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_33 = 1'b0;
    if(when_ArraySlice_l158_270) begin
      if(when_ArraySlice_l159_270) begin
        debug_6_33 = 1'b1;
      end else begin
        debug_6_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_270) begin
        debug_6_33 = 1'b1;
      end else begin
        debug_6_33 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_33 = 1'b0;
    if(when_ArraySlice_l158_271) begin
      if(when_ArraySlice_l159_271) begin
        debug_7_33 = 1'b1;
      end else begin
        debug_7_33 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_271) begin
        debug_7_33 = 1'b1;
      end else begin
        debug_7_33 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_264 = (_zz_when_ArraySlice_l158_264 <= _zz_when_ArraySlice_l158_264_3);
  assign when_ArraySlice_l159_264 = (_zz_when_ArraySlice_l159_264 <= _zz_when_ArraySlice_l159_264_1);
  assign _zz_realValue_0_264 = (_zz__zz_realValue_0_264 % _zz__zz_realValue_0_264_1);
  assign when_ArraySlice_l110_264 = (_zz_realValue_0_264 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_264) begin
      realValue_0_264 = (_zz_realValue_0_264_1 - _zz_realValue_0_264);
    end else begin
      realValue_0_264 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_264 = (_zz_when_ArraySlice_l166_264 <= _zz_when_ArraySlice_l166_264_1);
  assign when_ArraySlice_l158_265 = (_zz_when_ArraySlice_l158_265 <= _zz_when_ArraySlice_l158_265_3);
  assign when_ArraySlice_l159_265 = (_zz_when_ArraySlice_l159_265 <= _zz_when_ArraySlice_l159_265_2);
  assign _zz_realValue_0_265 = (_zz__zz_realValue_0_265 % _zz__zz_realValue_0_265_1);
  assign when_ArraySlice_l110_265 = (_zz_realValue_0_265 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_265) begin
      realValue_0_265 = (_zz_realValue_0_265_1 - _zz_realValue_0_265);
    end else begin
      realValue_0_265 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_265 = (_zz_when_ArraySlice_l166_265 <= _zz_when_ArraySlice_l166_265_2);
  assign when_ArraySlice_l158_266 = (_zz_when_ArraySlice_l158_266 <= _zz_when_ArraySlice_l158_266_3);
  assign when_ArraySlice_l159_266 = (_zz_when_ArraySlice_l159_266 <= _zz_when_ArraySlice_l159_266_2);
  assign _zz_realValue_0_266 = (_zz__zz_realValue_0_266 % _zz__zz_realValue_0_266_1);
  assign when_ArraySlice_l110_266 = (_zz_realValue_0_266 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_266) begin
      realValue_0_266 = (_zz_realValue_0_266_1 - _zz_realValue_0_266);
    end else begin
      realValue_0_266 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_266 = (_zz_when_ArraySlice_l166_266 <= _zz_when_ArraySlice_l166_266_2);
  assign when_ArraySlice_l158_267 = (_zz_when_ArraySlice_l158_267 <= _zz_when_ArraySlice_l158_267_3);
  assign when_ArraySlice_l159_267 = (_zz_when_ArraySlice_l159_267 <= _zz_when_ArraySlice_l159_267_2);
  assign _zz_realValue_0_267 = (_zz__zz_realValue_0_267 % _zz__zz_realValue_0_267_1);
  assign when_ArraySlice_l110_267 = (_zz_realValue_0_267 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_267) begin
      realValue_0_267 = (_zz_realValue_0_267_1 - _zz_realValue_0_267);
    end else begin
      realValue_0_267 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_267 = (_zz_when_ArraySlice_l166_267 <= _zz_when_ArraySlice_l166_267_2);
  assign when_ArraySlice_l158_268 = (_zz_when_ArraySlice_l158_268 <= _zz_when_ArraySlice_l158_268_3);
  assign when_ArraySlice_l159_268 = (_zz_when_ArraySlice_l159_268 <= _zz_when_ArraySlice_l159_268_2);
  assign _zz_realValue_0_268 = (_zz__zz_realValue_0_268 % _zz__zz_realValue_0_268_1);
  assign when_ArraySlice_l110_268 = (_zz_realValue_0_268 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_268) begin
      realValue_0_268 = (_zz_realValue_0_268_1 - _zz_realValue_0_268);
    end else begin
      realValue_0_268 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_268 = (_zz_when_ArraySlice_l166_268 <= _zz_when_ArraySlice_l166_268_2);
  assign when_ArraySlice_l158_269 = (_zz_when_ArraySlice_l158_269 <= _zz_when_ArraySlice_l158_269_3);
  assign when_ArraySlice_l159_269 = (_zz_when_ArraySlice_l159_269 <= _zz_when_ArraySlice_l159_269_2);
  assign _zz_realValue_0_269 = (_zz__zz_realValue_0_269 % _zz__zz_realValue_0_269_1);
  assign when_ArraySlice_l110_269 = (_zz_realValue_0_269 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_269) begin
      realValue_0_269 = (_zz_realValue_0_269_1 - _zz_realValue_0_269);
    end else begin
      realValue_0_269 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_269 = (_zz_when_ArraySlice_l166_269 <= _zz_when_ArraySlice_l166_269_2);
  assign when_ArraySlice_l158_270 = (_zz_when_ArraySlice_l158_270 <= _zz_when_ArraySlice_l158_270_3);
  assign when_ArraySlice_l159_270 = (_zz_when_ArraySlice_l159_270 <= _zz_when_ArraySlice_l159_270_2);
  assign _zz_realValue_0_270 = (_zz__zz_realValue_0_270 % _zz__zz_realValue_0_270_1);
  assign when_ArraySlice_l110_270 = (_zz_realValue_0_270 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_270) begin
      realValue_0_270 = (_zz_realValue_0_270_1 - _zz_realValue_0_270);
    end else begin
      realValue_0_270 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_270 = (_zz_when_ArraySlice_l166_270 <= _zz_when_ArraySlice_l166_270_2);
  assign when_ArraySlice_l158_271 = (_zz_when_ArraySlice_l158_271 <= _zz_when_ArraySlice_l158_271_3);
  assign when_ArraySlice_l159_271 = (_zz_when_ArraySlice_l159_271 <= _zz_when_ArraySlice_l159_271_2);
  assign _zz_realValue_0_271 = (_zz__zz_realValue_0_271 % _zz__zz_realValue_0_271_1);
  assign when_ArraySlice_l110_271 = (_zz_realValue_0_271 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_271) begin
      realValue_0_271 = (_zz_realValue_0_271_1 - _zz_realValue_0_271);
    end else begin
      realValue_0_271 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_271 = (_zz_when_ArraySlice_l166_271 <= _zz_when_ArraySlice_l166_271_2);
  assign when_ArraySlice_l282_2 = (! ((((((_zz_when_ArraySlice_l282_2_1 && _zz_when_ArraySlice_l282_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l282_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_2_4 && _zz_when_ArraySlice_l282_2_5) && (debug_4_33 == _zz_when_ArraySlice_l282_2_6)) && (debug_5_33 == 1'b1)) && (debug_6_33 == 1'b1)) && (debug_7_33 == 1'b1))));
  assign when_ArraySlice_l285_2 = (_zz_when_ArraySlice_l285_2_1 <= _zz_when_ArraySlice_l285_2_2);
  assign when_ArraySlice_l288_2 = (_zz_when_ArraySlice_l288_2_1 <= _zz_when_ArraySlice_l288_2_2);
  assign outputStreamArrayData_2_fire_10 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l295_2 = ((_zz_when_ArraySlice_l295_2 == 13'h0) && outputStreamArrayData_2_fire_10);
  assign outputStreamArrayData_2_fire_11 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l306_2 = ((handshakeTimes_2_value == _zz_when_ArraySlice_l306_2_1) && outputStreamArrayData_2_fire_11);
  assign _zz_realValue1_0_32 = (_zz__zz_realValue1_0_32 % _zz__zz_realValue1_0_32_1);
  assign when_ArraySlice_l95_32 = (_zz_realValue1_0_32 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_32) begin
      realValue1_0_32 = (_zz_realValue1_0_32_1 - _zz_realValue1_0_32);
    end else begin
      realValue1_0_32 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_2 = (_zz_when_ArraySlice_l307_2_1 < _zz_when_ArraySlice_l307_2_3);
  always @(*) begin
    debug_0_34 = 1'b0;
    if(when_ArraySlice_l158_272) begin
      if(when_ArraySlice_l159_272) begin
        debug_0_34 = 1'b1;
      end else begin
        debug_0_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_272) begin
        debug_0_34 = 1'b1;
      end else begin
        debug_0_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_34 = 1'b0;
    if(when_ArraySlice_l158_273) begin
      if(when_ArraySlice_l159_273) begin
        debug_1_34 = 1'b1;
      end else begin
        debug_1_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_273) begin
        debug_1_34 = 1'b1;
      end else begin
        debug_1_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_34 = 1'b0;
    if(when_ArraySlice_l158_274) begin
      if(when_ArraySlice_l159_274) begin
        debug_2_34 = 1'b1;
      end else begin
        debug_2_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_274) begin
        debug_2_34 = 1'b1;
      end else begin
        debug_2_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_34 = 1'b0;
    if(when_ArraySlice_l158_275) begin
      if(when_ArraySlice_l159_275) begin
        debug_3_34 = 1'b1;
      end else begin
        debug_3_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_275) begin
        debug_3_34 = 1'b1;
      end else begin
        debug_3_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_34 = 1'b0;
    if(when_ArraySlice_l158_276) begin
      if(when_ArraySlice_l159_276) begin
        debug_4_34 = 1'b1;
      end else begin
        debug_4_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_276) begin
        debug_4_34 = 1'b1;
      end else begin
        debug_4_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_34 = 1'b0;
    if(when_ArraySlice_l158_277) begin
      if(when_ArraySlice_l159_277) begin
        debug_5_34 = 1'b1;
      end else begin
        debug_5_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_277) begin
        debug_5_34 = 1'b1;
      end else begin
        debug_5_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_34 = 1'b0;
    if(when_ArraySlice_l158_278) begin
      if(when_ArraySlice_l159_278) begin
        debug_6_34 = 1'b1;
      end else begin
        debug_6_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_278) begin
        debug_6_34 = 1'b1;
      end else begin
        debug_6_34 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_34 = 1'b0;
    if(when_ArraySlice_l158_279) begin
      if(when_ArraySlice_l159_279) begin
        debug_7_34 = 1'b1;
      end else begin
        debug_7_34 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_279) begin
        debug_7_34 = 1'b1;
      end else begin
        debug_7_34 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_272 = (_zz_when_ArraySlice_l158_272 <= _zz_when_ArraySlice_l158_272_3);
  assign when_ArraySlice_l159_272 = (_zz_when_ArraySlice_l159_272 <= _zz_when_ArraySlice_l159_272_1);
  assign _zz_realValue_0_272 = (_zz__zz_realValue_0_272 % _zz__zz_realValue_0_272_1);
  assign when_ArraySlice_l110_272 = (_zz_realValue_0_272 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_272) begin
      realValue_0_272 = (_zz_realValue_0_272_1 - _zz_realValue_0_272);
    end else begin
      realValue_0_272 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_272 = (_zz_when_ArraySlice_l166_272 <= _zz_when_ArraySlice_l166_272_1);
  assign when_ArraySlice_l158_273 = (_zz_when_ArraySlice_l158_273 <= _zz_when_ArraySlice_l158_273_3);
  assign when_ArraySlice_l159_273 = (_zz_when_ArraySlice_l159_273 <= _zz_when_ArraySlice_l159_273_2);
  assign _zz_realValue_0_273 = (_zz__zz_realValue_0_273 % _zz__zz_realValue_0_273_1);
  assign when_ArraySlice_l110_273 = (_zz_realValue_0_273 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_273) begin
      realValue_0_273 = (_zz_realValue_0_273_1 - _zz_realValue_0_273);
    end else begin
      realValue_0_273 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_273 = (_zz_when_ArraySlice_l166_273 <= _zz_when_ArraySlice_l166_273_2);
  assign when_ArraySlice_l158_274 = (_zz_when_ArraySlice_l158_274 <= _zz_when_ArraySlice_l158_274_3);
  assign when_ArraySlice_l159_274 = (_zz_when_ArraySlice_l159_274 <= _zz_when_ArraySlice_l159_274_2);
  assign _zz_realValue_0_274 = (_zz__zz_realValue_0_274 % _zz__zz_realValue_0_274_1);
  assign when_ArraySlice_l110_274 = (_zz_realValue_0_274 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_274) begin
      realValue_0_274 = (_zz_realValue_0_274_1 - _zz_realValue_0_274);
    end else begin
      realValue_0_274 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_274 = (_zz_when_ArraySlice_l166_274 <= _zz_when_ArraySlice_l166_274_2);
  assign when_ArraySlice_l158_275 = (_zz_when_ArraySlice_l158_275 <= _zz_when_ArraySlice_l158_275_3);
  assign when_ArraySlice_l159_275 = (_zz_when_ArraySlice_l159_275 <= _zz_when_ArraySlice_l159_275_2);
  assign _zz_realValue_0_275 = (_zz__zz_realValue_0_275 % _zz__zz_realValue_0_275_1);
  assign when_ArraySlice_l110_275 = (_zz_realValue_0_275 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_275) begin
      realValue_0_275 = (_zz_realValue_0_275_1 - _zz_realValue_0_275);
    end else begin
      realValue_0_275 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_275 = (_zz_when_ArraySlice_l166_275 <= _zz_when_ArraySlice_l166_275_2);
  assign when_ArraySlice_l158_276 = (_zz_when_ArraySlice_l158_276 <= _zz_when_ArraySlice_l158_276_3);
  assign when_ArraySlice_l159_276 = (_zz_when_ArraySlice_l159_276 <= _zz_when_ArraySlice_l159_276_2);
  assign _zz_realValue_0_276 = (_zz__zz_realValue_0_276 % _zz__zz_realValue_0_276_1);
  assign when_ArraySlice_l110_276 = (_zz_realValue_0_276 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_276) begin
      realValue_0_276 = (_zz_realValue_0_276_1 - _zz_realValue_0_276);
    end else begin
      realValue_0_276 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_276 = (_zz_when_ArraySlice_l166_276 <= _zz_when_ArraySlice_l166_276_2);
  assign when_ArraySlice_l158_277 = (_zz_when_ArraySlice_l158_277 <= _zz_when_ArraySlice_l158_277_3);
  assign when_ArraySlice_l159_277 = (_zz_when_ArraySlice_l159_277 <= _zz_when_ArraySlice_l159_277_2);
  assign _zz_realValue_0_277 = (_zz__zz_realValue_0_277 % _zz__zz_realValue_0_277_1);
  assign when_ArraySlice_l110_277 = (_zz_realValue_0_277 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_277) begin
      realValue_0_277 = (_zz_realValue_0_277_1 - _zz_realValue_0_277);
    end else begin
      realValue_0_277 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_277 = (_zz_when_ArraySlice_l166_277 <= _zz_when_ArraySlice_l166_277_2);
  assign when_ArraySlice_l158_278 = (_zz_when_ArraySlice_l158_278 <= _zz_when_ArraySlice_l158_278_3);
  assign when_ArraySlice_l159_278 = (_zz_when_ArraySlice_l159_278 <= _zz_when_ArraySlice_l159_278_2);
  assign _zz_realValue_0_278 = (_zz__zz_realValue_0_278 % _zz__zz_realValue_0_278_1);
  assign when_ArraySlice_l110_278 = (_zz_realValue_0_278 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_278) begin
      realValue_0_278 = (_zz_realValue_0_278_1 - _zz_realValue_0_278);
    end else begin
      realValue_0_278 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_278 = (_zz_when_ArraySlice_l166_278 <= _zz_when_ArraySlice_l166_278_2);
  assign when_ArraySlice_l158_279 = (_zz_when_ArraySlice_l158_279 <= _zz_when_ArraySlice_l158_279_3);
  assign when_ArraySlice_l159_279 = (_zz_when_ArraySlice_l159_279 <= _zz_when_ArraySlice_l159_279_2);
  assign _zz_realValue_0_279 = (_zz__zz_realValue_0_279 % _zz__zz_realValue_0_279_1);
  assign when_ArraySlice_l110_279 = (_zz_realValue_0_279 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_279) begin
      realValue_0_279 = (_zz_realValue_0_279_1 - _zz_realValue_0_279);
    end else begin
      realValue_0_279 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_279 = (_zz_when_ArraySlice_l166_279 <= _zz_when_ArraySlice_l166_279_2);
  assign when_ArraySlice_l314_2 = (! ((((((_zz_when_ArraySlice_l314_2_1 && _zz_when_ArraySlice_l314_2_2) && (holdReadOp_4 == _zz_when_ArraySlice_l314_2_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_2_4 && _zz_when_ArraySlice_l314_2_5) && (debug_4_34 == _zz_when_ArraySlice_l314_2_6)) && (debug_5_34 == 1'b1)) && (debug_6_34 == 1'b1)) && (debug_7_34 == 1'b1))));
  assign outputStreamArrayData_2_fire_12 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l318_2 = ((_zz_when_ArraySlice_l318_2 == 13'h0) && outputStreamArrayData_2_fire_12);
  assign when_ArraySlice_l304_2 = (allowPadding_2 && (_zz_when_ArraySlice_l304_2_1 <= _zz_when_ArraySlice_l304_2_2));
  assign outputStreamArrayData_2_fire_13 = (outputStreamArrayData_2_valid && outputStreamArrayData_2_ready);
  assign when_ArraySlice_l325_2 = (handshakeTimes_2_value == _zz_when_ArraySlice_l325_2_1);
  assign when_ArraySlice_l233_3 = (_zz_when_ArraySlice_l233_3_1 < _zz_when_ArraySlice_l233_3_4);
  assign when_ArraySlice_l234_3 = ((! holdReadOp_3) && (_zz_when_ArraySlice_l234_3_1 != 7'h0));
  assign _zz_outputStreamArrayData_3_valid_1 = (selectReadFifo_3 + _zz__zz_outputStreamArrayData_3_valid_1_1);
  assign _zz_14 = ({127'd0,1'b1} <<< _zz__zz_14);
  assign _zz_io_pop_ready_11 = outputStreamArrayData_3_ready;
  assign when_ArraySlice_l239_3 = (! holdReadOp_3);
  assign outputStreamArrayData_3_fire_7 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l240_3 = ((7'h01 < _zz_when_ArraySlice_l240_3_1) && outputStreamArrayData_3_fire_7);
  assign when_ArraySlice_l241_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l241_3);
  assign when_ArraySlice_l244_3 = (_zz_when_ArraySlice_l244_3 == 13'h0);
  assign outputStreamArrayData_3_fire_8 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l249_3 = ((_zz_when_ArraySlice_l249_3_1 == 7'h01) && outputStreamArrayData_3_fire_8);
  assign when_ArraySlice_l250_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l250_3);
  assign _zz_realValue1_0_33 = (_zz__zz_realValue1_0_33 % _zz__zz_realValue1_0_33_1);
  assign when_ArraySlice_l95_33 = (_zz_realValue1_0_33 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_33) begin
      realValue1_0_33 = (_zz_realValue1_0_33_1 - _zz_realValue1_0_33);
    end else begin
      realValue1_0_33 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_3 = (_zz_when_ArraySlice_l252_3 < _zz_when_ArraySlice_l252_3_2);
  always @(*) begin
    debug_0_35 = 1'b0;
    if(when_ArraySlice_l158_280) begin
      if(when_ArraySlice_l159_280) begin
        debug_0_35 = 1'b1;
      end else begin
        debug_0_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_280) begin
        debug_0_35 = 1'b1;
      end else begin
        debug_0_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_35 = 1'b0;
    if(when_ArraySlice_l158_281) begin
      if(when_ArraySlice_l159_281) begin
        debug_1_35 = 1'b1;
      end else begin
        debug_1_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_281) begin
        debug_1_35 = 1'b1;
      end else begin
        debug_1_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_35 = 1'b0;
    if(when_ArraySlice_l158_282) begin
      if(when_ArraySlice_l159_282) begin
        debug_2_35 = 1'b1;
      end else begin
        debug_2_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_282) begin
        debug_2_35 = 1'b1;
      end else begin
        debug_2_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_35 = 1'b0;
    if(when_ArraySlice_l158_283) begin
      if(when_ArraySlice_l159_283) begin
        debug_3_35 = 1'b1;
      end else begin
        debug_3_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_283) begin
        debug_3_35 = 1'b1;
      end else begin
        debug_3_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_35 = 1'b0;
    if(when_ArraySlice_l158_284) begin
      if(when_ArraySlice_l159_284) begin
        debug_4_35 = 1'b1;
      end else begin
        debug_4_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_284) begin
        debug_4_35 = 1'b1;
      end else begin
        debug_4_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_35 = 1'b0;
    if(when_ArraySlice_l158_285) begin
      if(when_ArraySlice_l159_285) begin
        debug_5_35 = 1'b1;
      end else begin
        debug_5_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_285) begin
        debug_5_35 = 1'b1;
      end else begin
        debug_5_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_35 = 1'b0;
    if(when_ArraySlice_l158_286) begin
      if(when_ArraySlice_l159_286) begin
        debug_6_35 = 1'b1;
      end else begin
        debug_6_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_286) begin
        debug_6_35 = 1'b1;
      end else begin
        debug_6_35 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_35 = 1'b0;
    if(when_ArraySlice_l158_287) begin
      if(when_ArraySlice_l159_287) begin
        debug_7_35 = 1'b1;
      end else begin
        debug_7_35 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_287) begin
        debug_7_35 = 1'b1;
      end else begin
        debug_7_35 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_280 = (_zz_when_ArraySlice_l158_280 <= _zz_when_ArraySlice_l158_280_3);
  assign when_ArraySlice_l159_280 = (_zz_when_ArraySlice_l159_280 <= _zz_when_ArraySlice_l159_280_1);
  assign _zz_realValue_0_280 = (_zz__zz_realValue_0_280 % _zz__zz_realValue_0_280_1);
  assign when_ArraySlice_l110_280 = (_zz_realValue_0_280 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_280) begin
      realValue_0_280 = (_zz_realValue_0_280_1 - _zz_realValue_0_280);
    end else begin
      realValue_0_280 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_280 = (_zz_when_ArraySlice_l166_280 <= _zz_when_ArraySlice_l166_280_1);
  assign when_ArraySlice_l158_281 = (_zz_when_ArraySlice_l158_281 <= _zz_when_ArraySlice_l158_281_3);
  assign when_ArraySlice_l159_281 = (_zz_when_ArraySlice_l159_281 <= _zz_when_ArraySlice_l159_281_2);
  assign _zz_realValue_0_281 = (_zz__zz_realValue_0_281 % _zz__zz_realValue_0_281_1);
  assign when_ArraySlice_l110_281 = (_zz_realValue_0_281 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_281) begin
      realValue_0_281 = (_zz_realValue_0_281_1 - _zz_realValue_0_281);
    end else begin
      realValue_0_281 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_281 = (_zz_when_ArraySlice_l166_281 <= _zz_when_ArraySlice_l166_281_2);
  assign when_ArraySlice_l158_282 = (_zz_when_ArraySlice_l158_282 <= _zz_when_ArraySlice_l158_282_3);
  assign when_ArraySlice_l159_282 = (_zz_when_ArraySlice_l159_282 <= _zz_when_ArraySlice_l159_282_2);
  assign _zz_realValue_0_282 = (_zz__zz_realValue_0_282 % _zz__zz_realValue_0_282_1);
  assign when_ArraySlice_l110_282 = (_zz_realValue_0_282 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_282) begin
      realValue_0_282 = (_zz_realValue_0_282_1 - _zz_realValue_0_282);
    end else begin
      realValue_0_282 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_282 = (_zz_when_ArraySlice_l166_282 <= _zz_when_ArraySlice_l166_282_2);
  assign when_ArraySlice_l158_283 = (_zz_when_ArraySlice_l158_283 <= _zz_when_ArraySlice_l158_283_3);
  assign when_ArraySlice_l159_283 = (_zz_when_ArraySlice_l159_283 <= _zz_when_ArraySlice_l159_283_2);
  assign _zz_realValue_0_283 = (_zz__zz_realValue_0_283 % _zz__zz_realValue_0_283_1);
  assign when_ArraySlice_l110_283 = (_zz_realValue_0_283 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_283) begin
      realValue_0_283 = (_zz_realValue_0_283_1 - _zz_realValue_0_283);
    end else begin
      realValue_0_283 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_283 = (_zz_when_ArraySlice_l166_283 <= _zz_when_ArraySlice_l166_283_2);
  assign when_ArraySlice_l158_284 = (_zz_when_ArraySlice_l158_284 <= _zz_when_ArraySlice_l158_284_3);
  assign when_ArraySlice_l159_284 = (_zz_when_ArraySlice_l159_284 <= _zz_when_ArraySlice_l159_284_2);
  assign _zz_realValue_0_284 = (_zz__zz_realValue_0_284 % _zz__zz_realValue_0_284_1);
  assign when_ArraySlice_l110_284 = (_zz_realValue_0_284 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_284) begin
      realValue_0_284 = (_zz_realValue_0_284_1 - _zz_realValue_0_284);
    end else begin
      realValue_0_284 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_284 = (_zz_when_ArraySlice_l166_284 <= _zz_when_ArraySlice_l166_284_2);
  assign when_ArraySlice_l158_285 = (_zz_when_ArraySlice_l158_285 <= _zz_when_ArraySlice_l158_285_3);
  assign when_ArraySlice_l159_285 = (_zz_when_ArraySlice_l159_285 <= _zz_when_ArraySlice_l159_285_2);
  assign _zz_realValue_0_285 = (_zz__zz_realValue_0_285 % _zz__zz_realValue_0_285_1);
  assign when_ArraySlice_l110_285 = (_zz_realValue_0_285 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_285) begin
      realValue_0_285 = (_zz_realValue_0_285_1 - _zz_realValue_0_285);
    end else begin
      realValue_0_285 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_285 = (_zz_when_ArraySlice_l166_285 <= _zz_when_ArraySlice_l166_285_2);
  assign when_ArraySlice_l158_286 = (_zz_when_ArraySlice_l158_286 <= _zz_when_ArraySlice_l158_286_3);
  assign when_ArraySlice_l159_286 = (_zz_when_ArraySlice_l159_286 <= _zz_when_ArraySlice_l159_286_2);
  assign _zz_realValue_0_286 = (_zz__zz_realValue_0_286 % _zz__zz_realValue_0_286_1);
  assign when_ArraySlice_l110_286 = (_zz_realValue_0_286 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_286) begin
      realValue_0_286 = (_zz_realValue_0_286_1 - _zz_realValue_0_286);
    end else begin
      realValue_0_286 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_286 = (_zz_when_ArraySlice_l166_286 <= _zz_when_ArraySlice_l166_286_2);
  assign when_ArraySlice_l158_287 = (_zz_when_ArraySlice_l158_287 <= _zz_when_ArraySlice_l158_287_3);
  assign when_ArraySlice_l159_287 = (_zz_when_ArraySlice_l159_287 <= _zz_when_ArraySlice_l159_287_2);
  assign _zz_realValue_0_287 = (_zz__zz_realValue_0_287 % _zz__zz_realValue_0_287_1);
  assign when_ArraySlice_l110_287 = (_zz_realValue_0_287 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_287) begin
      realValue_0_287 = (_zz_realValue_0_287_1 - _zz_realValue_0_287);
    end else begin
      realValue_0_287 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_287 = (_zz_when_ArraySlice_l166_287 <= _zz_when_ArraySlice_l166_287_2);
  assign when_ArraySlice_l257_3 = (! ((((((_zz_when_ArraySlice_l257_3_1 && _zz_when_ArraySlice_l257_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l257_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_3_4 && _zz_when_ArraySlice_l257_3_5) && (debug_4_35 == _zz_when_ArraySlice_l257_3_6)) && (debug_5_35 == 1'b1)) && (debug_6_35 == 1'b1)) && (debug_7_35 == 1'b1))));
  assign when_ArraySlice_l260_3 = (_zz_when_ArraySlice_l260_3_1 <= _zz_when_ArraySlice_l260_3_2);
  assign when_ArraySlice_l263_3 = (_zz_when_ArraySlice_l263_3_1 <= _zz_when_ArraySlice_l263_3_2);
  assign when_ArraySlice_l270_3 = (_zz_when_ArraySlice_l270_3 == 13'h0);
  assign when_ArraySlice_l274_3 = (_zz_when_ArraySlice_l274_3_1 == 7'h0);
  assign outputStreamArrayData_3_fire_9 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l275_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l275_3_1) && outputStreamArrayData_3_fire_9);
  assign _zz_realValue1_0_34 = (_zz__zz_realValue1_0_34 % _zz__zz_realValue1_0_34_1);
  assign when_ArraySlice_l95_34 = (_zz_realValue1_0_34 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_34) begin
      realValue1_0_34 = (_zz_realValue1_0_34_1 - _zz_realValue1_0_34);
    end else begin
      realValue1_0_34 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_3 = (_zz_when_ArraySlice_l277_3 < _zz_when_ArraySlice_l277_3_2);
  always @(*) begin
    debug_0_36 = 1'b0;
    if(when_ArraySlice_l158_288) begin
      if(when_ArraySlice_l159_288) begin
        debug_0_36 = 1'b1;
      end else begin
        debug_0_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_288) begin
        debug_0_36 = 1'b1;
      end else begin
        debug_0_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_36 = 1'b0;
    if(when_ArraySlice_l158_289) begin
      if(when_ArraySlice_l159_289) begin
        debug_1_36 = 1'b1;
      end else begin
        debug_1_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_289) begin
        debug_1_36 = 1'b1;
      end else begin
        debug_1_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_36 = 1'b0;
    if(when_ArraySlice_l158_290) begin
      if(when_ArraySlice_l159_290) begin
        debug_2_36 = 1'b1;
      end else begin
        debug_2_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_290) begin
        debug_2_36 = 1'b1;
      end else begin
        debug_2_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_36 = 1'b0;
    if(when_ArraySlice_l158_291) begin
      if(when_ArraySlice_l159_291) begin
        debug_3_36 = 1'b1;
      end else begin
        debug_3_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_291) begin
        debug_3_36 = 1'b1;
      end else begin
        debug_3_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_36 = 1'b0;
    if(when_ArraySlice_l158_292) begin
      if(when_ArraySlice_l159_292) begin
        debug_4_36 = 1'b1;
      end else begin
        debug_4_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_292) begin
        debug_4_36 = 1'b1;
      end else begin
        debug_4_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_36 = 1'b0;
    if(when_ArraySlice_l158_293) begin
      if(when_ArraySlice_l159_293) begin
        debug_5_36 = 1'b1;
      end else begin
        debug_5_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_293) begin
        debug_5_36 = 1'b1;
      end else begin
        debug_5_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_36 = 1'b0;
    if(when_ArraySlice_l158_294) begin
      if(when_ArraySlice_l159_294) begin
        debug_6_36 = 1'b1;
      end else begin
        debug_6_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_294) begin
        debug_6_36 = 1'b1;
      end else begin
        debug_6_36 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_36 = 1'b0;
    if(when_ArraySlice_l158_295) begin
      if(when_ArraySlice_l159_295) begin
        debug_7_36 = 1'b1;
      end else begin
        debug_7_36 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_295) begin
        debug_7_36 = 1'b1;
      end else begin
        debug_7_36 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_288 = (_zz_when_ArraySlice_l158_288 <= _zz_when_ArraySlice_l158_288_3);
  assign when_ArraySlice_l159_288 = (_zz_when_ArraySlice_l159_288 <= _zz_when_ArraySlice_l159_288_1);
  assign _zz_realValue_0_288 = (_zz__zz_realValue_0_288 % _zz__zz_realValue_0_288_1);
  assign when_ArraySlice_l110_288 = (_zz_realValue_0_288 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_288) begin
      realValue_0_288 = (_zz_realValue_0_288_1 - _zz_realValue_0_288);
    end else begin
      realValue_0_288 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_288 = (_zz_when_ArraySlice_l166_288 <= _zz_when_ArraySlice_l166_288_1);
  assign when_ArraySlice_l158_289 = (_zz_when_ArraySlice_l158_289 <= _zz_when_ArraySlice_l158_289_3);
  assign when_ArraySlice_l159_289 = (_zz_when_ArraySlice_l159_289 <= _zz_when_ArraySlice_l159_289_2);
  assign _zz_realValue_0_289 = (_zz__zz_realValue_0_289 % _zz__zz_realValue_0_289_1);
  assign when_ArraySlice_l110_289 = (_zz_realValue_0_289 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_289) begin
      realValue_0_289 = (_zz_realValue_0_289_1 - _zz_realValue_0_289);
    end else begin
      realValue_0_289 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_289 = (_zz_when_ArraySlice_l166_289 <= _zz_when_ArraySlice_l166_289_2);
  assign when_ArraySlice_l158_290 = (_zz_when_ArraySlice_l158_290 <= _zz_when_ArraySlice_l158_290_3);
  assign when_ArraySlice_l159_290 = (_zz_when_ArraySlice_l159_290 <= _zz_when_ArraySlice_l159_290_2);
  assign _zz_realValue_0_290 = (_zz__zz_realValue_0_290 % _zz__zz_realValue_0_290_1);
  assign when_ArraySlice_l110_290 = (_zz_realValue_0_290 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_290) begin
      realValue_0_290 = (_zz_realValue_0_290_1 - _zz_realValue_0_290);
    end else begin
      realValue_0_290 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_290 = (_zz_when_ArraySlice_l166_290 <= _zz_when_ArraySlice_l166_290_2);
  assign when_ArraySlice_l158_291 = (_zz_when_ArraySlice_l158_291 <= _zz_when_ArraySlice_l158_291_3);
  assign when_ArraySlice_l159_291 = (_zz_when_ArraySlice_l159_291 <= _zz_when_ArraySlice_l159_291_2);
  assign _zz_realValue_0_291 = (_zz__zz_realValue_0_291 % _zz__zz_realValue_0_291_1);
  assign when_ArraySlice_l110_291 = (_zz_realValue_0_291 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_291) begin
      realValue_0_291 = (_zz_realValue_0_291_1 - _zz_realValue_0_291);
    end else begin
      realValue_0_291 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_291 = (_zz_when_ArraySlice_l166_291 <= _zz_when_ArraySlice_l166_291_2);
  assign when_ArraySlice_l158_292 = (_zz_when_ArraySlice_l158_292 <= _zz_when_ArraySlice_l158_292_3);
  assign when_ArraySlice_l159_292 = (_zz_when_ArraySlice_l159_292 <= _zz_when_ArraySlice_l159_292_2);
  assign _zz_realValue_0_292 = (_zz__zz_realValue_0_292 % _zz__zz_realValue_0_292_1);
  assign when_ArraySlice_l110_292 = (_zz_realValue_0_292 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_292) begin
      realValue_0_292 = (_zz_realValue_0_292_1 - _zz_realValue_0_292);
    end else begin
      realValue_0_292 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_292 = (_zz_when_ArraySlice_l166_292 <= _zz_when_ArraySlice_l166_292_2);
  assign when_ArraySlice_l158_293 = (_zz_when_ArraySlice_l158_293 <= _zz_when_ArraySlice_l158_293_3);
  assign when_ArraySlice_l159_293 = (_zz_when_ArraySlice_l159_293 <= _zz_when_ArraySlice_l159_293_2);
  assign _zz_realValue_0_293 = (_zz__zz_realValue_0_293 % _zz__zz_realValue_0_293_1);
  assign when_ArraySlice_l110_293 = (_zz_realValue_0_293 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_293) begin
      realValue_0_293 = (_zz_realValue_0_293_1 - _zz_realValue_0_293);
    end else begin
      realValue_0_293 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_293 = (_zz_when_ArraySlice_l166_293 <= _zz_when_ArraySlice_l166_293_2);
  assign when_ArraySlice_l158_294 = (_zz_when_ArraySlice_l158_294 <= _zz_when_ArraySlice_l158_294_3);
  assign when_ArraySlice_l159_294 = (_zz_when_ArraySlice_l159_294 <= _zz_when_ArraySlice_l159_294_2);
  assign _zz_realValue_0_294 = (_zz__zz_realValue_0_294 % _zz__zz_realValue_0_294_1);
  assign when_ArraySlice_l110_294 = (_zz_realValue_0_294 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_294) begin
      realValue_0_294 = (_zz_realValue_0_294_1 - _zz_realValue_0_294);
    end else begin
      realValue_0_294 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_294 = (_zz_when_ArraySlice_l166_294 <= _zz_when_ArraySlice_l166_294_2);
  assign when_ArraySlice_l158_295 = (_zz_when_ArraySlice_l158_295 <= _zz_when_ArraySlice_l158_295_3);
  assign when_ArraySlice_l159_295 = (_zz_when_ArraySlice_l159_295 <= _zz_when_ArraySlice_l159_295_2);
  assign _zz_realValue_0_295 = (_zz__zz_realValue_0_295 % _zz__zz_realValue_0_295_1);
  assign when_ArraySlice_l110_295 = (_zz_realValue_0_295 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_295) begin
      realValue_0_295 = (_zz_realValue_0_295_1 - _zz_realValue_0_295);
    end else begin
      realValue_0_295 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_295 = (_zz_when_ArraySlice_l166_295 <= _zz_when_ArraySlice_l166_295_2);
  assign when_ArraySlice_l282_3 = (! ((((((_zz_when_ArraySlice_l282_3_1 && _zz_when_ArraySlice_l282_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l282_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_3_4 && _zz_when_ArraySlice_l282_3_5) && (debug_4_36 == _zz_when_ArraySlice_l282_3_6)) && (debug_5_36 == 1'b1)) && (debug_6_36 == 1'b1)) && (debug_7_36 == 1'b1))));
  assign when_ArraySlice_l285_3 = (_zz_when_ArraySlice_l285_3_1 <= _zz_when_ArraySlice_l285_3_2);
  assign when_ArraySlice_l288_3 = (_zz_when_ArraySlice_l288_3_1 <= _zz_when_ArraySlice_l288_3_2);
  assign outputStreamArrayData_3_fire_10 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l295_3 = ((_zz_when_ArraySlice_l295_3 == 13'h0) && outputStreamArrayData_3_fire_10);
  assign outputStreamArrayData_3_fire_11 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l306_3 = ((handshakeTimes_3_value == _zz_when_ArraySlice_l306_3) && outputStreamArrayData_3_fire_11);
  assign _zz_realValue1_0_35 = (_zz__zz_realValue1_0_35 % _zz__zz_realValue1_0_35_1);
  assign when_ArraySlice_l95_35 = (_zz_realValue1_0_35 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_35) begin
      realValue1_0_35 = (_zz_realValue1_0_35_1 - _zz_realValue1_0_35);
    end else begin
      realValue1_0_35 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_3 = (_zz_when_ArraySlice_l307_3 < _zz_when_ArraySlice_l307_3_2);
  always @(*) begin
    debug_0_37 = 1'b0;
    if(when_ArraySlice_l158_296) begin
      if(when_ArraySlice_l159_296) begin
        debug_0_37 = 1'b1;
      end else begin
        debug_0_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_296) begin
        debug_0_37 = 1'b1;
      end else begin
        debug_0_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_37 = 1'b0;
    if(when_ArraySlice_l158_297) begin
      if(when_ArraySlice_l159_297) begin
        debug_1_37 = 1'b1;
      end else begin
        debug_1_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_297) begin
        debug_1_37 = 1'b1;
      end else begin
        debug_1_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_37 = 1'b0;
    if(when_ArraySlice_l158_298) begin
      if(when_ArraySlice_l159_298) begin
        debug_2_37 = 1'b1;
      end else begin
        debug_2_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_298) begin
        debug_2_37 = 1'b1;
      end else begin
        debug_2_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_37 = 1'b0;
    if(when_ArraySlice_l158_299) begin
      if(when_ArraySlice_l159_299) begin
        debug_3_37 = 1'b1;
      end else begin
        debug_3_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_299) begin
        debug_3_37 = 1'b1;
      end else begin
        debug_3_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_37 = 1'b0;
    if(when_ArraySlice_l158_300) begin
      if(when_ArraySlice_l159_300) begin
        debug_4_37 = 1'b1;
      end else begin
        debug_4_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_300) begin
        debug_4_37 = 1'b1;
      end else begin
        debug_4_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_37 = 1'b0;
    if(when_ArraySlice_l158_301) begin
      if(when_ArraySlice_l159_301) begin
        debug_5_37 = 1'b1;
      end else begin
        debug_5_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_301) begin
        debug_5_37 = 1'b1;
      end else begin
        debug_5_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_37 = 1'b0;
    if(when_ArraySlice_l158_302) begin
      if(when_ArraySlice_l159_302) begin
        debug_6_37 = 1'b1;
      end else begin
        debug_6_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_302) begin
        debug_6_37 = 1'b1;
      end else begin
        debug_6_37 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_37 = 1'b0;
    if(when_ArraySlice_l158_303) begin
      if(when_ArraySlice_l159_303) begin
        debug_7_37 = 1'b1;
      end else begin
        debug_7_37 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_303) begin
        debug_7_37 = 1'b1;
      end else begin
        debug_7_37 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_296 = (_zz_when_ArraySlice_l158_296 <= _zz_when_ArraySlice_l158_296_3);
  assign when_ArraySlice_l159_296 = (_zz_when_ArraySlice_l159_296 <= _zz_when_ArraySlice_l159_296_1);
  assign _zz_realValue_0_296 = (_zz__zz_realValue_0_296 % _zz__zz_realValue_0_296_1);
  assign when_ArraySlice_l110_296 = (_zz_realValue_0_296 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_296) begin
      realValue_0_296 = (_zz_realValue_0_296_1 - _zz_realValue_0_296);
    end else begin
      realValue_0_296 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_296 = (_zz_when_ArraySlice_l166_296 <= _zz_when_ArraySlice_l166_296_1);
  assign when_ArraySlice_l158_297 = (_zz_when_ArraySlice_l158_297 <= _zz_when_ArraySlice_l158_297_3);
  assign when_ArraySlice_l159_297 = (_zz_when_ArraySlice_l159_297 <= _zz_when_ArraySlice_l159_297_2);
  assign _zz_realValue_0_297 = (_zz__zz_realValue_0_297 % _zz__zz_realValue_0_297_1);
  assign when_ArraySlice_l110_297 = (_zz_realValue_0_297 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_297) begin
      realValue_0_297 = (_zz_realValue_0_297_1 - _zz_realValue_0_297);
    end else begin
      realValue_0_297 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_297 = (_zz_when_ArraySlice_l166_297 <= _zz_when_ArraySlice_l166_297_2);
  assign when_ArraySlice_l158_298 = (_zz_when_ArraySlice_l158_298 <= _zz_when_ArraySlice_l158_298_3);
  assign when_ArraySlice_l159_298 = (_zz_when_ArraySlice_l159_298 <= _zz_when_ArraySlice_l159_298_2);
  assign _zz_realValue_0_298 = (_zz__zz_realValue_0_298 % _zz__zz_realValue_0_298_1);
  assign when_ArraySlice_l110_298 = (_zz_realValue_0_298 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_298) begin
      realValue_0_298 = (_zz_realValue_0_298_1 - _zz_realValue_0_298);
    end else begin
      realValue_0_298 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_298 = (_zz_when_ArraySlice_l166_298 <= _zz_when_ArraySlice_l166_298_2);
  assign when_ArraySlice_l158_299 = (_zz_when_ArraySlice_l158_299 <= _zz_when_ArraySlice_l158_299_3);
  assign when_ArraySlice_l159_299 = (_zz_when_ArraySlice_l159_299 <= _zz_when_ArraySlice_l159_299_2);
  assign _zz_realValue_0_299 = (_zz__zz_realValue_0_299 % _zz__zz_realValue_0_299_1);
  assign when_ArraySlice_l110_299 = (_zz_realValue_0_299 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_299) begin
      realValue_0_299 = (_zz_realValue_0_299_1 - _zz_realValue_0_299);
    end else begin
      realValue_0_299 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_299 = (_zz_when_ArraySlice_l166_299 <= _zz_when_ArraySlice_l166_299_2);
  assign when_ArraySlice_l158_300 = (_zz_when_ArraySlice_l158_300 <= _zz_when_ArraySlice_l158_300_3);
  assign when_ArraySlice_l159_300 = (_zz_when_ArraySlice_l159_300 <= _zz_when_ArraySlice_l159_300_2);
  assign _zz_realValue_0_300 = (_zz__zz_realValue_0_300 % _zz__zz_realValue_0_300_1);
  assign when_ArraySlice_l110_300 = (_zz_realValue_0_300 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_300) begin
      realValue_0_300 = (_zz_realValue_0_300_1 - _zz_realValue_0_300);
    end else begin
      realValue_0_300 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_300 = (_zz_when_ArraySlice_l166_300 <= _zz_when_ArraySlice_l166_300_2);
  assign when_ArraySlice_l158_301 = (_zz_when_ArraySlice_l158_301 <= _zz_when_ArraySlice_l158_301_3);
  assign when_ArraySlice_l159_301 = (_zz_when_ArraySlice_l159_301 <= _zz_when_ArraySlice_l159_301_2);
  assign _zz_realValue_0_301 = (_zz__zz_realValue_0_301 % _zz__zz_realValue_0_301_1);
  assign when_ArraySlice_l110_301 = (_zz_realValue_0_301 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_301) begin
      realValue_0_301 = (_zz_realValue_0_301_1 - _zz_realValue_0_301);
    end else begin
      realValue_0_301 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_301 = (_zz_when_ArraySlice_l166_301 <= _zz_when_ArraySlice_l166_301_2);
  assign when_ArraySlice_l158_302 = (_zz_when_ArraySlice_l158_302 <= _zz_when_ArraySlice_l158_302_3);
  assign when_ArraySlice_l159_302 = (_zz_when_ArraySlice_l159_302 <= _zz_when_ArraySlice_l159_302_2);
  assign _zz_realValue_0_302 = (_zz__zz_realValue_0_302 % _zz__zz_realValue_0_302_1);
  assign when_ArraySlice_l110_302 = (_zz_realValue_0_302 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_302) begin
      realValue_0_302 = (_zz_realValue_0_302_1 - _zz_realValue_0_302);
    end else begin
      realValue_0_302 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_302 = (_zz_when_ArraySlice_l166_302 <= _zz_when_ArraySlice_l166_302_2);
  assign when_ArraySlice_l158_303 = (_zz_when_ArraySlice_l158_303 <= _zz_when_ArraySlice_l158_303_3);
  assign when_ArraySlice_l159_303 = (_zz_when_ArraySlice_l159_303 <= _zz_when_ArraySlice_l159_303_2);
  assign _zz_realValue_0_303 = (_zz__zz_realValue_0_303 % _zz__zz_realValue_0_303_1);
  assign when_ArraySlice_l110_303 = (_zz_realValue_0_303 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_303) begin
      realValue_0_303 = (_zz_realValue_0_303_1 - _zz_realValue_0_303);
    end else begin
      realValue_0_303 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_303 = (_zz_when_ArraySlice_l166_303 <= _zz_when_ArraySlice_l166_303_2);
  assign when_ArraySlice_l314_3 = (! ((((((_zz_when_ArraySlice_l314_3_1 && _zz_when_ArraySlice_l314_3_2) && (holdReadOp_4 == _zz_when_ArraySlice_l314_3_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_3_4 && _zz_when_ArraySlice_l314_3_5) && (debug_4_37 == _zz_when_ArraySlice_l314_3_6)) && (debug_5_37 == 1'b1)) && (debug_6_37 == 1'b1)) && (debug_7_37 == 1'b1))));
  assign outputStreamArrayData_3_fire_12 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l318_3 = ((_zz_when_ArraySlice_l318_3 == 13'h0) && outputStreamArrayData_3_fire_12);
  assign when_ArraySlice_l304_3 = (allowPadding_3 && (_zz_when_ArraySlice_l304_3_1 <= _zz_when_ArraySlice_l304_3_2));
  assign outputStreamArrayData_3_fire_13 = (outputStreamArrayData_3_valid && outputStreamArrayData_3_ready);
  assign when_ArraySlice_l325_3 = (handshakeTimes_3_value == _zz_when_ArraySlice_l325_3);
  assign when_ArraySlice_l233_4 = (_zz_when_ArraySlice_l233_4 < _zz_when_ArraySlice_l233_4_3);
  assign when_ArraySlice_l234_4 = ((! holdReadOp_4) && (_zz_when_ArraySlice_l234_4_1 != 7'h0));
  assign _zz_outputStreamArrayData_4_valid_1 = (selectReadFifo_4 + _zz__zz_outputStreamArrayData_4_valid_1_1);
  assign _zz_15 = ({127'd0,1'b1} <<< _zz__zz_15);
  assign _zz_io_pop_ready_12 = outputStreamArrayData_4_ready;
  assign when_ArraySlice_l239_4 = (! holdReadOp_4);
  assign outputStreamArrayData_4_fire_7 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l240_4 = ((7'h01 < _zz_when_ArraySlice_l240_4_1) && outputStreamArrayData_4_fire_7);
  assign when_ArraySlice_l241_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l241_4);
  assign when_ArraySlice_l244_4 = (_zz_when_ArraySlice_l244_4 == 13'h0);
  assign outputStreamArrayData_4_fire_8 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l249_4 = ((_zz_when_ArraySlice_l249_4_1 == 7'h01) && outputStreamArrayData_4_fire_8);
  assign when_ArraySlice_l250_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l250_4);
  assign _zz_realValue1_0_36 = (_zz__zz_realValue1_0_36 % _zz__zz_realValue1_0_36_1);
  assign when_ArraySlice_l95_36 = (_zz_realValue1_0_36 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_36) begin
      realValue1_0_36 = (_zz_realValue1_0_36_1 - _zz_realValue1_0_36);
    end else begin
      realValue1_0_36 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_4 = (_zz_when_ArraySlice_l252_4 < _zz_when_ArraySlice_l252_4_2);
  always @(*) begin
    debug_0_38 = 1'b0;
    if(when_ArraySlice_l158_304) begin
      if(when_ArraySlice_l159_304) begin
        debug_0_38 = 1'b1;
      end else begin
        debug_0_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_304) begin
        debug_0_38 = 1'b1;
      end else begin
        debug_0_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_38 = 1'b0;
    if(when_ArraySlice_l158_305) begin
      if(when_ArraySlice_l159_305) begin
        debug_1_38 = 1'b1;
      end else begin
        debug_1_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_305) begin
        debug_1_38 = 1'b1;
      end else begin
        debug_1_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_38 = 1'b0;
    if(when_ArraySlice_l158_306) begin
      if(when_ArraySlice_l159_306) begin
        debug_2_38 = 1'b1;
      end else begin
        debug_2_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_306) begin
        debug_2_38 = 1'b1;
      end else begin
        debug_2_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_38 = 1'b0;
    if(when_ArraySlice_l158_307) begin
      if(when_ArraySlice_l159_307) begin
        debug_3_38 = 1'b1;
      end else begin
        debug_3_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_307) begin
        debug_3_38 = 1'b1;
      end else begin
        debug_3_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_38 = 1'b0;
    if(when_ArraySlice_l158_308) begin
      if(when_ArraySlice_l159_308) begin
        debug_4_38 = 1'b1;
      end else begin
        debug_4_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_308) begin
        debug_4_38 = 1'b1;
      end else begin
        debug_4_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_38 = 1'b0;
    if(when_ArraySlice_l158_309) begin
      if(when_ArraySlice_l159_309) begin
        debug_5_38 = 1'b1;
      end else begin
        debug_5_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_309) begin
        debug_5_38 = 1'b1;
      end else begin
        debug_5_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_38 = 1'b0;
    if(when_ArraySlice_l158_310) begin
      if(when_ArraySlice_l159_310) begin
        debug_6_38 = 1'b1;
      end else begin
        debug_6_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_310) begin
        debug_6_38 = 1'b1;
      end else begin
        debug_6_38 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_38 = 1'b0;
    if(when_ArraySlice_l158_311) begin
      if(when_ArraySlice_l159_311) begin
        debug_7_38 = 1'b1;
      end else begin
        debug_7_38 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_311) begin
        debug_7_38 = 1'b1;
      end else begin
        debug_7_38 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_304 = (_zz_when_ArraySlice_l158_304 <= _zz_when_ArraySlice_l158_304_3);
  assign when_ArraySlice_l159_304 = (_zz_when_ArraySlice_l159_304 <= _zz_when_ArraySlice_l159_304_1);
  assign _zz_realValue_0_304 = (_zz__zz_realValue_0_304 % _zz__zz_realValue_0_304_1);
  assign when_ArraySlice_l110_304 = (_zz_realValue_0_304 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_304) begin
      realValue_0_304 = (_zz_realValue_0_304_1 - _zz_realValue_0_304);
    end else begin
      realValue_0_304 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_304 = (_zz_when_ArraySlice_l166_304 <= _zz_when_ArraySlice_l166_304_1);
  assign when_ArraySlice_l158_305 = (_zz_when_ArraySlice_l158_305 <= _zz_when_ArraySlice_l158_305_3);
  assign when_ArraySlice_l159_305 = (_zz_when_ArraySlice_l159_305 <= _zz_when_ArraySlice_l159_305_2);
  assign _zz_realValue_0_305 = (_zz__zz_realValue_0_305 % _zz__zz_realValue_0_305_1);
  assign when_ArraySlice_l110_305 = (_zz_realValue_0_305 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_305) begin
      realValue_0_305 = (_zz_realValue_0_305_1 - _zz_realValue_0_305);
    end else begin
      realValue_0_305 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_305 = (_zz_when_ArraySlice_l166_305 <= _zz_when_ArraySlice_l166_305_2);
  assign when_ArraySlice_l158_306 = (_zz_when_ArraySlice_l158_306 <= _zz_when_ArraySlice_l158_306_3);
  assign when_ArraySlice_l159_306 = (_zz_when_ArraySlice_l159_306 <= _zz_when_ArraySlice_l159_306_2);
  assign _zz_realValue_0_306 = (_zz__zz_realValue_0_306 % _zz__zz_realValue_0_306_1);
  assign when_ArraySlice_l110_306 = (_zz_realValue_0_306 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_306) begin
      realValue_0_306 = (_zz_realValue_0_306_1 - _zz_realValue_0_306);
    end else begin
      realValue_0_306 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_306 = (_zz_when_ArraySlice_l166_306 <= _zz_when_ArraySlice_l166_306_2);
  assign when_ArraySlice_l158_307 = (_zz_when_ArraySlice_l158_307 <= _zz_when_ArraySlice_l158_307_3);
  assign when_ArraySlice_l159_307 = (_zz_when_ArraySlice_l159_307 <= _zz_when_ArraySlice_l159_307_2);
  assign _zz_realValue_0_307 = (_zz__zz_realValue_0_307 % _zz__zz_realValue_0_307_1);
  assign when_ArraySlice_l110_307 = (_zz_realValue_0_307 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_307) begin
      realValue_0_307 = (_zz_realValue_0_307_1 - _zz_realValue_0_307);
    end else begin
      realValue_0_307 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_307 = (_zz_when_ArraySlice_l166_307 <= _zz_when_ArraySlice_l166_307_2);
  assign when_ArraySlice_l158_308 = (_zz_when_ArraySlice_l158_308 <= _zz_when_ArraySlice_l158_308_3);
  assign when_ArraySlice_l159_308 = (_zz_when_ArraySlice_l159_308 <= _zz_when_ArraySlice_l159_308_2);
  assign _zz_realValue_0_308 = (_zz__zz_realValue_0_308 % _zz__zz_realValue_0_308_1);
  assign when_ArraySlice_l110_308 = (_zz_realValue_0_308 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_308) begin
      realValue_0_308 = (_zz_realValue_0_308_1 - _zz_realValue_0_308);
    end else begin
      realValue_0_308 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_308 = (_zz_when_ArraySlice_l166_308 <= _zz_when_ArraySlice_l166_308_2);
  assign when_ArraySlice_l158_309 = (_zz_when_ArraySlice_l158_309 <= _zz_when_ArraySlice_l158_309_3);
  assign when_ArraySlice_l159_309 = (_zz_when_ArraySlice_l159_309 <= _zz_when_ArraySlice_l159_309_2);
  assign _zz_realValue_0_309 = (_zz__zz_realValue_0_309 % _zz__zz_realValue_0_309_1);
  assign when_ArraySlice_l110_309 = (_zz_realValue_0_309 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_309) begin
      realValue_0_309 = (_zz_realValue_0_309_1 - _zz_realValue_0_309);
    end else begin
      realValue_0_309 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_309 = (_zz_when_ArraySlice_l166_309 <= _zz_when_ArraySlice_l166_309_2);
  assign when_ArraySlice_l158_310 = (_zz_when_ArraySlice_l158_310 <= _zz_when_ArraySlice_l158_310_3);
  assign when_ArraySlice_l159_310 = (_zz_when_ArraySlice_l159_310 <= _zz_when_ArraySlice_l159_310_2);
  assign _zz_realValue_0_310 = (_zz__zz_realValue_0_310 % _zz__zz_realValue_0_310_1);
  assign when_ArraySlice_l110_310 = (_zz_realValue_0_310 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_310) begin
      realValue_0_310 = (_zz_realValue_0_310_1 - _zz_realValue_0_310);
    end else begin
      realValue_0_310 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_310 = (_zz_when_ArraySlice_l166_310 <= _zz_when_ArraySlice_l166_310_2);
  assign when_ArraySlice_l158_311 = (_zz_when_ArraySlice_l158_311 <= _zz_when_ArraySlice_l158_311_3);
  assign when_ArraySlice_l159_311 = (_zz_when_ArraySlice_l159_311 <= _zz_when_ArraySlice_l159_311_2);
  assign _zz_realValue_0_311 = (_zz__zz_realValue_0_311 % _zz__zz_realValue_0_311_1);
  assign when_ArraySlice_l110_311 = (_zz_realValue_0_311 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_311) begin
      realValue_0_311 = (_zz_realValue_0_311_1 - _zz_realValue_0_311);
    end else begin
      realValue_0_311 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_311 = (_zz_when_ArraySlice_l166_311 <= _zz_when_ArraySlice_l166_311_2);
  assign when_ArraySlice_l257_4 = (! ((((((_zz_when_ArraySlice_l257_4_1 && _zz_when_ArraySlice_l257_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l257_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_4_4 && _zz_when_ArraySlice_l257_4_5) && (debug_4_38 == _zz_when_ArraySlice_l257_4_6)) && (debug_5_38 == 1'b1)) && (debug_6_38 == 1'b1)) && (debug_7_38 == 1'b1))));
  assign when_ArraySlice_l260_4 = (_zz_when_ArraySlice_l260_4_1 <= _zz_when_ArraySlice_l260_4_2);
  assign when_ArraySlice_l263_4 = (_zz_when_ArraySlice_l263_4_1 <= _zz_when_ArraySlice_l263_4_2);
  assign when_ArraySlice_l270_4 = (_zz_when_ArraySlice_l270_4 == 13'h0);
  assign when_ArraySlice_l274_4 = (_zz_when_ArraySlice_l274_4_1 == 7'h0);
  assign outputStreamArrayData_4_fire_9 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l275_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l275_4_1) && outputStreamArrayData_4_fire_9);
  assign _zz_realValue1_0_37 = (_zz__zz_realValue1_0_37 % _zz__zz_realValue1_0_37_1);
  assign when_ArraySlice_l95_37 = (_zz_realValue1_0_37 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_37) begin
      realValue1_0_37 = (_zz_realValue1_0_37_1 - _zz_realValue1_0_37);
    end else begin
      realValue1_0_37 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_4 = (_zz_when_ArraySlice_l277_4 < _zz_when_ArraySlice_l277_4_2);
  always @(*) begin
    debug_0_39 = 1'b0;
    if(when_ArraySlice_l158_312) begin
      if(when_ArraySlice_l159_312) begin
        debug_0_39 = 1'b1;
      end else begin
        debug_0_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_312) begin
        debug_0_39 = 1'b1;
      end else begin
        debug_0_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_39 = 1'b0;
    if(when_ArraySlice_l158_313) begin
      if(when_ArraySlice_l159_313) begin
        debug_1_39 = 1'b1;
      end else begin
        debug_1_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_313) begin
        debug_1_39 = 1'b1;
      end else begin
        debug_1_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_39 = 1'b0;
    if(when_ArraySlice_l158_314) begin
      if(when_ArraySlice_l159_314) begin
        debug_2_39 = 1'b1;
      end else begin
        debug_2_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_314) begin
        debug_2_39 = 1'b1;
      end else begin
        debug_2_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_39 = 1'b0;
    if(when_ArraySlice_l158_315) begin
      if(when_ArraySlice_l159_315) begin
        debug_3_39 = 1'b1;
      end else begin
        debug_3_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_315) begin
        debug_3_39 = 1'b1;
      end else begin
        debug_3_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_39 = 1'b0;
    if(when_ArraySlice_l158_316) begin
      if(when_ArraySlice_l159_316) begin
        debug_4_39 = 1'b1;
      end else begin
        debug_4_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_316) begin
        debug_4_39 = 1'b1;
      end else begin
        debug_4_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_39 = 1'b0;
    if(when_ArraySlice_l158_317) begin
      if(when_ArraySlice_l159_317) begin
        debug_5_39 = 1'b1;
      end else begin
        debug_5_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_317) begin
        debug_5_39 = 1'b1;
      end else begin
        debug_5_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_39 = 1'b0;
    if(when_ArraySlice_l158_318) begin
      if(when_ArraySlice_l159_318) begin
        debug_6_39 = 1'b1;
      end else begin
        debug_6_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_318) begin
        debug_6_39 = 1'b1;
      end else begin
        debug_6_39 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_39 = 1'b0;
    if(when_ArraySlice_l158_319) begin
      if(when_ArraySlice_l159_319) begin
        debug_7_39 = 1'b1;
      end else begin
        debug_7_39 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_319) begin
        debug_7_39 = 1'b1;
      end else begin
        debug_7_39 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_312 = (_zz_when_ArraySlice_l158_312 <= _zz_when_ArraySlice_l158_312_3);
  assign when_ArraySlice_l159_312 = (_zz_when_ArraySlice_l159_312 <= _zz_when_ArraySlice_l159_312_1);
  assign _zz_realValue_0_312 = (_zz__zz_realValue_0_312 % _zz__zz_realValue_0_312_1);
  assign when_ArraySlice_l110_312 = (_zz_realValue_0_312 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_312) begin
      realValue_0_312 = (_zz_realValue_0_312_1 - _zz_realValue_0_312);
    end else begin
      realValue_0_312 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_312 = (_zz_when_ArraySlice_l166_312 <= _zz_when_ArraySlice_l166_312_1);
  assign when_ArraySlice_l158_313 = (_zz_when_ArraySlice_l158_313 <= _zz_when_ArraySlice_l158_313_3);
  assign when_ArraySlice_l159_313 = (_zz_when_ArraySlice_l159_313 <= _zz_when_ArraySlice_l159_313_2);
  assign _zz_realValue_0_313 = (_zz__zz_realValue_0_313 % _zz__zz_realValue_0_313_1);
  assign when_ArraySlice_l110_313 = (_zz_realValue_0_313 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_313) begin
      realValue_0_313 = (_zz_realValue_0_313_1 - _zz_realValue_0_313);
    end else begin
      realValue_0_313 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_313 = (_zz_when_ArraySlice_l166_313 <= _zz_when_ArraySlice_l166_313_2);
  assign when_ArraySlice_l158_314 = (_zz_when_ArraySlice_l158_314 <= _zz_when_ArraySlice_l158_314_3);
  assign when_ArraySlice_l159_314 = (_zz_when_ArraySlice_l159_314 <= _zz_when_ArraySlice_l159_314_2);
  assign _zz_realValue_0_314 = (_zz__zz_realValue_0_314 % _zz__zz_realValue_0_314_1);
  assign when_ArraySlice_l110_314 = (_zz_realValue_0_314 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_314) begin
      realValue_0_314 = (_zz_realValue_0_314_1 - _zz_realValue_0_314);
    end else begin
      realValue_0_314 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_314 = (_zz_when_ArraySlice_l166_314 <= _zz_when_ArraySlice_l166_314_2);
  assign when_ArraySlice_l158_315 = (_zz_when_ArraySlice_l158_315 <= _zz_when_ArraySlice_l158_315_3);
  assign when_ArraySlice_l159_315 = (_zz_when_ArraySlice_l159_315 <= _zz_when_ArraySlice_l159_315_2);
  assign _zz_realValue_0_315 = (_zz__zz_realValue_0_315 % _zz__zz_realValue_0_315_1);
  assign when_ArraySlice_l110_315 = (_zz_realValue_0_315 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_315) begin
      realValue_0_315 = (_zz_realValue_0_315_1 - _zz_realValue_0_315);
    end else begin
      realValue_0_315 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_315 = (_zz_when_ArraySlice_l166_315 <= _zz_when_ArraySlice_l166_315_2);
  assign when_ArraySlice_l158_316 = (_zz_when_ArraySlice_l158_316 <= _zz_when_ArraySlice_l158_316_3);
  assign when_ArraySlice_l159_316 = (_zz_when_ArraySlice_l159_316 <= _zz_when_ArraySlice_l159_316_2);
  assign _zz_realValue_0_316 = (_zz__zz_realValue_0_316 % _zz__zz_realValue_0_316_1);
  assign when_ArraySlice_l110_316 = (_zz_realValue_0_316 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_316) begin
      realValue_0_316 = (_zz_realValue_0_316_1 - _zz_realValue_0_316);
    end else begin
      realValue_0_316 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_316 = (_zz_when_ArraySlice_l166_316 <= _zz_when_ArraySlice_l166_316_2);
  assign when_ArraySlice_l158_317 = (_zz_when_ArraySlice_l158_317 <= _zz_when_ArraySlice_l158_317_3);
  assign when_ArraySlice_l159_317 = (_zz_when_ArraySlice_l159_317 <= _zz_when_ArraySlice_l159_317_2);
  assign _zz_realValue_0_317 = (_zz__zz_realValue_0_317 % _zz__zz_realValue_0_317_1);
  assign when_ArraySlice_l110_317 = (_zz_realValue_0_317 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_317) begin
      realValue_0_317 = (_zz_realValue_0_317_1 - _zz_realValue_0_317);
    end else begin
      realValue_0_317 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_317 = (_zz_when_ArraySlice_l166_317 <= _zz_when_ArraySlice_l166_317_2);
  assign when_ArraySlice_l158_318 = (_zz_when_ArraySlice_l158_318 <= _zz_when_ArraySlice_l158_318_3);
  assign when_ArraySlice_l159_318 = (_zz_when_ArraySlice_l159_318 <= _zz_when_ArraySlice_l159_318_2);
  assign _zz_realValue_0_318 = (_zz__zz_realValue_0_318 % _zz__zz_realValue_0_318_1);
  assign when_ArraySlice_l110_318 = (_zz_realValue_0_318 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_318) begin
      realValue_0_318 = (_zz_realValue_0_318_1 - _zz_realValue_0_318);
    end else begin
      realValue_0_318 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_318 = (_zz_when_ArraySlice_l166_318 <= _zz_when_ArraySlice_l166_318_2);
  assign when_ArraySlice_l158_319 = (_zz_when_ArraySlice_l158_319 <= _zz_when_ArraySlice_l158_319_3);
  assign when_ArraySlice_l159_319 = (_zz_when_ArraySlice_l159_319 <= _zz_when_ArraySlice_l159_319_2);
  assign _zz_realValue_0_319 = (_zz__zz_realValue_0_319 % _zz__zz_realValue_0_319_1);
  assign when_ArraySlice_l110_319 = (_zz_realValue_0_319 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_319) begin
      realValue_0_319 = (_zz_realValue_0_319_1 - _zz_realValue_0_319);
    end else begin
      realValue_0_319 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_319 = (_zz_when_ArraySlice_l166_319 <= _zz_when_ArraySlice_l166_319_2);
  assign when_ArraySlice_l282_4 = (! ((((((_zz_when_ArraySlice_l282_4_1 && _zz_when_ArraySlice_l282_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l282_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_4_4 && _zz_when_ArraySlice_l282_4_5) && (debug_4_39 == _zz_when_ArraySlice_l282_4_6)) && (debug_5_39 == 1'b1)) && (debug_6_39 == 1'b1)) && (debug_7_39 == 1'b1))));
  assign when_ArraySlice_l285_4 = (_zz_when_ArraySlice_l285_4_1 <= _zz_when_ArraySlice_l285_4_2);
  assign when_ArraySlice_l288_4 = (_zz_when_ArraySlice_l288_4_1 <= _zz_when_ArraySlice_l288_4_2);
  assign outputStreamArrayData_4_fire_10 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l295_4 = ((_zz_when_ArraySlice_l295_4 == 13'h0) && outputStreamArrayData_4_fire_10);
  assign outputStreamArrayData_4_fire_11 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l306_4 = ((handshakeTimes_4_value == _zz_when_ArraySlice_l306_4) && outputStreamArrayData_4_fire_11);
  assign _zz_realValue1_0_38 = (_zz__zz_realValue1_0_38 % _zz__zz_realValue1_0_38_1);
  assign when_ArraySlice_l95_38 = (_zz_realValue1_0_38 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_38) begin
      realValue1_0_38 = (_zz_realValue1_0_38_1 - _zz_realValue1_0_38);
    end else begin
      realValue1_0_38 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_4 = (_zz_when_ArraySlice_l307_4 < _zz_when_ArraySlice_l307_4_2);
  always @(*) begin
    debug_0_40 = 1'b0;
    if(when_ArraySlice_l158_320) begin
      if(when_ArraySlice_l159_320) begin
        debug_0_40 = 1'b1;
      end else begin
        debug_0_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_320) begin
        debug_0_40 = 1'b1;
      end else begin
        debug_0_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_40 = 1'b0;
    if(when_ArraySlice_l158_321) begin
      if(when_ArraySlice_l159_321) begin
        debug_1_40 = 1'b1;
      end else begin
        debug_1_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_321) begin
        debug_1_40 = 1'b1;
      end else begin
        debug_1_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_40 = 1'b0;
    if(when_ArraySlice_l158_322) begin
      if(when_ArraySlice_l159_322) begin
        debug_2_40 = 1'b1;
      end else begin
        debug_2_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_322) begin
        debug_2_40 = 1'b1;
      end else begin
        debug_2_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_40 = 1'b0;
    if(when_ArraySlice_l158_323) begin
      if(when_ArraySlice_l159_323) begin
        debug_3_40 = 1'b1;
      end else begin
        debug_3_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_323) begin
        debug_3_40 = 1'b1;
      end else begin
        debug_3_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_40 = 1'b0;
    if(when_ArraySlice_l158_324) begin
      if(when_ArraySlice_l159_324) begin
        debug_4_40 = 1'b1;
      end else begin
        debug_4_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_324) begin
        debug_4_40 = 1'b1;
      end else begin
        debug_4_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_40 = 1'b0;
    if(when_ArraySlice_l158_325) begin
      if(when_ArraySlice_l159_325) begin
        debug_5_40 = 1'b1;
      end else begin
        debug_5_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_325) begin
        debug_5_40 = 1'b1;
      end else begin
        debug_5_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_40 = 1'b0;
    if(when_ArraySlice_l158_326) begin
      if(when_ArraySlice_l159_326) begin
        debug_6_40 = 1'b1;
      end else begin
        debug_6_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_326) begin
        debug_6_40 = 1'b1;
      end else begin
        debug_6_40 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_40 = 1'b0;
    if(when_ArraySlice_l158_327) begin
      if(when_ArraySlice_l159_327) begin
        debug_7_40 = 1'b1;
      end else begin
        debug_7_40 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_327) begin
        debug_7_40 = 1'b1;
      end else begin
        debug_7_40 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_320 = (_zz_when_ArraySlice_l158_320 <= _zz_when_ArraySlice_l158_320_3);
  assign when_ArraySlice_l159_320 = (_zz_when_ArraySlice_l159_320 <= _zz_when_ArraySlice_l159_320_1);
  assign _zz_realValue_0_320 = (_zz__zz_realValue_0_320 % _zz__zz_realValue_0_320_1);
  assign when_ArraySlice_l110_320 = (_zz_realValue_0_320 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_320) begin
      realValue_0_320 = (_zz_realValue_0_320_1 - _zz_realValue_0_320);
    end else begin
      realValue_0_320 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_320 = (_zz_when_ArraySlice_l166_320 <= _zz_when_ArraySlice_l166_320_1);
  assign when_ArraySlice_l158_321 = (_zz_when_ArraySlice_l158_321 <= _zz_when_ArraySlice_l158_321_3);
  assign when_ArraySlice_l159_321 = (_zz_when_ArraySlice_l159_321 <= _zz_when_ArraySlice_l159_321_2);
  assign _zz_realValue_0_321 = (_zz__zz_realValue_0_321 % _zz__zz_realValue_0_321_1);
  assign when_ArraySlice_l110_321 = (_zz_realValue_0_321 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_321) begin
      realValue_0_321 = (_zz_realValue_0_321_1 - _zz_realValue_0_321);
    end else begin
      realValue_0_321 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_321 = (_zz_when_ArraySlice_l166_321 <= _zz_when_ArraySlice_l166_321_2);
  assign when_ArraySlice_l158_322 = (_zz_when_ArraySlice_l158_322 <= _zz_when_ArraySlice_l158_322_3);
  assign when_ArraySlice_l159_322 = (_zz_when_ArraySlice_l159_322 <= _zz_when_ArraySlice_l159_322_2);
  assign _zz_realValue_0_322 = (_zz__zz_realValue_0_322 % _zz__zz_realValue_0_322_1);
  assign when_ArraySlice_l110_322 = (_zz_realValue_0_322 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_322) begin
      realValue_0_322 = (_zz_realValue_0_322_1 - _zz_realValue_0_322);
    end else begin
      realValue_0_322 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_322 = (_zz_when_ArraySlice_l166_322 <= _zz_when_ArraySlice_l166_322_2);
  assign when_ArraySlice_l158_323 = (_zz_when_ArraySlice_l158_323 <= _zz_when_ArraySlice_l158_323_3);
  assign when_ArraySlice_l159_323 = (_zz_when_ArraySlice_l159_323 <= _zz_when_ArraySlice_l159_323_2);
  assign _zz_realValue_0_323 = (_zz__zz_realValue_0_323 % _zz__zz_realValue_0_323_1);
  assign when_ArraySlice_l110_323 = (_zz_realValue_0_323 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_323) begin
      realValue_0_323 = (_zz_realValue_0_323_1 - _zz_realValue_0_323);
    end else begin
      realValue_0_323 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_323 = (_zz_when_ArraySlice_l166_323 <= _zz_when_ArraySlice_l166_323_2);
  assign when_ArraySlice_l158_324 = (_zz_when_ArraySlice_l158_324 <= _zz_when_ArraySlice_l158_324_3);
  assign when_ArraySlice_l159_324 = (_zz_when_ArraySlice_l159_324 <= _zz_when_ArraySlice_l159_324_2);
  assign _zz_realValue_0_324 = (_zz__zz_realValue_0_324 % _zz__zz_realValue_0_324_1);
  assign when_ArraySlice_l110_324 = (_zz_realValue_0_324 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_324) begin
      realValue_0_324 = (_zz_realValue_0_324_1 - _zz_realValue_0_324);
    end else begin
      realValue_0_324 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_324 = (_zz_when_ArraySlice_l166_324 <= _zz_when_ArraySlice_l166_324_2);
  assign when_ArraySlice_l158_325 = (_zz_when_ArraySlice_l158_325 <= _zz_when_ArraySlice_l158_325_3);
  assign when_ArraySlice_l159_325 = (_zz_when_ArraySlice_l159_325 <= _zz_when_ArraySlice_l159_325_2);
  assign _zz_realValue_0_325 = (_zz__zz_realValue_0_325 % _zz__zz_realValue_0_325_1);
  assign when_ArraySlice_l110_325 = (_zz_realValue_0_325 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_325) begin
      realValue_0_325 = (_zz_realValue_0_325_1 - _zz_realValue_0_325);
    end else begin
      realValue_0_325 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_325 = (_zz_when_ArraySlice_l166_325 <= _zz_when_ArraySlice_l166_325_2);
  assign when_ArraySlice_l158_326 = (_zz_when_ArraySlice_l158_326 <= _zz_when_ArraySlice_l158_326_3);
  assign when_ArraySlice_l159_326 = (_zz_when_ArraySlice_l159_326 <= _zz_when_ArraySlice_l159_326_2);
  assign _zz_realValue_0_326 = (_zz__zz_realValue_0_326 % _zz__zz_realValue_0_326_1);
  assign when_ArraySlice_l110_326 = (_zz_realValue_0_326 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_326) begin
      realValue_0_326 = (_zz_realValue_0_326_1 - _zz_realValue_0_326);
    end else begin
      realValue_0_326 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_326 = (_zz_when_ArraySlice_l166_326 <= _zz_when_ArraySlice_l166_326_2);
  assign when_ArraySlice_l158_327 = (_zz_when_ArraySlice_l158_327 <= _zz_when_ArraySlice_l158_327_3);
  assign when_ArraySlice_l159_327 = (_zz_when_ArraySlice_l159_327 <= _zz_when_ArraySlice_l159_327_2);
  assign _zz_realValue_0_327 = (_zz__zz_realValue_0_327 % _zz__zz_realValue_0_327_1);
  assign when_ArraySlice_l110_327 = (_zz_realValue_0_327 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_327) begin
      realValue_0_327 = (_zz_realValue_0_327_1 - _zz_realValue_0_327);
    end else begin
      realValue_0_327 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_327 = (_zz_when_ArraySlice_l166_327 <= _zz_when_ArraySlice_l166_327_2);
  assign when_ArraySlice_l314_4 = (! ((((((_zz_when_ArraySlice_l314_4_1 && _zz_when_ArraySlice_l314_4_2) && (holdReadOp_4 == _zz_when_ArraySlice_l314_4_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_4_4 && _zz_when_ArraySlice_l314_4_5) && (debug_4_40 == _zz_when_ArraySlice_l314_4_6)) && (debug_5_40 == 1'b1)) && (debug_6_40 == 1'b1)) && (debug_7_40 == 1'b1))));
  assign outputStreamArrayData_4_fire_12 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l318_4 = ((_zz_when_ArraySlice_l318_4 == 13'h0) && outputStreamArrayData_4_fire_12);
  assign when_ArraySlice_l304_4 = (allowPadding_4 && (_zz_when_ArraySlice_l304_4 <= _zz_when_ArraySlice_l304_4_1));
  assign outputStreamArrayData_4_fire_13 = (outputStreamArrayData_4_valid && outputStreamArrayData_4_ready);
  assign when_ArraySlice_l325_4 = (handshakeTimes_4_value == _zz_when_ArraySlice_l325_4);
  assign when_ArraySlice_l233_5 = (_zz_when_ArraySlice_l233_5 < _zz_when_ArraySlice_l233_5_3);
  assign when_ArraySlice_l234_5 = ((! holdReadOp_5) && (_zz_when_ArraySlice_l234_5 != 7'h0));
  assign _zz_outputStreamArrayData_5_valid_1 = (selectReadFifo_5 + _zz__zz_outputStreamArrayData_5_valid_1_1);
  assign _zz_16 = ({127'd0,1'b1} <<< _zz__zz_16);
  assign _zz_io_pop_ready_13 = outputStreamArrayData_5_ready;
  assign when_ArraySlice_l239_5 = (! holdReadOp_5);
  assign outputStreamArrayData_5_fire_7 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l240_5 = ((7'h01 < _zz_when_ArraySlice_l240_5) && outputStreamArrayData_5_fire_7);
  assign when_ArraySlice_l241_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l241_5);
  assign when_ArraySlice_l244_5 = (_zz_when_ArraySlice_l244_5 == 13'h0);
  assign outputStreamArrayData_5_fire_8 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l249_5 = ((_zz_when_ArraySlice_l249_5 == 7'h01) && outputStreamArrayData_5_fire_8);
  assign when_ArraySlice_l250_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l250_5);
  assign _zz_realValue1_0_39 = (_zz__zz_realValue1_0_39 % _zz__zz_realValue1_0_39_1);
  assign when_ArraySlice_l95_39 = (_zz_realValue1_0_39 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_39) begin
      realValue1_0_39 = (_zz_realValue1_0_39_1 - _zz_realValue1_0_39);
    end else begin
      realValue1_0_39 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_5 = (_zz_when_ArraySlice_l252_5 < _zz_when_ArraySlice_l252_5_2);
  always @(*) begin
    debug_0_41 = 1'b0;
    if(when_ArraySlice_l158_328) begin
      if(when_ArraySlice_l159_328) begin
        debug_0_41 = 1'b1;
      end else begin
        debug_0_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_328) begin
        debug_0_41 = 1'b1;
      end else begin
        debug_0_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_41 = 1'b0;
    if(when_ArraySlice_l158_329) begin
      if(when_ArraySlice_l159_329) begin
        debug_1_41 = 1'b1;
      end else begin
        debug_1_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_329) begin
        debug_1_41 = 1'b1;
      end else begin
        debug_1_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_41 = 1'b0;
    if(when_ArraySlice_l158_330) begin
      if(when_ArraySlice_l159_330) begin
        debug_2_41 = 1'b1;
      end else begin
        debug_2_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_330) begin
        debug_2_41 = 1'b1;
      end else begin
        debug_2_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_41 = 1'b0;
    if(when_ArraySlice_l158_331) begin
      if(when_ArraySlice_l159_331) begin
        debug_3_41 = 1'b1;
      end else begin
        debug_3_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_331) begin
        debug_3_41 = 1'b1;
      end else begin
        debug_3_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_41 = 1'b0;
    if(when_ArraySlice_l158_332) begin
      if(when_ArraySlice_l159_332) begin
        debug_4_41 = 1'b1;
      end else begin
        debug_4_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_332) begin
        debug_4_41 = 1'b1;
      end else begin
        debug_4_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_41 = 1'b0;
    if(when_ArraySlice_l158_333) begin
      if(when_ArraySlice_l159_333) begin
        debug_5_41 = 1'b1;
      end else begin
        debug_5_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_333) begin
        debug_5_41 = 1'b1;
      end else begin
        debug_5_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_41 = 1'b0;
    if(when_ArraySlice_l158_334) begin
      if(when_ArraySlice_l159_334) begin
        debug_6_41 = 1'b1;
      end else begin
        debug_6_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_334) begin
        debug_6_41 = 1'b1;
      end else begin
        debug_6_41 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_41 = 1'b0;
    if(when_ArraySlice_l158_335) begin
      if(when_ArraySlice_l159_335) begin
        debug_7_41 = 1'b1;
      end else begin
        debug_7_41 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_335) begin
        debug_7_41 = 1'b1;
      end else begin
        debug_7_41 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_328 = (_zz_when_ArraySlice_l158_328 <= _zz_when_ArraySlice_l158_328_3);
  assign when_ArraySlice_l159_328 = (_zz_when_ArraySlice_l159_328 <= _zz_when_ArraySlice_l159_328_1);
  assign _zz_realValue_0_328 = (_zz__zz_realValue_0_328 % _zz__zz_realValue_0_328_1);
  assign when_ArraySlice_l110_328 = (_zz_realValue_0_328 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_328) begin
      realValue_0_328 = (_zz_realValue_0_328_1 - _zz_realValue_0_328);
    end else begin
      realValue_0_328 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_328 = (_zz_when_ArraySlice_l166_328 <= _zz_when_ArraySlice_l166_328_1);
  assign when_ArraySlice_l158_329 = (_zz_when_ArraySlice_l158_329 <= _zz_when_ArraySlice_l158_329_3);
  assign when_ArraySlice_l159_329 = (_zz_when_ArraySlice_l159_329 <= _zz_when_ArraySlice_l159_329_2);
  assign _zz_realValue_0_329 = (_zz__zz_realValue_0_329 % _zz__zz_realValue_0_329_1);
  assign when_ArraySlice_l110_329 = (_zz_realValue_0_329 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_329) begin
      realValue_0_329 = (_zz_realValue_0_329_1 - _zz_realValue_0_329);
    end else begin
      realValue_0_329 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_329 = (_zz_when_ArraySlice_l166_329 <= _zz_when_ArraySlice_l166_329_2);
  assign when_ArraySlice_l158_330 = (_zz_when_ArraySlice_l158_330 <= _zz_when_ArraySlice_l158_330_3);
  assign when_ArraySlice_l159_330 = (_zz_when_ArraySlice_l159_330 <= _zz_when_ArraySlice_l159_330_2);
  assign _zz_realValue_0_330 = (_zz__zz_realValue_0_330 % _zz__zz_realValue_0_330_1);
  assign when_ArraySlice_l110_330 = (_zz_realValue_0_330 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_330) begin
      realValue_0_330 = (_zz_realValue_0_330_1 - _zz_realValue_0_330);
    end else begin
      realValue_0_330 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_330 = (_zz_when_ArraySlice_l166_330 <= _zz_when_ArraySlice_l166_330_2);
  assign when_ArraySlice_l158_331 = (_zz_when_ArraySlice_l158_331 <= _zz_when_ArraySlice_l158_331_3);
  assign when_ArraySlice_l159_331 = (_zz_when_ArraySlice_l159_331 <= _zz_when_ArraySlice_l159_331_2);
  assign _zz_realValue_0_331 = (_zz__zz_realValue_0_331 % _zz__zz_realValue_0_331_1);
  assign when_ArraySlice_l110_331 = (_zz_realValue_0_331 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_331) begin
      realValue_0_331 = (_zz_realValue_0_331_1 - _zz_realValue_0_331);
    end else begin
      realValue_0_331 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_331 = (_zz_when_ArraySlice_l166_331 <= _zz_when_ArraySlice_l166_331_2);
  assign when_ArraySlice_l158_332 = (_zz_when_ArraySlice_l158_332 <= _zz_when_ArraySlice_l158_332_3);
  assign when_ArraySlice_l159_332 = (_zz_when_ArraySlice_l159_332 <= _zz_when_ArraySlice_l159_332_2);
  assign _zz_realValue_0_332 = (_zz__zz_realValue_0_332 % _zz__zz_realValue_0_332_1);
  assign when_ArraySlice_l110_332 = (_zz_realValue_0_332 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_332) begin
      realValue_0_332 = (_zz_realValue_0_332_1 - _zz_realValue_0_332);
    end else begin
      realValue_0_332 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_332 = (_zz_when_ArraySlice_l166_332 <= _zz_when_ArraySlice_l166_332_2);
  assign when_ArraySlice_l158_333 = (_zz_when_ArraySlice_l158_333 <= _zz_when_ArraySlice_l158_333_3);
  assign when_ArraySlice_l159_333 = (_zz_when_ArraySlice_l159_333 <= _zz_when_ArraySlice_l159_333_2);
  assign _zz_realValue_0_333 = (_zz__zz_realValue_0_333 % _zz__zz_realValue_0_333_1);
  assign when_ArraySlice_l110_333 = (_zz_realValue_0_333 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_333) begin
      realValue_0_333 = (_zz_realValue_0_333_1 - _zz_realValue_0_333);
    end else begin
      realValue_0_333 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_333 = (_zz_when_ArraySlice_l166_333 <= _zz_when_ArraySlice_l166_333_2);
  assign when_ArraySlice_l158_334 = (_zz_when_ArraySlice_l158_334 <= _zz_when_ArraySlice_l158_334_3);
  assign when_ArraySlice_l159_334 = (_zz_when_ArraySlice_l159_334 <= _zz_when_ArraySlice_l159_334_2);
  assign _zz_realValue_0_334 = (_zz__zz_realValue_0_334 % _zz__zz_realValue_0_334_1);
  assign when_ArraySlice_l110_334 = (_zz_realValue_0_334 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_334) begin
      realValue_0_334 = (_zz_realValue_0_334_1 - _zz_realValue_0_334);
    end else begin
      realValue_0_334 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_334 = (_zz_when_ArraySlice_l166_334 <= _zz_when_ArraySlice_l166_334_2);
  assign when_ArraySlice_l158_335 = (_zz_when_ArraySlice_l158_335 <= _zz_when_ArraySlice_l158_335_3);
  assign when_ArraySlice_l159_335 = (_zz_when_ArraySlice_l159_335 <= _zz_when_ArraySlice_l159_335_2);
  assign _zz_realValue_0_335 = (_zz__zz_realValue_0_335 % _zz__zz_realValue_0_335_1);
  assign when_ArraySlice_l110_335 = (_zz_realValue_0_335 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_335) begin
      realValue_0_335 = (_zz_realValue_0_335_1 - _zz_realValue_0_335);
    end else begin
      realValue_0_335 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_335 = (_zz_when_ArraySlice_l166_335 <= _zz_when_ArraySlice_l166_335_2);
  assign when_ArraySlice_l257_5 = (! ((((((_zz_when_ArraySlice_l257_5_1 && _zz_when_ArraySlice_l257_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l257_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_5_4 && _zz_when_ArraySlice_l257_5_5) && (debug_4_41 == _zz_when_ArraySlice_l257_5_6)) && (debug_5_41 == 1'b1)) && (debug_6_41 == 1'b1)) && (debug_7_41 == 1'b1))));
  assign when_ArraySlice_l260_5 = (_zz_when_ArraySlice_l260_5_1 <= _zz_when_ArraySlice_l260_5_2);
  assign when_ArraySlice_l263_5 = (_zz_when_ArraySlice_l263_5 <= _zz_when_ArraySlice_l263_5_1);
  assign when_ArraySlice_l270_5 = (_zz_when_ArraySlice_l270_5 == 13'h0);
  assign when_ArraySlice_l274_5 = (_zz_when_ArraySlice_l274_5 == 7'h0);
  assign outputStreamArrayData_5_fire_9 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l275_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l275_5) && outputStreamArrayData_5_fire_9);
  assign _zz_realValue1_0_40 = (_zz__zz_realValue1_0_40 % _zz__zz_realValue1_0_40_1);
  assign when_ArraySlice_l95_40 = (_zz_realValue1_0_40 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_40) begin
      realValue1_0_40 = (_zz_realValue1_0_40_1 - _zz_realValue1_0_40);
    end else begin
      realValue1_0_40 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_5 = (_zz_when_ArraySlice_l277_5 < _zz_when_ArraySlice_l277_5_2);
  always @(*) begin
    debug_0_42 = 1'b0;
    if(when_ArraySlice_l158_336) begin
      if(when_ArraySlice_l159_336) begin
        debug_0_42 = 1'b1;
      end else begin
        debug_0_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_336) begin
        debug_0_42 = 1'b1;
      end else begin
        debug_0_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_42 = 1'b0;
    if(when_ArraySlice_l158_337) begin
      if(when_ArraySlice_l159_337) begin
        debug_1_42 = 1'b1;
      end else begin
        debug_1_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_337) begin
        debug_1_42 = 1'b1;
      end else begin
        debug_1_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_42 = 1'b0;
    if(when_ArraySlice_l158_338) begin
      if(when_ArraySlice_l159_338) begin
        debug_2_42 = 1'b1;
      end else begin
        debug_2_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_338) begin
        debug_2_42 = 1'b1;
      end else begin
        debug_2_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_42 = 1'b0;
    if(when_ArraySlice_l158_339) begin
      if(when_ArraySlice_l159_339) begin
        debug_3_42 = 1'b1;
      end else begin
        debug_3_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_339) begin
        debug_3_42 = 1'b1;
      end else begin
        debug_3_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_42 = 1'b0;
    if(when_ArraySlice_l158_340) begin
      if(when_ArraySlice_l159_340) begin
        debug_4_42 = 1'b1;
      end else begin
        debug_4_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_340) begin
        debug_4_42 = 1'b1;
      end else begin
        debug_4_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_42 = 1'b0;
    if(when_ArraySlice_l158_341) begin
      if(when_ArraySlice_l159_341) begin
        debug_5_42 = 1'b1;
      end else begin
        debug_5_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_341) begin
        debug_5_42 = 1'b1;
      end else begin
        debug_5_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_42 = 1'b0;
    if(when_ArraySlice_l158_342) begin
      if(when_ArraySlice_l159_342) begin
        debug_6_42 = 1'b1;
      end else begin
        debug_6_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_342) begin
        debug_6_42 = 1'b1;
      end else begin
        debug_6_42 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_42 = 1'b0;
    if(when_ArraySlice_l158_343) begin
      if(when_ArraySlice_l159_343) begin
        debug_7_42 = 1'b1;
      end else begin
        debug_7_42 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_343) begin
        debug_7_42 = 1'b1;
      end else begin
        debug_7_42 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_336 = (_zz_when_ArraySlice_l158_336 <= _zz_when_ArraySlice_l158_336_3);
  assign when_ArraySlice_l159_336 = (_zz_when_ArraySlice_l159_336 <= _zz_when_ArraySlice_l159_336_1);
  assign _zz_realValue_0_336 = (_zz__zz_realValue_0_336 % _zz__zz_realValue_0_336_1);
  assign when_ArraySlice_l110_336 = (_zz_realValue_0_336 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_336) begin
      realValue_0_336 = (_zz_realValue_0_336_1 - _zz_realValue_0_336);
    end else begin
      realValue_0_336 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_336 = (_zz_when_ArraySlice_l166_336 <= _zz_when_ArraySlice_l166_336_1);
  assign when_ArraySlice_l158_337 = (_zz_when_ArraySlice_l158_337 <= _zz_when_ArraySlice_l158_337_3);
  assign when_ArraySlice_l159_337 = (_zz_when_ArraySlice_l159_337 <= _zz_when_ArraySlice_l159_337_2);
  assign _zz_realValue_0_337 = (_zz__zz_realValue_0_337 % _zz__zz_realValue_0_337_1);
  assign when_ArraySlice_l110_337 = (_zz_realValue_0_337 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_337) begin
      realValue_0_337 = (_zz_realValue_0_337_1 - _zz_realValue_0_337);
    end else begin
      realValue_0_337 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_337 = (_zz_when_ArraySlice_l166_337 <= _zz_when_ArraySlice_l166_337_2);
  assign when_ArraySlice_l158_338 = (_zz_when_ArraySlice_l158_338 <= _zz_when_ArraySlice_l158_338_3);
  assign when_ArraySlice_l159_338 = (_zz_when_ArraySlice_l159_338 <= _zz_when_ArraySlice_l159_338_2);
  assign _zz_realValue_0_338 = (_zz__zz_realValue_0_338 % _zz__zz_realValue_0_338_1);
  assign when_ArraySlice_l110_338 = (_zz_realValue_0_338 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_338) begin
      realValue_0_338 = (_zz_realValue_0_338_1 - _zz_realValue_0_338);
    end else begin
      realValue_0_338 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_338 = (_zz_when_ArraySlice_l166_338 <= _zz_when_ArraySlice_l166_338_2);
  assign when_ArraySlice_l158_339 = (_zz_when_ArraySlice_l158_339 <= _zz_when_ArraySlice_l158_339_3);
  assign when_ArraySlice_l159_339 = (_zz_when_ArraySlice_l159_339 <= _zz_when_ArraySlice_l159_339_2);
  assign _zz_realValue_0_339 = (_zz__zz_realValue_0_339 % _zz__zz_realValue_0_339_1);
  assign when_ArraySlice_l110_339 = (_zz_realValue_0_339 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_339) begin
      realValue_0_339 = (_zz_realValue_0_339_1 - _zz_realValue_0_339);
    end else begin
      realValue_0_339 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_339 = (_zz_when_ArraySlice_l166_339 <= _zz_when_ArraySlice_l166_339_2);
  assign when_ArraySlice_l158_340 = (_zz_when_ArraySlice_l158_340 <= _zz_when_ArraySlice_l158_340_3);
  assign when_ArraySlice_l159_340 = (_zz_when_ArraySlice_l159_340 <= _zz_when_ArraySlice_l159_340_2);
  assign _zz_realValue_0_340 = (_zz__zz_realValue_0_340 % _zz__zz_realValue_0_340_1);
  assign when_ArraySlice_l110_340 = (_zz_realValue_0_340 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_340) begin
      realValue_0_340 = (_zz_realValue_0_340_1 - _zz_realValue_0_340);
    end else begin
      realValue_0_340 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_340 = (_zz_when_ArraySlice_l166_340 <= _zz_when_ArraySlice_l166_340_2);
  assign when_ArraySlice_l158_341 = (_zz_when_ArraySlice_l158_341 <= _zz_when_ArraySlice_l158_341_3);
  assign when_ArraySlice_l159_341 = (_zz_when_ArraySlice_l159_341 <= _zz_when_ArraySlice_l159_341_2);
  assign _zz_realValue_0_341 = (_zz__zz_realValue_0_341 % _zz__zz_realValue_0_341_1);
  assign when_ArraySlice_l110_341 = (_zz_realValue_0_341 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_341) begin
      realValue_0_341 = (_zz_realValue_0_341_1 - _zz_realValue_0_341);
    end else begin
      realValue_0_341 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_341 = (_zz_when_ArraySlice_l166_341 <= _zz_when_ArraySlice_l166_341_2);
  assign when_ArraySlice_l158_342 = (_zz_when_ArraySlice_l158_342 <= _zz_when_ArraySlice_l158_342_3);
  assign when_ArraySlice_l159_342 = (_zz_when_ArraySlice_l159_342 <= _zz_when_ArraySlice_l159_342_2);
  assign _zz_realValue_0_342 = (_zz__zz_realValue_0_342 % _zz__zz_realValue_0_342_1);
  assign when_ArraySlice_l110_342 = (_zz_realValue_0_342 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_342) begin
      realValue_0_342 = (_zz_realValue_0_342_1 - _zz_realValue_0_342);
    end else begin
      realValue_0_342 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_342 = (_zz_when_ArraySlice_l166_342 <= _zz_when_ArraySlice_l166_342_2);
  assign when_ArraySlice_l158_343 = (_zz_when_ArraySlice_l158_343 <= _zz_when_ArraySlice_l158_343_3);
  assign when_ArraySlice_l159_343 = (_zz_when_ArraySlice_l159_343 <= _zz_when_ArraySlice_l159_343_2);
  assign _zz_realValue_0_343 = (_zz__zz_realValue_0_343 % _zz__zz_realValue_0_343_1);
  assign when_ArraySlice_l110_343 = (_zz_realValue_0_343 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_343) begin
      realValue_0_343 = (_zz_realValue_0_343_1 - _zz_realValue_0_343);
    end else begin
      realValue_0_343 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_343 = (_zz_when_ArraySlice_l166_343 <= _zz_when_ArraySlice_l166_343_2);
  assign when_ArraySlice_l282_5 = (! ((((((_zz_when_ArraySlice_l282_5_1 && _zz_when_ArraySlice_l282_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l282_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_5_4 && _zz_when_ArraySlice_l282_5_5) && (debug_4_42 == _zz_when_ArraySlice_l282_5_6)) && (debug_5_42 == 1'b1)) && (debug_6_42 == 1'b1)) && (debug_7_42 == 1'b1))));
  assign when_ArraySlice_l285_5 = (_zz_when_ArraySlice_l285_5_1 <= _zz_when_ArraySlice_l285_5_2);
  assign when_ArraySlice_l288_5 = (_zz_when_ArraySlice_l288_5 <= _zz_when_ArraySlice_l288_5_1);
  assign outputStreamArrayData_5_fire_10 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l295_5 = ((_zz_when_ArraySlice_l295_5 == 13'h0) && outputStreamArrayData_5_fire_10);
  assign outputStreamArrayData_5_fire_11 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l306_5 = ((handshakeTimes_5_value == _zz_when_ArraySlice_l306_5) && outputStreamArrayData_5_fire_11);
  assign _zz_realValue1_0_41 = (_zz__zz_realValue1_0_41 % _zz__zz_realValue1_0_41_1);
  assign when_ArraySlice_l95_41 = (_zz_realValue1_0_41 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_41) begin
      realValue1_0_41 = (_zz_realValue1_0_41_1 - _zz_realValue1_0_41);
    end else begin
      realValue1_0_41 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_5 = (_zz_when_ArraySlice_l307_5 < _zz_when_ArraySlice_l307_5_2);
  always @(*) begin
    debug_0_43 = 1'b0;
    if(when_ArraySlice_l158_344) begin
      if(when_ArraySlice_l159_344) begin
        debug_0_43 = 1'b1;
      end else begin
        debug_0_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_344) begin
        debug_0_43 = 1'b1;
      end else begin
        debug_0_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_43 = 1'b0;
    if(when_ArraySlice_l158_345) begin
      if(when_ArraySlice_l159_345) begin
        debug_1_43 = 1'b1;
      end else begin
        debug_1_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_345) begin
        debug_1_43 = 1'b1;
      end else begin
        debug_1_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_43 = 1'b0;
    if(when_ArraySlice_l158_346) begin
      if(when_ArraySlice_l159_346) begin
        debug_2_43 = 1'b1;
      end else begin
        debug_2_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_346) begin
        debug_2_43 = 1'b1;
      end else begin
        debug_2_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_43 = 1'b0;
    if(when_ArraySlice_l158_347) begin
      if(when_ArraySlice_l159_347) begin
        debug_3_43 = 1'b1;
      end else begin
        debug_3_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_347) begin
        debug_3_43 = 1'b1;
      end else begin
        debug_3_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_43 = 1'b0;
    if(when_ArraySlice_l158_348) begin
      if(when_ArraySlice_l159_348) begin
        debug_4_43 = 1'b1;
      end else begin
        debug_4_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_348) begin
        debug_4_43 = 1'b1;
      end else begin
        debug_4_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_43 = 1'b0;
    if(when_ArraySlice_l158_349) begin
      if(when_ArraySlice_l159_349) begin
        debug_5_43 = 1'b1;
      end else begin
        debug_5_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_349) begin
        debug_5_43 = 1'b1;
      end else begin
        debug_5_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_43 = 1'b0;
    if(when_ArraySlice_l158_350) begin
      if(when_ArraySlice_l159_350) begin
        debug_6_43 = 1'b1;
      end else begin
        debug_6_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_350) begin
        debug_6_43 = 1'b1;
      end else begin
        debug_6_43 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_43 = 1'b0;
    if(when_ArraySlice_l158_351) begin
      if(when_ArraySlice_l159_351) begin
        debug_7_43 = 1'b1;
      end else begin
        debug_7_43 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_351) begin
        debug_7_43 = 1'b1;
      end else begin
        debug_7_43 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_344 = (_zz_when_ArraySlice_l158_344 <= _zz_when_ArraySlice_l158_344_3);
  assign when_ArraySlice_l159_344 = (_zz_when_ArraySlice_l159_344 <= _zz_when_ArraySlice_l159_344_1);
  assign _zz_realValue_0_344 = (_zz__zz_realValue_0_344 % _zz__zz_realValue_0_344_1);
  assign when_ArraySlice_l110_344 = (_zz_realValue_0_344 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_344) begin
      realValue_0_344 = (_zz_realValue_0_344_1 - _zz_realValue_0_344);
    end else begin
      realValue_0_344 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_344 = (_zz_when_ArraySlice_l166_344 <= _zz_when_ArraySlice_l166_344_1);
  assign when_ArraySlice_l158_345 = (_zz_when_ArraySlice_l158_345 <= _zz_when_ArraySlice_l158_345_3);
  assign when_ArraySlice_l159_345 = (_zz_when_ArraySlice_l159_345 <= _zz_when_ArraySlice_l159_345_2);
  assign _zz_realValue_0_345 = (_zz__zz_realValue_0_345 % _zz__zz_realValue_0_345_1);
  assign when_ArraySlice_l110_345 = (_zz_realValue_0_345 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_345) begin
      realValue_0_345 = (_zz_realValue_0_345_1 - _zz_realValue_0_345);
    end else begin
      realValue_0_345 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_345 = (_zz_when_ArraySlice_l166_345 <= _zz_when_ArraySlice_l166_345_2);
  assign when_ArraySlice_l158_346 = (_zz_when_ArraySlice_l158_346 <= _zz_when_ArraySlice_l158_346_3);
  assign when_ArraySlice_l159_346 = (_zz_when_ArraySlice_l159_346 <= _zz_when_ArraySlice_l159_346_2);
  assign _zz_realValue_0_346 = (_zz__zz_realValue_0_346 % _zz__zz_realValue_0_346_1);
  assign when_ArraySlice_l110_346 = (_zz_realValue_0_346 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_346) begin
      realValue_0_346 = (_zz_realValue_0_346_1 - _zz_realValue_0_346);
    end else begin
      realValue_0_346 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_346 = (_zz_when_ArraySlice_l166_346 <= _zz_when_ArraySlice_l166_346_2);
  assign when_ArraySlice_l158_347 = (_zz_when_ArraySlice_l158_347 <= _zz_when_ArraySlice_l158_347_3);
  assign when_ArraySlice_l159_347 = (_zz_when_ArraySlice_l159_347 <= _zz_when_ArraySlice_l159_347_2);
  assign _zz_realValue_0_347 = (_zz__zz_realValue_0_347 % _zz__zz_realValue_0_347_1);
  assign when_ArraySlice_l110_347 = (_zz_realValue_0_347 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_347) begin
      realValue_0_347 = (_zz_realValue_0_347_1 - _zz_realValue_0_347);
    end else begin
      realValue_0_347 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_347 = (_zz_when_ArraySlice_l166_347 <= _zz_when_ArraySlice_l166_347_2);
  assign when_ArraySlice_l158_348 = (_zz_when_ArraySlice_l158_348 <= _zz_when_ArraySlice_l158_348_3);
  assign when_ArraySlice_l159_348 = (_zz_when_ArraySlice_l159_348 <= _zz_when_ArraySlice_l159_348_2);
  assign _zz_realValue_0_348 = (_zz__zz_realValue_0_348 % _zz__zz_realValue_0_348_1);
  assign when_ArraySlice_l110_348 = (_zz_realValue_0_348 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_348) begin
      realValue_0_348 = (_zz_realValue_0_348_1 - _zz_realValue_0_348);
    end else begin
      realValue_0_348 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_348 = (_zz_when_ArraySlice_l166_348 <= _zz_when_ArraySlice_l166_348_2);
  assign when_ArraySlice_l158_349 = (_zz_when_ArraySlice_l158_349 <= _zz_when_ArraySlice_l158_349_3);
  assign when_ArraySlice_l159_349 = (_zz_when_ArraySlice_l159_349 <= _zz_when_ArraySlice_l159_349_2);
  assign _zz_realValue_0_349 = (_zz__zz_realValue_0_349 % _zz__zz_realValue_0_349_1);
  assign when_ArraySlice_l110_349 = (_zz_realValue_0_349 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_349) begin
      realValue_0_349 = (_zz_realValue_0_349_1 - _zz_realValue_0_349);
    end else begin
      realValue_0_349 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_349 = (_zz_when_ArraySlice_l166_349 <= _zz_when_ArraySlice_l166_349_2);
  assign when_ArraySlice_l158_350 = (_zz_when_ArraySlice_l158_350 <= _zz_when_ArraySlice_l158_350_3);
  assign when_ArraySlice_l159_350 = (_zz_when_ArraySlice_l159_350 <= _zz_when_ArraySlice_l159_350_2);
  assign _zz_realValue_0_350 = (_zz__zz_realValue_0_350 % _zz__zz_realValue_0_350_1);
  assign when_ArraySlice_l110_350 = (_zz_realValue_0_350 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_350) begin
      realValue_0_350 = (_zz_realValue_0_350_1 - _zz_realValue_0_350);
    end else begin
      realValue_0_350 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_350 = (_zz_when_ArraySlice_l166_350 <= _zz_when_ArraySlice_l166_350_2);
  assign when_ArraySlice_l158_351 = (_zz_when_ArraySlice_l158_351 <= _zz_when_ArraySlice_l158_351_3);
  assign when_ArraySlice_l159_351 = (_zz_when_ArraySlice_l159_351 <= _zz_when_ArraySlice_l159_351_2);
  assign _zz_realValue_0_351 = (_zz__zz_realValue_0_351 % _zz__zz_realValue_0_351_1);
  assign when_ArraySlice_l110_351 = (_zz_realValue_0_351 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_351) begin
      realValue_0_351 = (_zz_realValue_0_351_1 - _zz_realValue_0_351);
    end else begin
      realValue_0_351 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_351 = (_zz_when_ArraySlice_l166_351 <= _zz_when_ArraySlice_l166_351_2);
  assign when_ArraySlice_l314_5 = (! ((((((_zz_when_ArraySlice_l314_5_1 && _zz_when_ArraySlice_l314_5_2) && (holdReadOp_4 == _zz_when_ArraySlice_l314_5_3)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_5_4 && _zz_when_ArraySlice_l314_5_5) && (debug_4_43 == _zz_when_ArraySlice_l314_5_6)) && (debug_5_43 == 1'b1)) && (debug_6_43 == 1'b1)) && (debug_7_43 == 1'b1))));
  assign outputStreamArrayData_5_fire_12 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l318_5 = ((_zz_when_ArraySlice_l318_5 == 13'h0) && outputStreamArrayData_5_fire_12);
  assign when_ArraySlice_l304_5 = (allowPadding_5 && (_zz_when_ArraySlice_l304_5 <= _zz_when_ArraySlice_l304_5_1));
  assign outputStreamArrayData_5_fire_13 = (outputStreamArrayData_5_valid && outputStreamArrayData_5_ready);
  assign when_ArraySlice_l325_5 = (handshakeTimes_5_value == _zz_when_ArraySlice_l325_5);
  assign when_ArraySlice_l233_6 = (_zz_when_ArraySlice_l233_6 < _zz_when_ArraySlice_l233_6_3);
  assign when_ArraySlice_l234_6 = ((! holdReadOp_6) && (_zz_when_ArraySlice_l234_6 != 7'h0));
  assign _zz_outputStreamArrayData_6_valid_1 = (selectReadFifo_6 + _zz__zz_outputStreamArrayData_6_valid_1_1);
  assign _zz_17 = ({127'd0,1'b1} <<< _zz__zz_17);
  assign _zz_io_pop_ready_14 = outputStreamArrayData_6_ready;
  assign when_ArraySlice_l239_6 = (! holdReadOp_6);
  assign outputStreamArrayData_6_fire_7 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l240_6 = ((7'h01 < _zz_when_ArraySlice_l240_6) && outputStreamArrayData_6_fire_7);
  assign when_ArraySlice_l241_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l241_6);
  assign when_ArraySlice_l244_6 = (_zz_when_ArraySlice_l244_6 == 13'h0);
  assign outputStreamArrayData_6_fire_8 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l249_6 = ((_zz_when_ArraySlice_l249_6 == 7'h01) && outputStreamArrayData_6_fire_8);
  assign when_ArraySlice_l250_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l250_6);
  assign _zz_realValue1_0_42 = (_zz__zz_realValue1_0_42 % _zz__zz_realValue1_0_42_1);
  assign when_ArraySlice_l95_42 = (_zz_realValue1_0_42 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_42) begin
      realValue1_0_42 = (_zz_realValue1_0_42_1 - _zz_realValue1_0_42);
    end else begin
      realValue1_0_42 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_6 = (_zz_when_ArraySlice_l252_6 < _zz_when_ArraySlice_l252_6_2);
  always @(*) begin
    debug_0_44 = 1'b0;
    if(when_ArraySlice_l158_352) begin
      if(when_ArraySlice_l159_352) begin
        debug_0_44 = 1'b1;
      end else begin
        debug_0_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_352) begin
        debug_0_44 = 1'b1;
      end else begin
        debug_0_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_44 = 1'b0;
    if(when_ArraySlice_l158_353) begin
      if(when_ArraySlice_l159_353) begin
        debug_1_44 = 1'b1;
      end else begin
        debug_1_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_353) begin
        debug_1_44 = 1'b1;
      end else begin
        debug_1_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_44 = 1'b0;
    if(when_ArraySlice_l158_354) begin
      if(when_ArraySlice_l159_354) begin
        debug_2_44 = 1'b1;
      end else begin
        debug_2_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_354) begin
        debug_2_44 = 1'b1;
      end else begin
        debug_2_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_44 = 1'b0;
    if(when_ArraySlice_l158_355) begin
      if(when_ArraySlice_l159_355) begin
        debug_3_44 = 1'b1;
      end else begin
        debug_3_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_355) begin
        debug_3_44 = 1'b1;
      end else begin
        debug_3_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_44 = 1'b0;
    if(when_ArraySlice_l158_356) begin
      if(when_ArraySlice_l159_356) begin
        debug_4_44 = 1'b1;
      end else begin
        debug_4_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_356) begin
        debug_4_44 = 1'b1;
      end else begin
        debug_4_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_44 = 1'b0;
    if(when_ArraySlice_l158_357) begin
      if(when_ArraySlice_l159_357) begin
        debug_5_44 = 1'b1;
      end else begin
        debug_5_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_357) begin
        debug_5_44 = 1'b1;
      end else begin
        debug_5_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_44 = 1'b0;
    if(when_ArraySlice_l158_358) begin
      if(when_ArraySlice_l159_358) begin
        debug_6_44 = 1'b1;
      end else begin
        debug_6_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_358) begin
        debug_6_44 = 1'b1;
      end else begin
        debug_6_44 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_44 = 1'b0;
    if(when_ArraySlice_l158_359) begin
      if(when_ArraySlice_l159_359) begin
        debug_7_44 = 1'b1;
      end else begin
        debug_7_44 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_359) begin
        debug_7_44 = 1'b1;
      end else begin
        debug_7_44 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_352 = (_zz_when_ArraySlice_l158_352 <= _zz_when_ArraySlice_l158_352_3);
  assign when_ArraySlice_l159_352 = (_zz_when_ArraySlice_l159_352 <= _zz_when_ArraySlice_l159_352_1);
  assign _zz_realValue_0_352 = (_zz__zz_realValue_0_352 % _zz__zz_realValue_0_352_1);
  assign when_ArraySlice_l110_352 = (_zz_realValue_0_352 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_352) begin
      realValue_0_352 = (_zz_realValue_0_352_1 - _zz_realValue_0_352);
    end else begin
      realValue_0_352 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_352 = (_zz_when_ArraySlice_l166_352 <= _zz_when_ArraySlice_l166_352_1);
  assign when_ArraySlice_l158_353 = (_zz_when_ArraySlice_l158_353 <= _zz_when_ArraySlice_l158_353_3);
  assign when_ArraySlice_l159_353 = (_zz_when_ArraySlice_l159_353 <= _zz_when_ArraySlice_l159_353_2);
  assign _zz_realValue_0_353 = (_zz__zz_realValue_0_353 % _zz__zz_realValue_0_353_1);
  assign when_ArraySlice_l110_353 = (_zz_realValue_0_353 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_353) begin
      realValue_0_353 = (_zz_realValue_0_353_1 - _zz_realValue_0_353);
    end else begin
      realValue_0_353 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_353 = (_zz_when_ArraySlice_l166_353 <= _zz_when_ArraySlice_l166_353_2);
  assign when_ArraySlice_l158_354 = (_zz_when_ArraySlice_l158_354 <= _zz_when_ArraySlice_l158_354_3);
  assign when_ArraySlice_l159_354 = (_zz_when_ArraySlice_l159_354 <= _zz_when_ArraySlice_l159_354_2);
  assign _zz_realValue_0_354 = (_zz__zz_realValue_0_354 % _zz__zz_realValue_0_354_1);
  assign when_ArraySlice_l110_354 = (_zz_realValue_0_354 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_354) begin
      realValue_0_354 = (_zz_realValue_0_354_1 - _zz_realValue_0_354);
    end else begin
      realValue_0_354 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_354 = (_zz_when_ArraySlice_l166_354 <= _zz_when_ArraySlice_l166_354_2);
  assign when_ArraySlice_l158_355 = (_zz_when_ArraySlice_l158_355 <= _zz_when_ArraySlice_l158_355_3);
  assign when_ArraySlice_l159_355 = (_zz_when_ArraySlice_l159_355 <= _zz_when_ArraySlice_l159_355_2);
  assign _zz_realValue_0_355 = (_zz__zz_realValue_0_355 % _zz__zz_realValue_0_355_1);
  assign when_ArraySlice_l110_355 = (_zz_realValue_0_355 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_355) begin
      realValue_0_355 = (_zz_realValue_0_355_1 - _zz_realValue_0_355);
    end else begin
      realValue_0_355 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_355 = (_zz_when_ArraySlice_l166_355 <= _zz_when_ArraySlice_l166_355_2);
  assign when_ArraySlice_l158_356 = (_zz_when_ArraySlice_l158_356 <= _zz_when_ArraySlice_l158_356_3);
  assign when_ArraySlice_l159_356 = (_zz_when_ArraySlice_l159_356 <= _zz_when_ArraySlice_l159_356_2);
  assign _zz_realValue_0_356 = (_zz__zz_realValue_0_356 % _zz__zz_realValue_0_356_1);
  assign when_ArraySlice_l110_356 = (_zz_realValue_0_356 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_356) begin
      realValue_0_356 = (_zz_realValue_0_356_1 - _zz_realValue_0_356);
    end else begin
      realValue_0_356 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_356 = (_zz_when_ArraySlice_l166_356 <= _zz_when_ArraySlice_l166_356_2);
  assign when_ArraySlice_l158_357 = (_zz_when_ArraySlice_l158_357 <= _zz_when_ArraySlice_l158_357_3);
  assign when_ArraySlice_l159_357 = (_zz_when_ArraySlice_l159_357 <= _zz_when_ArraySlice_l159_357_2);
  assign _zz_realValue_0_357 = (_zz__zz_realValue_0_357 % _zz__zz_realValue_0_357_1);
  assign when_ArraySlice_l110_357 = (_zz_realValue_0_357 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_357) begin
      realValue_0_357 = (_zz_realValue_0_357_1 - _zz_realValue_0_357);
    end else begin
      realValue_0_357 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_357 = (_zz_when_ArraySlice_l166_357 <= _zz_when_ArraySlice_l166_357_2);
  assign when_ArraySlice_l158_358 = (_zz_when_ArraySlice_l158_358 <= _zz_when_ArraySlice_l158_358_3);
  assign when_ArraySlice_l159_358 = (_zz_when_ArraySlice_l159_358 <= _zz_when_ArraySlice_l159_358_2);
  assign _zz_realValue_0_358 = (_zz__zz_realValue_0_358 % _zz__zz_realValue_0_358_1);
  assign when_ArraySlice_l110_358 = (_zz_realValue_0_358 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_358) begin
      realValue_0_358 = (_zz_realValue_0_358_1 - _zz_realValue_0_358);
    end else begin
      realValue_0_358 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_358 = (_zz_when_ArraySlice_l166_358 <= _zz_when_ArraySlice_l166_358_2);
  assign when_ArraySlice_l158_359 = (_zz_when_ArraySlice_l158_359 <= _zz_when_ArraySlice_l158_359_3);
  assign when_ArraySlice_l159_359 = (_zz_when_ArraySlice_l159_359 <= _zz_when_ArraySlice_l159_359_2);
  assign _zz_realValue_0_359 = (_zz__zz_realValue_0_359 % _zz__zz_realValue_0_359_1);
  assign when_ArraySlice_l110_359 = (_zz_realValue_0_359 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_359) begin
      realValue_0_359 = (_zz_realValue_0_359_1 - _zz_realValue_0_359);
    end else begin
      realValue_0_359 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_359 = (_zz_when_ArraySlice_l166_359 <= _zz_when_ArraySlice_l166_359_2);
  assign when_ArraySlice_l257_6 = (! ((((((_zz_when_ArraySlice_l257_6 && _zz_when_ArraySlice_l257_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l257_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_6_3 && _zz_when_ArraySlice_l257_6_4) && (debug_4_44 == _zz_when_ArraySlice_l257_6_5)) && (debug_5_44 == 1'b1)) && (debug_6_44 == 1'b1)) && (debug_7_44 == 1'b1))));
  assign when_ArraySlice_l260_6 = (_zz_when_ArraySlice_l260_6_1 <= _zz_when_ArraySlice_l260_6_2);
  assign when_ArraySlice_l263_6 = (_zz_when_ArraySlice_l263_6 <= _zz_when_ArraySlice_l263_6_1);
  assign when_ArraySlice_l270_6 = (_zz_when_ArraySlice_l270_6 == 13'h0);
  assign when_ArraySlice_l274_6 = (_zz_when_ArraySlice_l274_6 == 7'h0);
  assign outputStreamArrayData_6_fire_9 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l275_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l275_6) && outputStreamArrayData_6_fire_9);
  assign _zz_realValue1_0_43 = (_zz__zz_realValue1_0_43 % _zz__zz_realValue1_0_43_1);
  assign when_ArraySlice_l95_43 = (_zz_realValue1_0_43 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_43) begin
      realValue1_0_43 = (_zz_realValue1_0_43_1 - _zz_realValue1_0_43);
    end else begin
      realValue1_0_43 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_6 = (_zz_when_ArraySlice_l277_6 < _zz_when_ArraySlice_l277_6_2);
  always @(*) begin
    debug_0_45 = 1'b0;
    if(when_ArraySlice_l158_360) begin
      if(when_ArraySlice_l159_360) begin
        debug_0_45 = 1'b1;
      end else begin
        debug_0_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_360) begin
        debug_0_45 = 1'b1;
      end else begin
        debug_0_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_45 = 1'b0;
    if(when_ArraySlice_l158_361) begin
      if(when_ArraySlice_l159_361) begin
        debug_1_45 = 1'b1;
      end else begin
        debug_1_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_361) begin
        debug_1_45 = 1'b1;
      end else begin
        debug_1_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_45 = 1'b0;
    if(when_ArraySlice_l158_362) begin
      if(when_ArraySlice_l159_362) begin
        debug_2_45 = 1'b1;
      end else begin
        debug_2_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_362) begin
        debug_2_45 = 1'b1;
      end else begin
        debug_2_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_45 = 1'b0;
    if(when_ArraySlice_l158_363) begin
      if(when_ArraySlice_l159_363) begin
        debug_3_45 = 1'b1;
      end else begin
        debug_3_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_363) begin
        debug_3_45 = 1'b1;
      end else begin
        debug_3_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_45 = 1'b0;
    if(when_ArraySlice_l158_364) begin
      if(when_ArraySlice_l159_364) begin
        debug_4_45 = 1'b1;
      end else begin
        debug_4_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_364) begin
        debug_4_45 = 1'b1;
      end else begin
        debug_4_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_45 = 1'b0;
    if(when_ArraySlice_l158_365) begin
      if(when_ArraySlice_l159_365) begin
        debug_5_45 = 1'b1;
      end else begin
        debug_5_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_365) begin
        debug_5_45 = 1'b1;
      end else begin
        debug_5_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_45 = 1'b0;
    if(when_ArraySlice_l158_366) begin
      if(when_ArraySlice_l159_366) begin
        debug_6_45 = 1'b1;
      end else begin
        debug_6_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_366) begin
        debug_6_45 = 1'b1;
      end else begin
        debug_6_45 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_45 = 1'b0;
    if(when_ArraySlice_l158_367) begin
      if(when_ArraySlice_l159_367) begin
        debug_7_45 = 1'b1;
      end else begin
        debug_7_45 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_367) begin
        debug_7_45 = 1'b1;
      end else begin
        debug_7_45 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_360 = (_zz_when_ArraySlice_l158_360 <= _zz_when_ArraySlice_l158_360_3);
  assign when_ArraySlice_l159_360 = (_zz_when_ArraySlice_l159_360 <= _zz_when_ArraySlice_l159_360_1);
  assign _zz_realValue_0_360 = (_zz__zz_realValue_0_360 % _zz__zz_realValue_0_360_1);
  assign when_ArraySlice_l110_360 = (_zz_realValue_0_360 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_360) begin
      realValue_0_360 = (_zz_realValue_0_360_1 - _zz_realValue_0_360);
    end else begin
      realValue_0_360 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_360 = (_zz_when_ArraySlice_l166_360 <= _zz_when_ArraySlice_l166_360_1);
  assign when_ArraySlice_l158_361 = (_zz_when_ArraySlice_l158_361 <= _zz_when_ArraySlice_l158_361_3);
  assign when_ArraySlice_l159_361 = (_zz_when_ArraySlice_l159_361 <= _zz_when_ArraySlice_l159_361_2);
  assign _zz_realValue_0_361 = (_zz__zz_realValue_0_361 % _zz__zz_realValue_0_361_1);
  assign when_ArraySlice_l110_361 = (_zz_realValue_0_361 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_361) begin
      realValue_0_361 = (_zz_realValue_0_361_1 - _zz_realValue_0_361);
    end else begin
      realValue_0_361 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_361 = (_zz_when_ArraySlice_l166_361 <= _zz_when_ArraySlice_l166_361_2);
  assign when_ArraySlice_l158_362 = (_zz_when_ArraySlice_l158_362 <= _zz_when_ArraySlice_l158_362_3);
  assign when_ArraySlice_l159_362 = (_zz_when_ArraySlice_l159_362 <= _zz_when_ArraySlice_l159_362_2);
  assign _zz_realValue_0_362 = (_zz__zz_realValue_0_362 % _zz__zz_realValue_0_362_1);
  assign when_ArraySlice_l110_362 = (_zz_realValue_0_362 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_362) begin
      realValue_0_362 = (_zz_realValue_0_362_1 - _zz_realValue_0_362);
    end else begin
      realValue_0_362 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_362 = (_zz_when_ArraySlice_l166_362 <= _zz_when_ArraySlice_l166_362_2);
  assign when_ArraySlice_l158_363 = (_zz_when_ArraySlice_l158_363 <= _zz_when_ArraySlice_l158_363_3);
  assign when_ArraySlice_l159_363 = (_zz_when_ArraySlice_l159_363 <= _zz_when_ArraySlice_l159_363_2);
  assign _zz_realValue_0_363 = (_zz__zz_realValue_0_363 % _zz__zz_realValue_0_363_1);
  assign when_ArraySlice_l110_363 = (_zz_realValue_0_363 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_363) begin
      realValue_0_363 = (_zz_realValue_0_363_1 - _zz_realValue_0_363);
    end else begin
      realValue_0_363 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_363 = (_zz_when_ArraySlice_l166_363 <= _zz_when_ArraySlice_l166_363_2);
  assign when_ArraySlice_l158_364 = (_zz_when_ArraySlice_l158_364 <= _zz_when_ArraySlice_l158_364_3);
  assign when_ArraySlice_l159_364 = (_zz_when_ArraySlice_l159_364 <= _zz_when_ArraySlice_l159_364_2);
  assign _zz_realValue_0_364 = (_zz__zz_realValue_0_364 % _zz__zz_realValue_0_364_1);
  assign when_ArraySlice_l110_364 = (_zz_realValue_0_364 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_364) begin
      realValue_0_364 = (_zz_realValue_0_364_1 - _zz_realValue_0_364);
    end else begin
      realValue_0_364 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_364 = (_zz_when_ArraySlice_l166_364 <= _zz_when_ArraySlice_l166_364_2);
  assign when_ArraySlice_l158_365 = (_zz_when_ArraySlice_l158_365 <= _zz_when_ArraySlice_l158_365_3);
  assign when_ArraySlice_l159_365 = (_zz_when_ArraySlice_l159_365 <= _zz_when_ArraySlice_l159_365_2);
  assign _zz_realValue_0_365 = (_zz__zz_realValue_0_365 % _zz__zz_realValue_0_365_1);
  assign when_ArraySlice_l110_365 = (_zz_realValue_0_365 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_365) begin
      realValue_0_365 = (_zz_realValue_0_365_1 - _zz_realValue_0_365);
    end else begin
      realValue_0_365 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_365 = (_zz_when_ArraySlice_l166_365 <= _zz_when_ArraySlice_l166_365_2);
  assign when_ArraySlice_l158_366 = (_zz_when_ArraySlice_l158_366 <= _zz_when_ArraySlice_l158_366_3);
  assign when_ArraySlice_l159_366 = (_zz_when_ArraySlice_l159_366 <= _zz_when_ArraySlice_l159_366_2);
  assign _zz_realValue_0_366 = (_zz__zz_realValue_0_366 % _zz__zz_realValue_0_366_1);
  assign when_ArraySlice_l110_366 = (_zz_realValue_0_366 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_366) begin
      realValue_0_366 = (_zz_realValue_0_366_1 - _zz_realValue_0_366);
    end else begin
      realValue_0_366 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_366 = (_zz_when_ArraySlice_l166_366 <= _zz_when_ArraySlice_l166_366_2);
  assign when_ArraySlice_l158_367 = (_zz_when_ArraySlice_l158_367 <= _zz_when_ArraySlice_l158_367_3);
  assign when_ArraySlice_l159_367 = (_zz_when_ArraySlice_l159_367 <= _zz_when_ArraySlice_l159_367_2);
  assign _zz_realValue_0_367 = (_zz__zz_realValue_0_367 % _zz__zz_realValue_0_367_1);
  assign when_ArraySlice_l110_367 = (_zz_realValue_0_367 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_367) begin
      realValue_0_367 = (_zz_realValue_0_367_1 - _zz_realValue_0_367);
    end else begin
      realValue_0_367 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_367 = (_zz_when_ArraySlice_l166_367 <= _zz_when_ArraySlice_l166_367_2);
  assign when_ArraySlice_l282_6 = (! ((((((_zz_when_ArraySlice_l282_6 && _zz_when_ArraySlice_l282_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l282_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_6_3 && _zz_when_ArraySlice_l282_6_4) && (debug_4_45 == _zz_when_ArraySlice_l282_6_5)) && (debug_5_45 == 1'b1)) && (debug_6_45 == 1'b1)) && (debug_7_45 == 1'b1))));
  assign when_ArraySlice_l285_6 = (_zz_when_ArraySlice_l285_6_1 <= _zz_when_ArraySlice_l285_6_2);
  assign when_ArraySlice_l288_6 = (_zz_when_ArraySlice_l288_6 <= _zz_when_ArraySlice_l288_6_1);
  assign outputStreamArrayData_6_fire_10 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l295_6 = ((_zz_when_ArraySlice_l295_6 == 13'h0) && outputStreamArrayData_6_fire_10);
  assign outputStreamArrayData_6_fire_11 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l306_6 = ((handshakeTimes_6_value == _zz_when_ArraySlice_l306_6) && outputStreamArrayData_6_fire_11);
  assign _zz_realValue1_0_44 = (_zz__zz_realValue1_0_44 % _zz__zz_realValue1_0_44_1);
  assign when_ArraySlice_l95_44 = (_zz_realValue1_0_44 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_44) begin
      realValue1_0_44 = (_zz_realValue1_0_44_1 - _zz_realValue1_0_44);
    end else begin
      realValue1_0_44 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_6 = (_zz_when_ArraySlice_l307_6 < _zz_when_ArraySlice_l307_6_2);
  always @(*) begin
    debug_0_46 = 1'b0;
    if(when_ArraySlice_l158_368) begin
      if(when_ArraySlice_l159_368) begin
        debug_0_46 = 1'b1;
      end else begin
        debug_0_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_368) begin
        debug_0_46 = 1'b1;
      end else begin
        debug_0_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_46 = 1'b0;
    if(when_ArraySlice_l158_369) begin
      if(when_ArraySlice_l159_369) begin
        debug_1_46 = 1'b1;
      end else begin
        debug_1_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_369) begin
        debug_1_46 = 1'b1;
      end else begin
        debug_1_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_46 = 1'b0;
    if(when_ArraySlice_l158_370) begin
      if(when_ArraySlice_l159_370) begin
        debug_2_46 = 1'b1;
      end else begin
        debug_2_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_370) begin
        debug_2_46 = 1'b1;
      end else begin
        debug_2_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_46 = 1'b0;
    if(when_ArraySlice_l158_371) begin
      if(when_ArraySlice_l159_371) begin
        debug_3_46 = 1'b1;
      end else begin
        debug_3_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_371) begin
        debug_3_46 = 1'b1;
      end else begin
        debug_3_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_46 = 1'b0;
    if(when_ArraySlice_l158_372) begin
      if(when_ArraySlice_l159_372) begin
        debug_4_46 = 1'b1;
      end else begin
        debug_4_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_372) begin
        debug_4_46 = 1'b1;
      end else begin
        debug_4_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_46 = 1'b0;
    if(when_ArraySlice_l158_373) begin
      if(when_ArraySlice_l159_373) begin
        debug_5_46 = 1'b1;
      end else begin
        debug_5_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_373) begin
        debug_5_46 = 1'b1;
      end else begin
        debug_5_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_46 = 1'b0;
    if(when_ArraySlice_l158_374) begin
      if(when_ArraySlice_l159_374) begin
        debug_6_46 = 1'b1;
      end else begin
        debug_6_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_374) begin
        debug_6_46 = 1'b1;
      end else begin
        debug_6_46 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_46 = 1'b0;
    if(when_ArraySlice_l158_375) begin
      if(when_ArraySlice_l159_375) begin
        debug_7_46 = 1'b1;
      end else begin
        debug_7_46 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_375) begin
        debug_7_46 = 1'b1;
      end else begin
        debug_7_46 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_368 = (_zz_when_ArraySlice_l158_368 <= _zz_when_ArraySlice_l158_368_3);
  assign when_ArraySlice_l159_368 = (_zz_when_ArraySlice_l159_368 <= _zz_when_ArraySlice_l159_368_1);
  assign _zz_realValue_0_368 = (_zz__zz_realValue_0_368 % _zz__zz_realValue_0_368_1);
  assign when_ArraySlice_l110_368 = (_zz_realValue_0_368 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_368) begin
      realValue_0_368 = (_zz_realValue_0_368_1 - _zz_realValue_0_368);
    end else begin
      realValue_0_368 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_368 = (_zz_when_ArraySlice_l166_368 <= _zz_when_ArraySlice_l166_368_1);
  assign when_ArraySlice_l158_369 = (_zz_when_ArraySlice_l158_369 <= _zz_when_ArraySlice_l158_369_3);
  assign when_ArraySlice_l159_369 = (_zz_when_ArraySlice_l159_369 <= _zz_when_ArraySlice_l159_369_2);
  assign _zz_realValue_0_369 = (_zz__zz_realValue_0_369 % _zz__zz_realValue_0_369_1);
  assign when_ArraySlice_l110_369 = (_zz_realValue_0_369 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_369) begin
      realValue_0_369 = (_zz_realValue_0_369_1 - _zz_realValue_0_369);
    end else begin
      realValue_0_369 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_369 = (_zz_when_ArraySlice_l166_369 <= _zz_when_ArraySlice_l166_369_2);
  assign when_ArraySlice_l158_370 = (_zz_when_ArraySlice_l158_370 <= _zz_when_ArraySlice_l158_370_3);
  assign when_ArraySlice_l159_370 = (_zz_when_ArraySlice_l159_370 <= _zz_when_ArraySlice_l159_370_2);
  assign _zz_realValue_0_370 = (_zz__zz_realValue_0_370 % _zz__zz_realValue_0_370_1);
  assign when_ArraySlice_l110_370 = (_zz_realValue_0_370 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_370) begin
      realValue_0_370 = (_zz_realValue_0_370_1 - _zz_realValue_0_370);
    end else begin
      realValue_0_370 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_370 = (_zz_when_ArraySlice_l166_370 <= _zz_when_ArraySlice_l166_370_2);
  assign when_ArraySlice_l158_371 = (_zz_when_ArraySlice_l158_371 <= _zz_when_ArraySlice_l158_371_3);
  assign when_ArraySlice_l159_371 = (_zz_when_ArraySlice_l159_371 <= _zz_when_ArraySlice_l159_371_2);
  assign _zz_realValue_0_371 = (_zz__zz_realValue_0_371 % _zz__zz_realValue_0_371_1);
  assign when_ArraySlice_l110_371 = (_zz_realValue_0_371 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_371) begin
      realValue_0_371 = (_zz_realValue_0_371_1 - _zz_realValue_0_371);
    end else begin
      realValue_0_371 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_371 = (_zz_when_ArraySlice_l166_371 <= _zz_when_ArraySlice_l166_371_2);
  assign when_ArraySlice_l158_372 = (_zz_when_ArraySlice_l158_372 <= _zz_when_ArraySlice_l158_372_3);
  assign when_ArraySlice_l159_372 = (_zz_when_ArraySlice_l159_372 <= _zz_when_ArraySlice_l159_372_2);
  assign _zz_realValue_0_372 = (_zz__zz_realValue_0_372 % _zz__zz_realValue_0_372_1);
  assign when_ArraySlice_l110_372 = (_zz_realValue_0_372 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_372) begin
      realValue_0_372 = (_zz_realValue_0_372_1 - _zz_realValue_0_372);
    end else begin
      realValue_0_372 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_372 = (_zz_when_ArraySlice_l166_372 <= _zz_when_ArraySlice_l166_372_2);
  assign when_ArraySlice_l158_373 = (_zz_when_ArraySlice_l158_373 <= _zz_when_ArraySlice_l158_373_3);
  assign when_ArraySlice_l159_373 = (_zz_when_ArraySlice_l159_373 <= _zz_when_ArraySlice_l159_373_2);
  assign _zz_realValue_0_373 = (_zz__zz_realValue_0_373 % _zz__zz_realValue_0_373_1);
  assign when_ArraySlice_l110_373 = (_zz_realValue_0_373 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_373) begin
      realValue_0_373 = (_zz_realValue_0_373_1 - _zz_realValue_0_373);
    end else begin
      realValue_0_373 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_373 = (_zz_when_ArraySlice_l166_373 <= _zz_when_ArraySlice_l166_373_2);
  assign when_ArraySlice_l158_374 = (_zz_when_ArraySlice_l158_374 <= _zz_when_ArraySlice_l158_374_3);
  assign when_ArraySlice_l159_374 = (_zz_when_ArraySlice_l159_374 <= _zz_when_ArraySlice_l159_374_2);
  assign _zz_realValue_0_374 = (_zz__zz_realValue_0_374 % _zz__zz_realValue_0_374_1);
  assign when_ArraySlice_l110_374 = (_zz_realValue_0_374 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_374) begin
      realValue_0_374 = (_zz_realValue_0_374_1 - _zz_realValue_0_374);
    end else begin
      realValue_0_374 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_374 = (_zz_when_ArraySlice_l166_374 <= _zz_when_ArraySlice_l166_374_2);
  assign when_ArraySlice_l158_375 = (_zz_when_ArraySlice_l158_375 <= _zz_when_ArraySlice_l158_375_3);
  assign when_ArraySlice_l159_375 = (_zz_when_ArraySlice_l159_375 <= _zz_when_ArraySlice_l159_375_2);
  assign _zz_realValue_0_375 = (_zz__zz_realValue_0_375 % _zz__zz_realValue_0_375_1);
  assign when_ArraySlice_l110_375 = (_zz_realValue_0_375 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_375) begin
      realValue_0_375 = (_zz_realValue_0_375_1 - _zz_realValue_0_375);
    end else begin
      realValue_0_375 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_375 = (_zz_when_ArraySlice_l166_375 <= _zz_when_ArraySlice_l166_375_2);
  assign when_ArraySlice_l314_6 = (! ((((((_zz_when_ArraySlice_l314_6 && _zz_when_ArraySlice_l314_6_1) && (holdReadOp_4 == _zz_when_ArraySlice_l314_6_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_6_3 && _zz_when_ArraySlice_l314_6_4) && (debug_4_46 == _zz_when_ArraySlice_l314_6_5)) && (debug_5_46 == 1'b1)) && (debug_6_46 == 1'b1)) && (debug_7_46 == 1'b1))));
  assign outputStreamArrayData_6_fire_12 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l318_6 = ((_zz_when_ArraySlice_l318_6 == 13'h0) && outputStreamArrayData_6_fire_12);
  assign when_ArraySlice_l304_6 = (allowPadding_6 && (_zz_when_ArraySlice_l304_6 <= _zz_when_ArraySlice_l304_6_1));
  assign outputStreamArrayData_6_fire_13 = (outputStreamArrayData_6_valid && outputStreamArrayData_6_ready);
  assign when_ArraySlice_l325_6 = (handshakeTimes_6_value == _zz_when_ArraySlice_l325_6);
  assign when_ArraySlice_l233_7 = (_zz_when_ArraySlice_l233_7 < _zz_when_ArraySlice_l233_7_3);
  assign when_ArraySlice_l234_7 = ((! holdReadOp_7) && (_zz_when_ArraySlice_l234_7 != 7'h0));
  assign _zz_outputStreamArrayData_7_valid_1 = (selectReadFifo_7 + _zz__zz_outputStreamArrayData_7_valid_1_1);
  assign _zz_18 = ({127'd0,1'b1} <<< _zz__zz_18);
  assign _zz_io_pop_ready_15 = outputStreamArrayData_7_ready;
  assign when_ArraySlice_l239_7 = (! holdReadOp_7);
  assign outputStreamArrayData_7_fire_7 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l240_7 = ((7'h01 < _zz_when_ArraySlice_l240_7) && outputStreamArrayData_7_fire_7);
  assign when_ArraySlice_l241_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l241_7);
  assign when_ArraySlice_l244_7 = (_zz_when_ArraySlice_l244_7 == 13'h0);
  assign outputStreamArrayData_7_fire_8 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l249_7 = ((_zz_when_ArraySlice_l249_7 == 7'h01) && outputStreamArrayData_7_fire_8);
  assign when_ArraySlice_l250_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l250_7);
  assign _zz_realValue1_0_45 = (_zz__zz_realValue1_0_45 % _zz__zz_realValue1_0_45_1);
  assign when_ArraySlice_l95_45 = (_zz_realValue1_0_45 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_45) begin
      realValue1_0_45 = (_zz_realValue1_0_45_1 - _zz_realValue1_0_45);
    end else begin
      realValue1_0_45 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l252_7 = (_zz_when_ArraySlice_l252_7 < _zz_when_ArraySlice_l252_7_2);
  always @(*) begin
    debug_0_47 = 1'b0;
    if(when_ArraySlice_l158_376) begin
      if(when_ArraySlice_l159_376) begin
        debug_0_47 = 1'b1;
      end else begin
        debug_0_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_376) begin
        debug_0_47 = 1'b1;
      end else begin
        debug_0_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_47 = 1'b0;
    if(when_ArraySlice_l158_377) begin
      if(when_ArraySlice_l159_377) begin
        debug_1_47 = 1'b1;
      end else begin
        debug_1_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_377) begin
        debug_1_47 = 1'b1;
      end else begin
        debug_1_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_47 = 1'b0;
    if(when_ArraySlice_l158_378) begin
      if(when_ArraySlice_l159_378) begin
        debug_2_47 = 1'b1;
      end else begin
        debug_2_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_378) begin
        debug_2_47 = 1'b1;
      end else begin
        debug_2_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_47 = 1'b0;
    if(when_ArraySlice_l158_379) begin
      if(when_ArraySlice_l159_379) begin
        debug_3_47 = 1'b1;
      end else begin
        debug_3_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_379) begin
        debug_3_47 = 1'b1;
      end else begin
        debug_3_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_47 = 1'b0;
    if(when_ArraySlice_l158_380) begin
      if(when_ArraySlice_l159_380) begin
        debug_4_47 = 1'b1;
      end else begin
        debug_4_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_380) begin
        debug_4_47 = 1'b1;
      end else begin
        debug_4_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_47 = 1'b0;
    if(when_ArraySlice_l158_381) begin
      if(when_ArraySlice_l159_381) begin
        debug_5_47 = 1'b1;
      end else begin
        debug_5_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_381) begin
        debug_5_47 = 1'b1;
      end else begin
        debug_5_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_47 = 1'b0;
    if(when_ArraySlice_l158_382) begin
      if(when_ArraySlice_l159_382) begin
        debug_6_47 = 1'b1;
      end else begin
        debug_6_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_382) begin
        debug_6_47 = 1'b1;
      end else begin
        debug_6_47 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_47 = 1'b0;
    if(when_ArraySlice_l158_383) begin
      if(when_ArraySlice_l159_383) begin
        debug_7_47 = 1'b1;
      end else begin
        debug_7_47 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_383) begin
        debug_7_47 = 1'b1;
      end else begin
        debug_7_47 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_376 = (_zz_when_ArraySlice_l158_376 <= _zz_when_ArraySlice_l158_376_3);
  assign when_ArraySlice_l159_376 = (_zz_when_ArraySlice_l159_376 <= _zz_when_ArraySlice_l159_376_1);
  assign _zz_realValue_0_376 = (_zz__zz_realValue_0_376 % _zz__zz_realValue_0_376_1);
  assign when_ArraySlice_l110_376 = (_zz_realValue_0_376 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_376) begin
      realValue_0_376 = (_zz_realValue_0_376_1 - _zz_realValue_0_376);
    end else begin
      realValue_0_376 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_376 = (_zz_when_ArraySlice_l166_376 <= _zz_when_ArraySlice_l166_376_1);
  assign when_ArraySlice_l158_377 = (_zz_when_ArraySlice_l158_377 <= _zz_when_ArraySlice_l158_377_3);
  assign when_ArraySlice_l159_377 = (_zz_when_ArraySlice_l159_377 <= _zz_when_ArraySlice_l159_377_2);
  assign _zz_realValue_0_377 = (_zz__zz_realValue_0_377 % _zz__zz_realValue_0_377_1);
  assign when_ArraySlice_l110_377 = (_zz_realValue_0_377 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_377) begin
      realValue_0_377 = (_zz_realValue_0_377_1 - _zz_realValue_0_377);
    end else begin
      realValue_0_377 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_377 = (_zz_when_ArraySlice_l166_377 <= _zz_when_ArraySlice_l166_377_2);
  assign when_ArraySlice_l158_378 = (_zz_when_ArraySlice_l158_378 <= _zz_when_ArraySlice_l158_378_3);
  assign when_ArraySlice_l159_378 = (_zz_when_ArraySlice_l159_378 <= _zz_when_ArraySlice_l159_378_2);
  assign _zz_realValue_0_378 = (_zz__zz_realValue_0_378 % _zz__zz_realValue_0_378_1);
  assign when_ArraySlice_l110_378 = (_zz_realValue_0_378 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_378) begin
      realValue_0_378 = (_zz_realValue_0_378_1 - _zz_realValue_0_378);
    end else begin
      realValue_0_378 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_378 = (_zz_when_ArraySlice_l166_378 <= _zz_when_ArraySlice_l166_378_2);
  assign when_ArraySlice_l158_379 = (_zz_when_ArraySlice_l158_379 <= _zz_when_ArraySlice_l158_379_3);
  assign when_ArraySlice_l159_379 = (_zz_when_ArraySlice_l159_379 <= _zz_when_ArraySlice_l159_379_2);
  assign _zz_realValue_0_379 = (_zz__zz_realValue_0_379 % _zz__zz_realValue_0_379_1);
  assign when_ArraySlice_l110_379 = (_zz_realValue_0_379 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_379) begin
      realValue_0_379 = (_zz_realValue_0_379_1 - _zz_realValue_0_379);
    end else begin
      realValue_0_379 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_379 = (_zz_when_ArraySlice_l166_379 <= _zz_when_ArraySlice_l166_379_2);
  assign when_ArraySlice_l158_380 = (_zz_when_ArraySlice_l158_380 <= _zz_when_ArraySlice_l158_380_3);
  assign when_ArraySlice_l159_380 = (_zz_when_ArraySlice_l159_380 <= _zz_when_ArraySlice_l159_380_2);
  assign _zz_realValue_0_380 = (_zz__zz_realValue_0_380 % _zz__zz_realValue_0_380_1);
  assign when_ArraySlice_l110_380 = (_zz_realValue_0_380 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_380) begin
      realValue_0_380 = (_zz_realValue_0_380_1 - _zz_realValue_0_380);
    end else begin
      realValue_0_380 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_380 = (_zz_when_ArraySlice_l166_380 <= _zz_when_ArraySlice_l166_380_2);
  assign when_ArraySlice_l158_381 = (_zz_when_ArraySlice_l158_381 <= _zz_when_ArraySlice_l158_381_3);
  assign when_ArraySlice_l159_381 = (_zz_when_ArraySlice_l159_381 <= _zz_when_ArraySlice_l159_381_2);
  assign _zz_realValue_0_381 = (_zz__zz_realValue_0_381 % _zz__zz_realValue_0_381_1);
  assign when_ArraySlice_l110_381 = (_zz_realValue_0_381 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_381) begin
      realValue_0_381 = (_zz_realValue_0_381_1 - _zz_realValue_0_381);
    end else begin
      realValue_0_381 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_381 = (_zz_when_ArraySlice_l166_381 <= _zz_when_ArraySlice_l166_381_2);
  assign when_ArraySlice_l158_382 = (_zz_when_ArraySlice_l158_382 <= _zz_when_ArraySlice_l158_382_3);
  assign when_ArraySlice_l159_382 = (_zz_when_ArraySlice_l159_382 <= _zz_when_ArraySlice_l159_382_2);
  assign _zz_realValue_0_382 = (_zz__zz_realValue_0_382 % _zz__zz_realValue_0_382_1);
  assign when_ArraySlice_l110_382 = (_zz_realValue_0_382 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_382) begin
      realValue_0_382 = (_zz_realValue_0_382_1 - _zz_realValue_0_382);
    end else begin
      realValue_0_382 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_382 = (_zz_when_ArraySlice_l166_382 <= _zz_when_ArraySlice_l166_382_2);
  assign when_ArraySlice_l158_383 = (_zz_when_ArraySlice_l158_383 <= _zz_when_ArraySlice_l158_383_3);
  assign when_ArraySlice_l159_383 = (_zz_when_ArraySlice_l159_383 <= _zz_when_ArraySlice_l159_383_2);
  assign _zz_realValue_0_383 = (_zz__zz_realValue_0_383 % _zz__zz_realValue_0_383_1);
  assign when_ArraySlice_l110_383 = (_zz_realValue_0_383 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_383) begin
      realValue_0_383 = (_zz_realValue_0_383_1 - _zz_realValue_0_383);
    end else begin
      realValue_0_383 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_383 = (_zz_when_ArraySlice_l166_383 <= _zz_when_ArraySlice_l166_383_2);
  assign when_ArraySlice_l257_7 = (! ((((((_zz_when_ArraySlice_l257_7 && _zz_when_ArraySlice_l257_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l257_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l257_7_3 && _zz_when_ArraySlice_l257_7_4) && (debug_4_47 == _zz_when_ArraySlice_l257_7_5)) && (debug_5_47 == 1'b1)) && (debug_6_47 == 1'b1)) && (debug_7_47 == 1'b1))));
  assign when_ArraySlice_l260_7 = (_zz_when_ArraySlice_l260_7_1 <= _zz_when_ArraySlice_l260_7_2);
  assign when_ArraySlice_l263_7 = (_zz_when_ArraySlice_l263_7 <= _zz_when_ArraySlice_l263_7_1);
  assign when_ArraySlice_l270_7 = (_zz_when_ArraySlice_l270_7 == 13'h0);
  assign when_ArraySlice_l274_7 = (_zz_when_ArraySlice_l274_7 == 7'h0);
  assign outputStreamArrayData_7_fire_9 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l275_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l275_7) && outputStreamArrayData_7_fire_9);
  assign _zz_realValue1_0_46 = (_zz__zz_realValue1_0_46 % _zz__zz_realValue1_0_46_1);
  assign when_ArraySlice_l95_46 = (_zz_realValue1_0_46 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_46) begin
      realValue1_0_46 = (_zz_realValue1_0_46_1 - _zz_realValue1_0_46);
    end else begin
      realValue1_0_46 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l277_7 = (_zz_when_ArraySlice_l277_7 < _zz_when_ArraySlice_l277_7_2);
  always @(*) begin
    debug_0_48 = 1'b0;
    if(when_ArraySlice_l158_384) begin
      if(when_ArraySlice_l159_384) begin
        debug_0_48 = 1'b1;
      end else begin
        debug_0_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_384) begin
        debug_0_48 = 1'b1;
      end else begin
        debug_0_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_48 = 1'b0;
    if(when_ArraySlice_l158_385) begin
      if(when_ArraySlice_l159_385) begin
        debug_1_48 = 1'b1;
      end else begin
        debug_1_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_385) begin
        debug_1_48 = 1'b1;
      end else begin
        debug_1_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_48 = 1'b0;
    if(when_ArraySlice_l158_386) begin
      if(when_ArraySlice_l159_386) begin
        debug_2_48 = 1'b1;
      end else begin
        debug_2_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_386) begin
        debug_2_48 = 1'b1;
      end else begin
        debug_2_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_48 = 1'b0;
    if(when_ArraySlice_l158_387) begin
      if(when_ArraySlice_l159_387) begin
        debug_3_48 = 1'b1;
      end else begin
        debug_3_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_387) begin
        debug_3_48 = 1'b1;
      end else begin
        debug_3_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_48 = 1'b0;
    if(when_ArraySlice_l158_388) begin
      if(when_ArraySlice_l159_388) begin
        debug_4_48 = 1'b1;
      end else begin
        debug_4_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_388) begin
        debug_4_48 = 1'b1;
      end else begin
        debug_4_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_48 = 1'b0;
    if(when_ArraySlice_l158_389) begin
      if(when_ArraySlice_l159_389) begin
        debug_5_48 = 1'b1;
      end else begin
        debug_5_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_389) begin
        debug_5_48 = 1'b1;
      end else begin
        debug_5_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_48 = 1'b0;
    if(when_ArraySlice_l158_390) begin
      if(when_ArraySlice_l159_390) begin
        debug_6_48 = 1'b1;
      end else begin
        debug_6_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_390) begin
        debug_6_48 = 1'b1;
      end else begin
        debug_6_48 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_48 = 1'b0;
    if(when_ArraySlice_l158_391) begin
      if(when_ArraySlice_l159_391) begin
        debug_7_48 = 1'b1;
      end else begin
        debug_7_48 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_391) begin
        debug_7_48 = 1'b1;
      end else begin
        debug_7_48 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_384 = (_zz_when_ArraySlice_l158_384 <= _zz_when_ArraySlice_l158_384_3);
  assign when_ArraySlice_l159_384 = (_zz_when_ArraySlice_l159_384 <= _zz_when_ArraySlice_l159_384_1);
  assign _zz_realValue_0_384 = (_zz__zz_realValue_0_384 % _zz__zz_realValue_0_384_1);
  assign when_ArraySlice_l110_384 = (_zz_realValue_0_384 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_384) begin
      realValue_0_384 = (_zz_realValue_0_384_1 - _zz_realValue_0_384);
    end else begin
      realValue_0_384 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_384 = (_zz_when_ArraySlice_l166_384 <= _zz_when_ArraySlice_l166_384_1);
  assign when_ArraySlice_l158_385 = (_zz_when_ArraySlice_l158_385 <= _zz_when_ArraySlice_l158_385_3);
  assign when_ArraySlice_l159_385 = (_zz_when_ArraySlice_l159_385 <= _zz_when_ArraySlice_l159_385_2);
  assign _zz_realValue_0_385 = (_zz__zz_realValue_0_385 % _zz__zz_realValue_0_385_1);
  assign when_ArraySlice_l110_385 = (_zz_realValue_0_385 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_385) begin
      realValue_0_385 = (_zz_realValue_0_385_1 - _zz_realValue_0_385);
    end else begin
      realValue_0_385 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_385 = (_zz_when_ArraySlice_l166_385 <= _zz_when_ArraySlice_l166_385_2);
  assign when_ArraySlice_l158_386 = (_zz_when_ArraySlice_l158_386 <= _zz_when_ArraySlice_l158_386_3);
  assign when_ArraySlice_l159_386 = (_zz_when_ArraySlice_l159_386 <= _zz_when_ArraySlice_l159_386_2);
  assign _zz_realValue_0_386 = (_zz__zz_realValue_0_386 % _zz__zz_realValue_0_386_1);
  assign when_ArraySlice_l110_386 = (_zz_realValue_0_386 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_386) begin
      realValue_0_386 = (_zz_realValue_0_386_1 - _zz_realValue_0_386);
    end else begin
      realValue_0_386 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_386 = (_zz_when_ArraySlice_l166_386 <= _zz_when_ArraySlice_l166_386_2);
  assign when_ArraySlice_l158_387 = (_zz_when_ArraySlice_l158_387 <= _zz_when_ArraySlice_l158_387_3);
  assign when_ArraySlice_l159_387 = (_zz_when_ArraySlice_l159_387 <= _zz_when_ArraySlice_l159_387_2);
  assign _zz_realValue_0_387 = (_zz__zz_realValue_0_387 % _zz__zz_realValue_0_387_1);
  assign when_ArraySlice_l110_387 = (_zz_realValue_0_387 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_387) begin
      realValue_0_387 = (_zz_realValue_0_387_1 - _zz_realValue_0_387);
    end else begin
      realValue_0_387 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_387 = (_zz_when_ArraySlice_l166_387 <= _zz_when_ArraySlice_l166_387_2);
  assign when_ArraySlice_l158_388 = (_zz_when_ArraySlice_l158_388 <= _zz_when_ArraySlice_l158_388_3);
  assign when_ArraySlice_l159_388 = (_zz_when_ArraySlice_l159_388 <= _zz_when_ArraySlice_l159_388_2);
  assign _zz_realValue_0_388 = (_zz__zz_realValue_0_388 % _zz__zz_realValue_0_388_1);
  assign when_ArraySlice_l110_388 = (_zz_realValue_0_388 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_388) begin
      realValue_0_388 = (_zz_realValue_0_388_1 - _zz_realValue_0_388);
    end else begin
      realValue_0_388 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_388 = (_zz_when_ArraySlice_l166_388 <= _zz_when_ArraySlice_l166_388_2);
  assign when_ArraySlice_l158_389 = (_zz_when_ArraySlice_l158_389 <= _zz_when_ArraySlice_l158_389_3);
  assign when_ArraySlice_l159_389 = (_zz_when_ArraySlice_l159_389 <= _zz_when_ArraySlice_l159_389_2);
  assign _zz_realValue_0_389 = (_zz__zz_realValue_0_389 % _zz__zz_realValue_0_389_1);
  assign when_ArraySlice_l110_389 = (_zz_realValue_0_389 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_389) begin
      realValue_0_389 = (_zz_realValue_0_389_1 - _zz_realValue_0_389);
    end else begin
      realValue_0_389 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_389 = (_zz_when_ArraySlice_l166_389 <= _zz_when_ArraySlice_l166_389_2);
  assign when_ArraySlice_l158_390 = (_zz_when_ArraySlice_l158_390 <= _zz_when_ArraySlice_l158_390_3);
  assign when_ArraySlice_l159_390 = (_zz_when_ArraySlice_l159_390 <= _zz_when_ArraySlice_l159_390_2);
  assign _zz_realValue_0_390 = (_zz__zz_realValue_0_390 % _zz__zz_realValue_0_390_1);
  assign when_ArraySlice_l110_390 = (_zz_realValue_0_390 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_390) begin
      realValue_0_390 = (_zz_realValue_0_390_1 - _zz_realValue_0_390);
    end else begin
      realValue_0_390 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_390 = (_zz_when_ArraySlice_l166_390 <= _zz_when_ArraySlice_l166_390_2);
  assign when_ArraySlice_l158_391 = (_zz_when_ArraySlice_l158_391 <= _zz_when_ArraySlice_l158_391_3);
  assign when_ArraySlice_l159_391 = (_zz_when_ArraySlice_l159_391 <= _zz_when_ArraySlice_l159_391_2);
  assign _zz_realValue_0_391 = (_zz__zz_realValue_0_391 % _zz__zz_realValue_0_391_1);
  assign when_ArraySlice_l110_391 = (_zz_realValue_0_391 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_391) begin
      realValue_0_391 = (_zz_realValue_0_391_1 - _zz_realValue_0_391);
    end else begin
      realValue_0_391 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_391 = (_zz_when_ArraySlice_l166_391 <= _zz_when_ArraySlice_l166_391_2);
  assign when_ArraySlice_l282_7 = (! ((((((_zz_when_ArraySlice_l282_7 && _zz_when_ArraySlice_l282_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l282_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l282_7_3 && _zz_when_ArraySlice_l282_7_4) && (debug_4_48 == _zz_when_ArraySlice_l282_7_5)) && (debug_5_48 == 1'b1)) && (debug_6_48 == 1'b1)) && (debug_7_48 == 1'b1))));
  assign when_ArraySlice_l285_7 = (_zz_when_ArraySlice_l285_7_1 <= _zz_when_ArraySlice_l285_7_2);
  assign when_ArraySlice_l288_7 = (_zz_when_ArraySlice_l288_7 <= _zz_when_ArraySlice_l288_7_1);
  assign outputStreamArrayData_7_fire_10 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l295_7 = ((_zz_when_ArraySlice_l295_7 == 13'h0) && outputStreamArrayData_7_fire_10);
  assign outputStreamArrayData_7_fire_11 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l306_7 = ((handshakeTimes_7_value == _zz_when_ArraySlice_l306_7) && outputStreamArrayData_7_fire_11);
  assign _zz_realValue1_0_47 = (_zz__zz_realValue1_0_47 % _zz__zz_realValue1_0_47_1);
  assign when_ArraySlice_l95_47 = (_zz_realValue1_0_47 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l95_47) begin
      realValue1_0_47 = (_zz_realValue1_0_47_1 - _zz_realValue1_0_47);
    end else begin
      realValue1_0_47 = {1'd0, hReg};
    end
  end

  assign when_ArraySlice_l307_7 = (_zz_when_ArraySlice_l307_7 < _zz_when_ArraySlice_l307_7_2);
  always @(*) begin
    debug_0_49 = 1'b0;
    if(when_ArraySlice_l158_392) begin
      if(when_ArraySlice_l159_392) begin
        debug_0_49 = 1'b1;
      end else begin
        debug_0_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_392) begin
        debug_0_49 = 1'b1;
      end else begin
        debug_0_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_49 = 1'b0;
    if(when_ArraySlice_l158_393) begin
      if(when_ArraySlice_l159_393) begin
        debug_1_49 = 1'b1;
      end else begin
        debug_1_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_393) begin
        debug_1_49 = 1'b1;
      end else begin
        debug_1_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_49 = 1'b0;
    if(when_ArraySlice_l158_394) begin
      if(when_ArraySlice_l159_394) begin
        debug_2_49 = 1'b1;
      end else begin
        debug_2_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_394) begin
        debug_2_49 = 1'b1;
      end else begin
        debug_2_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_49 = 1'b0;
    if(when_ArraySlice_l158_395) begin
      if(when_ArraySlice_l159_395) begin
        debug_3_49 = 1'b1;
      end else begin
        debug_3_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_395) begin
        debug_3_49 = 1'b1;
      end else begin
        debug_3_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_49 = 1'b0;
    if(when_ArraySlice_l158_396) begin
      if(when_ArraySlice_l159_396) begin
        debug_4_49 = 1'b1;
      end else begin
        debug_4_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_396) begin
        debug_4_49 = 1'b1;
      end else begin
        debug_4_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_49 = 1'b0;
    if(when_ArraySlice_l158_397) begin
      if(when_ArraySlice_l159_397) begin
        debug_5_49 = 1'b1;
      end else begin
        debug_5_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_397) begin
        debug_5_49 = 1'b1;
      end else begin
        debug_5_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_49 = 1'b0;
    if(when_ArraySlice_l158_398) begin
      if(when_ArraySlice_l159_398) begin
        debug_6_49 = 1'b1;
      end else begin
        debug_6_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_398) begin
        debug_6_49 = 1'b1;
      end else begin
        debug_6_49 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_49 = 1'b0;
    if(when_ArraySlice_l158_399) begin
      if(when_ArraySlice_l159_399) begin
        debug_7_49 = 1'b1;
      end else begin
        debug_7_49 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_399) begin
        debug_7_49 = 1'b1;
      end else begin
        debug_7_49 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_392 = (_zz_when_ArraySlice_l158_392 <= _zz_when_ArraySlice_l158_392_3);
  assign when_ArraySlice_l159_392 = (_zz_when_ArraySlice_l159_392 <= _zz_when_ArraySlice_l159_392_1);
  assign _zz_realValue_0_392 = (_zz__zz_realValue_0_392 % _zz__zz_realValue_0_392_1);
  assign when_ArraySlice_l110_392 = (_zz_realValue_0_392 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_392) begin
      realValue_0_392 = (_zz_realValue_0_392_1 - _zz_realValue_0_392);
    end else begin
      realValue_0_392 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_392 = (_zz_when_ArraySlice_l166_392 <= _zz_when_ArraySlice_l166_392_1);
  assign when_ArraySlice_l158_393 = (_zz_when_ArraySlice_l158_393 <= _zz_when_ArraySlice_l158_393_3);
  assign when_ArraySlice_l159_393 = (_zz_when_ArraySlice_l159_393 <= _zz_when_ArraySlice_l159_393_2);
  assign _zz_realValue_0_393 = (_zz__zz_realValue_0_393 % _zz__zz_realValue_0_393_1);
  assign when_ArraySlice_l110_393 = (_zz_realValue_0_393 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_393) begin
      realValue_0_393 = (_zz_realValue_0_393_1 - _zz_realValue_0_393);
    end else begin
      realValue_0_393 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_393 = (_zz_when_ArraySlice_l166_393 <= _zz_when_ArraySlice_l166_393_2);
  assign when_ArraySlice_l158_394 = (_zz_when_ArraySlice_l158_394 <= _zz_when_ArraySlice_l158_394_3);
  assign when_ArraySlice_l159_394 = (_zz_when_ArraySlice_l159_394 <= _zz_when_ArraySlice_l159_394_2);
  assign _zz_realValue_0_394 = (_zz__zz_realValue_0_394 % _zz__zz_realValue_0_394_1);
  assign when_ArraySlice_l110_394 = (_zz_realValue_0_394 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_394) begin
      realValue_0_394 = (_zz_realValue_0_394_1 - _zz_realValue_0_394);
    end else begin
      realValue_0_394 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_394 = (_zz_when_ArraySlice_l166_394 <= _zz_when_ArraySlice_l166_394_2);
  assign when_ArraySlice_l158_395 = (_zz_when_ArraySlice_l158_395 <= _zz_when_ArraySlice_l158_395_3);
  assign when_ArraySlice_l159_395 = (_zz_when_ArraySlice_l159_395 <= _zz_when_ArraySlice_l159_395_2);
  assign _zz_realValue_0_395 = (_zz__zz_realValue_0_395 % _zz__zz_realValue_0_395_1);
  assign when_ArraySlice_l110_395 = (_zz_realValue_0_395 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_395) begin
      realValue_0_395 = (_zz_realValue_0_395_1 - _zz_realValue_0_395);
    end else begin
      realValue_0_395 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_395 = (_zz_when_ArraySlice_l166_395 <= _zz_when_ArraySlice_l166_395_2);
  assign when_ArraySlice_l158_396 = (_zz_when_ArraySlice_l158_396 <= _zz_when_ArraySlice_l158_396_3);
  assign when_ArraySlice_l159_396 = (_zz_when_ArraySlice_l159_396 <= _zz_when_ArraySlice_l159_396_2);
  assign _zz_realValue_0_396 = (_zz__zz_realValue_0_396 % _zz__zz_realValue_0_396_1);
  assign when_ArraySlice_l110_396 = (_zz_realValue_0_396 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_396) begin
      realValue_0_396 = (_zz_realValue_0_396_1 - _zz_realValue_0_396);
    end else begin
      realValue_0_396 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_396 = (_zz_when_ArraySlice_l166_396 <= _zz_when_ArraySlice_l166_396_2);
  assign when_ArraySlice_l158_397 = (_zz_when_ArraySlice_l158_397 <= _zz_when_ArraySlice_l158_397_3);
  assign when_ArraySlice_l159_397 = (_zz_when_ArraySlice_l159_397 <= _zz_when_ArraySlice_l159_397_2);
  assign _zz_realValue_0_397 = (_zz__zz_realValue_0_397 % _zz__zz_realValue_0_397_1);
  assign when_ArraySlice_l110_397 = (_zz_realValue_0_397 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_397) begin
      realValue_0_397 = (_zz_realValue_0_397_1 - _zz_realValue_0_397);
    end else begin
      realValue_0_397 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_397 = (_zz_when_ArraySlice_l166_397 <= _zz_when_ArraySlice_l166_397_2);
  assign when_ArraySlice_l158_398 = (_zz_when_ArraySlice_l158_398 <= _zz_when_ArraySlice_l158_398_3);
  assign when_ArraySlice_l159_398 = (_zz_when_ArraySlice_l159_398 <= _zz_when_ArraySlice_l159_398_2);
  assign _zz_realValue_0_398 = (_zz__zz_realValue_0_398 % _zz__zz_realValue_0_398_1);
  assign when_ArraySlice_l110_398 = (_zz_realValue_0_398 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_398) begin
      realValue_0_398 = (_zz_realValue_0_398_1 - _zz_realValue_0_398);
    end else begin
      realValue_0_398 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_398 = (_zz_when_ArraySlice_l166_398 <= _zz_when_ArraySlice_l166_398_2);
  assign when_ArraySlice_l158_399 = (_zz_when_ArraySlice_l158_399 <= _zz_when_ArraySlice_l158_399_3);
  assign when_ArraySlice_l159_399 = (_zz_when_ArraySlice_l159_399 <= _zz_when_ArraySlice_l159_399_2);
  assign _zz_realValue_0_399 = (_zz__zz_realValue_0_399 % _zz__zz_realValue_0_399_1);
  assign when_ArraySlice_l110_399 = (_zz_realValue_0_399 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_399) begin
      realValue_0_399 = (_zz_realValue_0_399_1 - _zz_realValue_0_399);
    end else begin
      realValue_0_399 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_399 = (_zz_when_ArraySlice_l166_399 <= _zz_when_ArraySlice_l166_399_2);
  assign when_ArraySlice_l314_7 = (! ((((((_zz_when_ArraySlice_l314_7 && _zz_when_ArraySlice_l314_7_1) && (holdReadOp_4 == _zz_when_ArraySlice_l314_7_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l314_7_3 && _zz_when_ArraySlice_l314_7_4) && (debug_4_49 == _zz_when_ArraySlice_l314_7_5)) && (debug_5_49 == 1'b1)) && (debug_6_49 == 1'b1)) && (debug_7_49 == 1'b1))));
  assign outputStreamArrayData_7_fire_12 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l318_7 = ((_zz_when_ArraySlice_l318_7 == 13'h0) && outputStreamArrayData_7_fire_12);
  assign when_ArraySlice_l304_7 = (allowPadding_7 && (_zz_when_ArraySlice_l304_7 <= _zz_when_ArraySlice_l304_7_1));
  assign outputStreamArrayData_7_fire_13 = (outputStreamArrayData_7_valid && outputStreamArrayData_7_ready);
  assign when_ArraySlice_l325_7 = (handshakeTimes_7_value == _zz_when_ArraySlice_l325_7);
  assign when_ArraySlice_l182 = (_zz_when_ArraySlice_l182 == _zz_when_ArraySlice_l182_1);
  assign when_ArraySlice_l183 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l182) begin
      if(when_ArraySlice_l183) begin
        _zz_when_ArraySlice_l336 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_1 = (_zz_when_ArraySlice_l182_1_1 == _zz_when_ArraySlice_l182_1_2);
  assign when_ArraySlice_l183_1 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l182_1) begin
      if(when_ArraySlice_l183_1) begin
        _zz_when_ArraySlice_l336_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_2 = (_zz_when_ArraySlice_l182_2_1 == _zz_when_ArraySlice_l182_2_2);
  assign when_ArraySlice_l183_2 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l182_2) begin
      if(when_ArraySlice_l183_2) begin
        _zz_when_ArraySlice_l336_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_3 = (_zz_when_ArraySlice_l182_3 == _zz_when_ArraySlice_l182_3_1);
  assign when_ArraySlice_l183_3 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l182_3) begin
      if(when_ArraySlice_l183_3) begin
        _zz_when_ArraySlice_l336_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_4 = (_zz_when_ArraySlice_l182_4 == _zz_when_ArraySlice_l182_4_1);
  assign when_ArraySlice_l183_4 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l182_4) begin
      if(when_ArraySlice_l183_4) begin
        _zz_when_ArraySlice_l336_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_5 = (_zz_when_ArraySlice_l182_5 == _zz_when_ArraySlice_l182_5_1);
  assign when_ArraySlice_l183_5 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l182_5) begin
      if(when_ArraySlice_l183_5) begin
        _zz_when_ArraySlice_l336_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_6 = (_zz_when_ArraySlice_l182_6 == _zz_when_ArraySlice_l182_6_1);
  assign when_ArraySlice_l183_6 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l182_6) begin
      if(when_ArraySlice_l183_6) begin
        _zz_when_ArraySlice_l336_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_7 = (_zz_when_ArraySlice_l182_7 == _zz_when_ArraySlice_l182_7_1);
  assign when_ArraySlice_l183_7 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l182_7) begin
      if(when_ArraySlice_l183_7) begin
        _zz_when_ArraySlice_l336_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l336_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l336_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l336 = (! ((((((((_zz_when_ArraySlice_l336 != _zz_when_ArraySlice_l336_8) || (_zz_when_ArraySlice_l336_1 != _zz_when_ArraySlice_l336_9)) || (_zz_when_ArraySlice_l336_2 != 1'b0)) || (_zz_when_ArraySlice_l336_3 != 1'b0)) || (_zz_when_ArraySlice_l336_4 != 1'b0)) || (_zz_when_ArraySlice_l336_5 != 1'b0)) || (_zz_when_ArraySlice_l336_6 != 1'b0)) || (_zz_when_ArraySlice_l336_7 != 1'b0)));
  assign when_ArraySlice_l337 = (_zz_when_ArraySlice_l337 < hReg);
  assign _zz_19 = ({127'd0,1'b1} <<< selectWriteFifo);
  assign _zz_20 = ({127'd0,1'b1} <<< selectWriteFifo);
  assign _zz_io_push_valid_1 = inputStreamArrayData_valid;
  assign _zz_io_push_payload_1 = inputStreamArrayData_payload;
  assign inputStreamArrayData_fire_1 = (inputStreamArrayData_valid && inputStreamArrayData_ready);
  assign when_ArraySlice_l341 = ((_zz_when_ArraySlice_l341 == _zz_when_ArraySlice_l341_1) && inputStreamArrayData_fire_1);
  assign when_ArraySlice_l342 = (selectWriteFifo == _zz_when_ArraySlice_l342);
  always @(*) begin
    debug_0_50 = 1'b0;
    if(when_ArraySlice_l158_400) begin
      if(when_ArraySlice_l159_400) begin
        debug_0_50 = 1'b1;
      end else begin
        debug_0_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_400) begin
        debug_0_50 = 1'b1;
      end else begin
        debug_0_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_50 = 1'b0;
    if(when_ArraySlice_l158_401) begin
      if(when_ArraySlice_l159_401) begin
        debug_1_50 = 1'b1;
      end else begin
        debug_1_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_401) begin
        debug_1_50 = 1'b1;
      end else begin
        debug_1_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_50 = 1'b0;
    if(when_ArraySlice_l158_402) begin
      if(when_ArraySlice_l159_402) begin
        debug_2_50 = 1'b1;
      end else begin
        debug_2_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_402) begin
        debug_2_50 = 1'b1;
      end else begin
        debug_2_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_50 = 1'b0;
    if(when_ArraySlice_l158_403) begin
      if(when_ArraySlice_l159_403) begin
        debug_3_50 = 1'b1;
      end else begin
        debug_3_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_403) begin
        debug_3_50 = 1'b1;
      end else begin
        debug_3_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_50 = 1'b0;
    if(when_ArraySlice_l158_404) begin
      if(when_ArraySlice_l159_404) begin
        debug_4_50 = 1'b1;
      end else begin
        debug_4_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_404) begin
        debug_4_50 = 1'b1;
      end else begin
        debug_4_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_50 = 1'b0;
    if(when_ArraySlice_l158_405) begin
      if(when_ArraySlice_l159_405) begin
        debug_5_50 = 1'b1;
      end else begin
        debug_5_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_405) begin
        debug_5_50 = 1'b1;
      end else begin
        debug_5_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_50 = 1'b0;
    if(when_ArraySlice_l158_406) begin
      if(when_ArraySlice_l159_406) begin
        debug_6_50 = 1'b1;
      end else begin
        debug_6_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_406) begin
        debug_6_50 = 1'b1;
      end else begin
        debug_6_50 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_50 = 1'b0;
    if(when_ArraySlice_l158_407) begin
      if(when_ArraySlice_l159_407) begin
        debug_7_50 = 1'b1;
      end else begin
        debug_7_50 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_407) begin
        debug_7_50 = 1'b1;
      end else begin
        debug_7_50 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_400 = (_zz_when_ArraySlice_l158_400 <= _zz_when_ArraySlice_l158_400_3);
  assign when_ArraySlice_l159_400 = (_zz_when_ArraySlice_l159_400 <= _zz_when_ArraySlice_l159_400_1);
  assign _zz_realValue_0_400 = (_zz__zz_realValue_0_400 % _zz__zz_realValue_0_400_1);
  assign when_ArraySlice_l110_400 = (_zz_realValue_0_400 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_400) begin
      realValue_0_400 = (_zz_realValue_0_400_1 - _zz_realValue_0_400);
    end else begin
      realValue_0_400 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_400 = (_zz_when_ArraySlice_l166_400 <= _zz_when_ArraySlice_l166_400_1);
  assign when_ArraySlice_l158_401 = (_zz_when_ArraySlice_l158_401 <= _zz_when_ArraySlice_l158_401_3);
  assign when_ArraySlice_l159_401 = (_zz_when_ArraySlice_l159_401 <= _zz_when_ArraySlice_l159_401_2);
  assign _zz_realValue_0_401 = (_zz__zz_realValue_0_401 % _zz__zz_realValue_0_401_1);
  assign when_ArraySlice_l110_401 = (_zz_realValue_0_401 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_401) begin
      realValue_0_401 = (_zz_realValue_0_401_1 - _zz_realValue_0_401);
    end else begin
      realValue_0_401 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_401 = (_zz_when_ArraySlice_l166_401 <= _zz_when_ArraySlice_l166_401_2);
  assign when_ArraySlice_l158_402 = (_zz_when_ArraySlice_l158_402 <= _zz_when_ArraySlice_l158_402_3);
  assign when_ArraySlice_l159_402 = (_zz_when_ArraySlice_l159_402 <= _zz_when_ArraySlice_l159_402_2);
  assign _zz_realValue_0_402 = (_zz__zz_realValue_0_402 % _zz__zz_realValue_0_402_1);
  assign when_ArraySlice_l110_402 = (_zz_realValue_0_402 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_402) begin
      realValue_0_402 = (_zz_realValue_0_402_1 - _zz_realValue_0_402);
    end else begin
      realValue_0_402 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_402 = (_zz_when_ArraySlice_l166_402 <= _zz_when_ArraySlice_l166_402_2);
  assign when_ArraySlice_l158_403 = (_zz_when_ArraySlice_l158_403 <= _zz_when_ArraySlice_l158_403_3);
  assign when_ArraySlice_l159_403 = (_zz_when_ArraySlice_l159_403 <= _zz_when_ArraySlice_l159_403_2);
  assign _zz_realValue_0_403 = (_zz__zz_realValue_0_403 % _zz__zz_realValue_0_403_1);
  assign when_ArraySlice_l110_403 = (_zz_realValue_0_403 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_403) begin
      realValue_0_403 = (_zz_realValue_0_403_1 - _zz_realValue_0_403);
    end else begin
      realValue_0_403 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_403 = (_zz_when_ArraySlice_l166_403 <= _zz_when_ArraySlice_l166_403_2);
  assign when_ArraySlice_l158_404 = (_zz_when_ArraySlice_l158_404 <= _zz_when_ArraySlice_l158_404_3);
  assign when_ArraySlice_l159_404 = (_zz_when_ArraySlice_l159_404 <= _zz_when_ArraySlice_l159_404_2);
  assign _zz_realValue_0_404 = (_zz__zz_realValue_0_404 % _zz__zz_realValue_0_404_1);
  assign when_ArraySlice_l110_404 = (_zz_realValue_0_404 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_404) begin
      realValue_0_404 = (_zz_realValue_0_404_1 - _zz_realValue_0_404);
    end else begin
      realValue_0_404 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_404 = (_zz_when_ArraySlice_l166_404 <= _zz_when_ArraySlice_l166_404_2);
  assign when_ArraySlice_l158_405 = (_zz_when_ArraySlice_l158_405 <= _zz_when_ArraySlice_l158_405_3);
  assign when_ArraySlice_l159_405 = (_zz_when_ArraySlice_l159_405 <= _zz_when_ArraySlice_l159_405_2);
  assign _zz_realValue_0_405 = (_zz__zz_realValue_0_405 % _zz__zz_realValue_0_405_1);
  assign when_ArraySlice_l110_405 = (_zz_realValue_0_405 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_405) begin
      realValue_0_405 = (_zz_realValue_0_405_1 - _zz_realValue_0_405);
    end else begin
      realValue_0_405 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_405 = (_zz_when_ArraySlice_l166_405 <= _zz_when_ArraySlice_l166_405_2);
  assign when_ArraySlice_l158_406 = (_zz_when_ArraySlice_l158_406 <= _zz_when_ArraySlice_l158_406_3);
  assign when_ArraySlice_l159_406 = (_zz_when_ArraySlice_l159_406 <= _zz_when_ArraySlice_l159_406_2);
  assign _zz_realValue_0_406 = (_zz__zz_realValue_0_406 % _zz__zz_realValue_0_406_1);
  assign when_ArraySlice_l110_406 = (_zz_realValue_0_406 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_406) begin
      realValue_0_406 = (_zz_realValue_0_406_1 - _zz_realValue_0_406);
    end else begin
      realValue_0_406 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_406 = (_zz_when_ArraySlice_l166_406 <= _zz_when_ArraySlice_l166_406_2);
  assign when_ArraySlice_l158_407 = (_zz_when_ArraySlice_l158_407 <= _zz_when_ArraySlice_l158_407_3);
  assign when_ArraySlice_l159_407 = (_zz_when_ArraySlice_l159_407 <= _zz_when_ArraySlice_l159_407_2);
  assign _zz_realValue_0_407 = (_zz__zz_realValue_0_407 % _zz__zz_realValue_0_407_1);
  assign when_ArraySlice_l110_407 = (_zz_realValue_0_407 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_407) begin
      realValue_0_407 = (_zz_realValue_0_407_1 - _zz_realValue_0_407);
    end else begin
      realValue_0_407 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_407 = (_zz_when_ArraySlice_l166_407 <= _zz_when_ArraySlice_l166_407_2);
  assign when_ArraySlice_l353 = ((((((_zz_when_ArraySlice_l353 && _zz_when_ArraySlice_l353_1) && (holdReadOp_4 == _zz_when_ArraySlice_l353_2)) && (holdReadOp_5 == 1'b1)) && (holdReadOp_6 == 1'b1)) && (holdReadOp_7 == 1'b1)) && (((((_zz_when_ArraySlice_l353_3 && _zz_when_ArraySlice_l353_4) && (debug_4_50 == _zz_when_ArraySlice_l353_5)) && (debug_5_50 == 1'b1)) && (debug_6_50 == 1'b1)) && (debug_7_50 == 1'b1)));
  always @(*) begin
    debug_0_51 = 1'b0;
    if(when_ArraySlice_l158_408) begin
      if(when_ArraySlice_l159_408) begin
        debug_0_51 = 1'b1;
      end else begin
        debug_0_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_408) begin
        debug_0_51 = 1'b1;
      end else begin
        debug_0_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_1_51 = 1'b0;
    if(when_ArraySlice_l158_409) begin
      if(when_ArraySlice_l159_409) begin
        debug_1_51 = 1'b1;
      end else begin
        debug_1_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_409) begin
        debug_1_51 = 1'b1;
      end else begin
        debug_1_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_2_51 = 1'b0;
    if(when_ArraySlice_l158_410) begin
      if(when_ArraySlice_l159_410) begin
        debug_2_51 = 1'b1;
      end else begin
        debug_2_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_410) begin
        debug_2_51 = 1'b1;
      end else begin
        debug_2_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_3_51 = 1'b0;
    if(when_ArraySlice_l158_411) begin
      if(when_ArraySlice_l159_411) begin
        debug_3_51 = 1'b1;
      end else begin
        debug_3_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_411) begin
        debug_3_51 = 1'b1;
      end else begin
        debug_3_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_4_51 = 1'b0;
    if(when_ArraySlice_l158_412) begin
      if(when_ArraySlice_l159_412) begin
        debug_4_51 = 1'b1;
      end else begin
        debug_4_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_412) begin
        debug_4_51 = 1'b1;
      end else begin
        debug_4_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_5_51 = 1'b0;
    if(when_ArraySlice_l158_413) begin
      if(when_ArraySlice_l159_413) begin
        debug_5_51 = 1'b1;
      end else begin
        debug_5_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_413) begin
        debug_5_51 = 1'b1;
      end else begin
        debug_5_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_6_51 = 1'b0;
    if(when_ArraySlice_l158_414) begin
      if(when_ArraySlice_l159_414) begin
        debug_6_51 = 1'b1;
      end else begin
        debug_6_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_414) begin
        debug_6_51 = 1'b1;
      end else begin
        debug_6_51 = 1'b0;
      end
    end
  end

  always @(*) begin
    debug_7_51 = 1'b0;
    if(when_ArraySlice_l158_415) begin
      if(when_ArraySlice_l159_415) begin
        debug_7_51 = 1'b1;
      end else begin
        debug_7_51 = 1'b0;
      end
    end else begin
      if(when_ArraySlice_l166_415) begin
        debug_7_51 = 1'b1;
      end else begin
        debug_7_51 = 1'b0;
      end
    end
  end

  assign when_ArraySlice_l158_408 = (_zz_when_ArraySlice_l158_408 <= _zz_when_ArraySlice_l158_408_3);
  assign when_ArraySlice_l159_408 = (_zz_when_ArraySlice_l159_408 <= _zz_when_ArraySlice_l159_408_1);
  assign _zz_realValue_0_408 = (_zz__zz_realValue_0_408 % _zz__zz_realValue_0_408_1);
  assign when_ArraySlice_l110_408 = (_zz_realValue_0_408 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_408) begin
      realValue_0_408 = (_zz_realValue_0_408_1 - _zz_realValue_0_408);
    end else begin
      realValue_0_408 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_408 = (_zz_when_ArraySlice_l166_408 <= _zz_when_ArraySlice_l166_408_1);
  assign when_ArraySlice_l158_409 = (_zz_when_ArraySlice_l158_409 <= _zz_when_ArraySlice_l158_409_3);
  assign when_ArraySlice_l159_409 = (_zz_when_ArraySlice_l159_409 <= _zz_when_ArraySlice_l159_409_2);
  assign _zz_realValue_0_409 = (_zz__zz_realValue_0_409 % _zz__zz_realValue_0_409_1);
  assign when_ArraySlice_l110_409 = (_zz_realValue_0_409 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_409) begin
      realValue_0_409 = (_zz_realValue_0_409_1 - _zz_realValue_0_409);
    end else begin
      realValue_0_409 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_409 = (_zz_when_ArraySlice_l166_409 <= _zz_when_ArraySlice_l166_409_2);
  assign when_ArraySlice_l158_410 = (_zz_when_ArraySlice_l158_410 <= _zz_when_ArraySlice_l158_410_3);
  assign when_ArraySlice_l159_410 = (_zz_when_ArraySlice_l159_410 <= _zz_when_ArraySlice_l159_410_2);
  assign _zz_realValue_0_410 = (_zz__zz_realValue_0_410 % _zz__zz_realValue_0_410_1);
  assign when_ArraySlice_l110_410 = (_zz_realValue_0_410 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_410) begin
      realValue_0_410 = (_zz_realValue_0_410_1 - _zz_realValue_0_410);
    end else begin
      realValue_0_410 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_410 = (_zz_when_ArraySlice_l166_410 <= _zz_when_ArraySlice_l166_410_2);
  assign when_ArraySlice_l158_411 = (_zz_when_ArraySlice_l158_411 <= _zz_when_ArraySlice_l158_411_3);
  assign when_ArraySlice_l159_411 = (_zz_when_ArraySlice_l159_411 <= _zz_when_ArraySlice_l159_411_2);
  assign _zz_realValue_0_411 = (_zz__zz_realValue_0_411 % _zz__zz_realValue_0_411_1);
  assign when_ArraySlice_l110_411 = (_zz_realValue_0_411 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_411) begin
      realValue_0_411 = (_zz_realValue_0_411_1 - _zz_realValue_0_411);
    end else begin
      realValue_0_411 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_411 = (_zz_when_ArraySlice_l166_411 <= _zz_when_ArraySlice_l166_411_2);
  assign when_ArraySlice_l158_412 = (_zz_when_ArraySlice_l158_412 <= _zz_when_ArraySlice_l158_412_3);
  assign when_ArraySlice_l159_412 = (_zz_when_ArraySlice_l159_412 <= _zz_when_ArraySlice_l159_412_2);
  assign _zz_realValue_0_412 = (_zz__zz_realValue_0_412 % _zz__zz_realValue_0_412_1);
  assign when_ArraySlice_l110_412 = (_zz_realValue_0_412 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_412) begin
      realValue_0_412 = (_zz_realValue_0_412_1 - _zz_realValue_0_412);
    end else begin
      realValue_0_412 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_412 = (_zz_when_ArraySlice_l166_412 <= _zz_when_ArraySlice_l166_412_2);
  assign when_ArraySlice_l158_413 = (_zz_when_ArraySlice_l158_413 <= _zz_when_ArraySlice_l158_413_3);
  assign when_ArraySlice_l159_413 = (_zz_when_ArraySlice_l159_413 <= _zz_when_ArraySlice_l159_413_2);
  assign _zz_realValue_0_413 = (_zz__zz_realValue_0_413 % _zz__zz_realValue_0_413_1);
  assign when_ArraySlice_l110_413 = (_zz_realValue_0_413 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_413) begin
      realValue_0_413 = (_zz_realValue_0_413_1 - _zz_realValue_0_413);
    end else begin
      realValue_0_413 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_413 = (_zz_when_ArraySlice_l166_413 <= _zz_when_ArraySlice_l166_413_2);
  assign when_ArraySlice_l158_414 = (_zz_when_ArraySlice_l158_414 <= _zz_when_ArraySlice_l158_414_3);
  assign when_ArraySlice_l159_414 = (_zz_when_ArraySlice_l159_414 <= _zz_when_ArraySlice_l159_414_2);
  assign _zz_realValue_0_414 = (_zz__zz_realValue_0_414 % _zz__zz_realValue_0_414_1);
  assign when_ArraySlice_l110_414 = (_zz_realValue_0_414 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_414) begin
      realValue_0_414 = (_zz_realValue_0_414_1 - _zz_realValue_0_414);
    end else begin
      realValue_0_414 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_414 = (_zz_when_ArraySlice_l166_414 <= _zz_when_ArraySlice_l166_414_2);
  assign when_ArraySlice_l158_415 = (_zz_when_ArraySlice_l158_415 <= _zz_when_ArraySlice_l158_415_3);
  assign when_ArraySlice_l159_415 = (_zz_when_ArraySlice_l159_415 <= _zz_when_ArraySlice_l159_415_2);
  assign _zz_realValue_0_415 = (_zz__zz_realValue_0_415 % _zz__zz_realValue_0_415_1);
  assign when_ArraySlice_l110_415 = (_zz_realValue_0_415 != 8'h0);
  always @(*) begin
    if(when_ArraySlice_l110_415) begin
      realValue_0_415 = (_zz_realValue_0_415_1 - _zz_realValue_0_415);
    end else begin
      realValue_0_415 = {1'd0, wReg};
    end
  end

  assign when_ArraySlice_l166_415 = (_zz_when_ArraySlice_l166_415 <= _zz_when_ArraySlice_l166_415_2);
  assign when_ArraySlice_l182_8 = (_zz_when_ArraySlice_l182_8 == _zz_when_ArraySlice_l182_8_1);
  assign when_ArraySlice_l183_8 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l182_8) begin
      if(when_ArraySlice_l183_8) begin
        _zz_when_ArraySlice_l357 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_9 = (_zz_when_ArraySlice_l182_9 == _zz_when_ArraySlice_l182_9_1);
  assign when_ArraySlice_l183_9 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l182_9) begin
      if(when_ArraySlice_l183_9) begin
        _zz_when_ArraySlice_l357_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_10 = (_zz_when_ArraySlice_l182_10 == _zz_when_ArraySlice_l182_10_1);
  assign when_ArraySlice_l183_10 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l182_10) begin
      if(when_ArraySlice_l183_10) begin
        _zz_when_ArraySlice_l357_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_11 = (_zz_when_ArraySlice_l182_11 == _zz_when_ArraySlice_l182_11_1);
  assign when_ArraySlice_l183_11 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l182_11) begin
      if(when_ArraySlice_l183_11) begin
        _zz_when_ArraySlice_l357_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_12 = (_zz_when_ArraySlice_l182_12 == _zz_when_ArraySlice_l182_12_1);
  assign when_ArraySlice_l183_12 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l182_12) begin
      if(when_ArraySlice_l183_12) begin
        _zz_when_ArraySlice_l357_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_13 = (_zz_when_ArraySlice_l182_13 == _zz_when_ArraySlice_l182_13_1);
  assign when_ArraySlice_l183_13 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l182_13) begin
      if(when_ArraySlice_l183_13) begin
        _zz_when_ArraySlice_l357_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_14 = (_zz_when_ArraySlice_l182_14 == _zz_when_ArraySlice_l182_14_1);
  assign when_ArraySlice_l183_14 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l182_14) begin
      if(when_ArraySlice_l183_14) begin
        _zz_when_ArraySlice_l357_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_15 = (_zz_when_ArraySlice_l182_15 == _zz_when_ArraySlice_l182_15_1);
  assign when_ArraySlice_l183_15 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l182_15) begin
      if(when_ArraySlice_l183_15) begin
        _zz_when_ArraySlice_l357_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l357_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l357_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l357 = (((((_zz_when_ArraySlice_l357_8 && _zz_when_ArraySlice_l357_12) && (holdReadOp_6 == _zz_when_ArraySlice_l357_13)) && (holdReadOp_7 == 1'b1)) && (! ((_zz_when_ArraySlice_l357_14 && _zz_when_ArraySlice_l357_18) && (debug_7_51 == _zz_when_ArraySlice_l357_19)))) && (! (((_zz_when_ArraySlice_l357_20 || _zz_when_ArraySlice_l357_24) || (_zz_when_ArraySlice_l357_6 != _zz_when_ArraySlice_l357_25)) || (_zz_when_ArraySlice_l357_7 != 1'b0))));
  assign when_ArraySlice_l182_16 = (_zz_when_ArraySlice_l182_16 == _zz_when_ArraySlice_l182_16_1);
  assign when_ArraySlice_l183_16 = (writeAround ^ readAround_0);
  always @(*) begin
    if(when_ArraySlice_l182_16) begin
      if(when_ArraySlice_l183_16) begin
        _zz_when_ArraySlice_l361 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_17 = (_zz_when_ArraySlice_l182_17 == _zz_when_ArraySlice_l182_17_1);
  assign when_ArraySlice_l183_17 = (writeAround ^ readAround_1);
  always @(*) begin
    if(when_ArraySlice_l182_17) begin
      if(when_ArraySlice_l183_17) begin
        _zz_when_ArraySlice_l361_1 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_1 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_1 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_18 = (_zz_when_ArraySlice_l182_18 == _zz_when_ArraySlice_l182_18_1);
  assign when_ArraySlice_l183_18 = (writeAround ^ readAround_2);
  always @(*) begin
    if(when_ArraySlice_l182_18) begin
      if(when_ArraySlice_l183_18) begin
        _zz_when_ArraySlice_l361_2 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_2 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_2 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_19 = (_zz_when_ArraySlice_l182_19 == _zz_when_ArraySlice_l182_19_1);
  assign when_ArraySlice_l183_19 = (writeAround ^ readAround_3);
  always @(*) begin
    if(when_ArraySlice_l182_19) begin
      if(when_ArraySlice_l183_19) begin
        _zz_when_ArraySlice_l361_3 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_3 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_3 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_20 = (_zz_when_ArraySlice_l182_20 == _zz_when_ArraySlice_l182_20_1);
  assign when_ArraySlice_l183_20 = (writeAround ^ readAround_4);
  always @(*) begin
    if(when_ArraySlice_l182_20) begin
      if(when_ArraySlice_l183_20) begin
        _zz_when_ArraySlice_l361_4 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_4 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_4 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_21 = (_zz_when_ArraySlice_l182_21 == _zz_when_ArraySlice_l182_21_1);
  assign when_ArraySlice_l183_21 = (writeAround ^ readAround_5);
  always @(*) begin
    if(when_ArraySlice_l182_21) begin
      if(when_ArraySlice_l183_21) begin
        _zz_when_ArraySlice_l361_5 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_5 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_5 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_22 = (_zz_when_ArraySlice_l182_22 == _zz_when_ArraySlice_l182_22_1);
  assign when_ArraySlice_l183_22 = (writeAround ^ readAround_6);
  always @(*) begin
    if(when_ArraySlice_l182_22) begin
      if(when_ArraySlice_l183_22) begin
        _zz_when_ArraySlice_l361_6 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_6 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_6 = 1'b0;
    end
  end

  assign when_ArraySlice_l182_23 = (_zz_when_ArraySlice_l182_23 == _zz_when_ArraySlice_l182_23_1);
  assign when_ArraySlice_l183_23 = (writeAround ^ readAround_7);
  always @(*) begin
    if(when_ArraySlice_l182_23) begin
      if(when_ArraySlice_l183_23) begin
        _zz_when_ArraySlice_l361_7 = 1'b1;
      end else begin
        _zz_when_ArraySlice_l361_7 = 1'b0;
      end
    end else begin
      _zz_when_ArraySlice_l361_7 = 1'b0;
    end
  end

  assign when_ArraySlice_l361 = ((((((((_zz_when_ArraySlice_l361 != 1'b0) || (_zz_when_ArraySlice_l361_1 != 1'b0)) || (_zz_when_ArraySlice_l361_2 != 1'b0)) || (_zz_when_ArraySlice_l361_3 != 1'b0)) || (_zz_when_ArraySlice_l361_4 != 1'b0)) || (_zz_when_ArraySlice_l361_5 != 1'b0)) || (_zz_when_ArraySlice_l361_6 != 1'b0)) || (_zz_when_ArraySlice_l361_7 != 1'b0));
  assign when_ArraySlice_l364 = (! allowPadding_0);
  assign when_ArraySlice_l364_1 = (! allowPadding_1);
  assign when_ArraySlice_l364_2 = (! allowPadding_2);
  assign when_ArraySlice_l364_3 = (! allowPadding_3);
  assign when_ArraySlice_l364_4 = (! allowPadding_4);
  assign when_ArraySlice_l364_5 = (! allowPadding_5);
  assign when_ArraySlice_l364_6 = (! allowPadding_6);
  assign when_ArraySlice_l364_7 = (! allowPadding_7);
  assign stateIndicate = arraySliceStateMachine_stateReg;
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      wReg <= 7'h7f;
      hReg <= 7'h7f;
      aReg <= 4'b1111;
      bReg <= 4'b1111;
      handshakeTimes_0_value <= 13'h0;
      handshakeTimes_1_value <= 13'h0;
      handshakeTimes_2_value <= 13'h0;
      handshakeTimes_3_value <= 13'h0;
      handshakeTimes_4_value <= 13'h0;
      handshakeTimes_5_value <= 13'h0;
      handshakeTimes_6_value <= 13'h0;
      handshakeTimes_7_value <= 13'h0;
      selectWriteFifo <= 7'h0;
      selectReadFifo_0 <= 8'h0;
      selectReadFifo_1 <= 8'h0;
      selectReadFifo_2 <= 8'h0;
      selectReadFifo_3 <= 8'h0;
      selectReadFifo_4 <= 8'h0;
      selectReadFifo_5 <= 8'h0;
      selectReadFifo_6 <= 8'h0;
      selectReadFifo_7 <= 8'h0;
      holdReadOp_0 <= 1'b0;
      holdReadOp_1 <= 1'b0;
      holdReadOp_2 <= 1'b0;
      holdReadOp_3 <= 1'b0;
      holdReadOp_4 <= 1'b0;
      holdReadOp_5 <= 1'b0;
      holdReadOp_6 <= 1'b0;
      holdReadOp_7 <= 1'b0;
      allowPadding_0 <= 1'b1;
      allowPadding_1 <= 1'b1;
      allowPadding_2 <= 1'b1;
      allowPadding_3 <= 1'b1;
      allowPadding_4 <= 1'b1;
      allowPadding_5 <= 1'b1;
      allowPadding_6 <= 1'b1;
      allowPadding_7 <= 1'b1;
      outSliceNumb_0_value <= 7'h0;
      outSliceNumb_1_value <= 7'h0;
      outSliceNumb_2_value <= 7'h0;
      outSliceNumb_3_value <= 7'h0;
      outSliceNumb_4_value <= 7'h0;
      outSliceNumb_5_value <= 7'h0;
      outSliceNumb_6_value <= 7'h0;
      outSliceNumb_7_value <= 7'h0;
      writeAround <= 1'b0;
      readAround_0 <= 1'b0;
      readAround_1 <= 1'b0;
      readAround_2 <= 1'b0;
      readAround_3 <= 1'b0;
      readAround_4 <= 1'b0;
      readAround_5 <= 1'b0;
      readAround_6 <= 1'b0;
      readAround_7 <= 1'b0;
      arraySliceStateMachine_stateReg <= arraySliceStateMachine_enumDef_BOOT;
    end else begin
      wReg <= inputFeatureMapWidth;
      hReg <= inputFeatureMapHeight;
      aReg <= outputFeatureMapHeight;
      bReg <= outputFeatureMapWidth;
      handshakeTimes_0_value <= handshakeTimes_0_valueNext;
      handshakeTimes_1_value <= handshakeTimes_1_valueNext;
      handshakeTimes_2_value <= handshakeTimes_2_valueNext;
      handshakeTimes_3_value <= handshakeTimes_3_valueNext;
      handshakeTimes_4_value <= handshakeTimes_4_valueNext;
      handshakeTimes_5_value <= handshakeTimes_5_valueNext;
      handshakeTimes_6_value <= handshakeTimes_6_valueNext;
      handshakeTimes_7_value <= handshakeTimes_7_valueNext;
      outSliceNumb_0_value <= outSliceNumb_0_valueNext;
      outSliceNumb_1_value <= outSliceNumb_1_valueNext;
      outSliceNumb_2_value <= outSliceNumb_2_valueNext;
      outSliceNumb_3_value <= outSliceNumb_3_valueNext;
      outSliceNumb_4_value <= outSliceNumb_4_valueNext;
      outSliceNumb_5_value <= outSliceNumb_5_valueNext;
      outSliceNumb_6_value <= outSliceNumb_6_valueNext;
      outSliceNumb_7_value <= outSliceNumb_7_valueNext;
      arraySliceStateMachine_stateReg <= arraySliceStateMachine_stateNext;
      case(arraySliceStateMachine_stateReg)
        arraySliceStateMachine_enumDef_writeDataOnly : begin
          if(when_ArraySlice_l208) begin
            if(when_ArraySlice_l209) begin
              selectWriteFifo <= 7'h0;
              writeAround <= (! writeAround);
            end else begin
              selectWriteFifo <= (selectWriteFifo + 7'h01);
            end
          end
          if(when_ArraySlice_l216) begin
            if(holdReadOp_0) begin
              holdReadOp_0 <= 1'b0;
            end
            if(when_ArraySlice_l222) begin
              allowPadding_0 <= 1'b1;
            end
            if(holdReadOp_1) begin
              holdReadOp_1 <= 1'b0;
            end
            if(when_ArraySlice_l222_1) begin
              allowPadding_1 <= 1'b1;
            end
            if(holdReadOp_2) begin
              holdReadOp_2 <= 1'b0;
            end
            if(when_ArraySlice_l222_2) begin
              allowPadding_2 <= 1'b1;
            end
            if(holdReadOp_3) begin
              holdReadOp_3 <= 1'b0;
            end
            if(when_ArraySlice_l222_3) begin
              allowPadding_3 <= 1'b1;
            end
            if(holdReadOp_4) begin
              holdReadOp_4 <= 1'b0;
            end
            if(when_ArraySlice_l222_4) begin
              allowPadding_4 <= 1'b1;
            end
            if(holdReadOp_5) begin
              holdReadOp_5 <= 1'b0;
            end
            if(when_ArraySlice_l222_5) begin
              allowPadding_5 <= 1'b1;
            end
            if(holdReadOp_6) begin
              holdReadOp_6 <= 1'b0;
            end
            if(when_ArraySlice_l222_6) begin
              allowPadding_6 <= 1'b1;
            end
            if(holdReadOp_7) begin
              holdReadOp_7 <= 1'b0;
            end
            if(when_ArraySlice_l222_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        arraySliceStateMachine_enumDef_readDataOnly : begin
          if(when_ArraySlice_l376) begin
            if(when_ArraySlice_l382) begin
              if(when_ArraySlice_l383) begin
                if(when_ArraySlice_l384) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392) begin
                if(when_ArraySlice_l393) begin
                  if(when_ArraySlice_l395) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_2 + _zz_selectReadFifo_0_4);
                  end else begin
                    if(when_ArraySlice_l400) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l403) begin
                      allowPadding_0 <= 1'b0;
                    end
                    if(when_ArraySlice_l406) begin
                      selectReadFifo_0 <= 8'h0;
                      readAround_0 <= (! readAround_0);
                    end else begin
                      selectReadFifo_0 <= (_zz_selectReadFifo_0_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417) begin
                if(when_ArraySlice_l418) begin
                  if(when_ArraySlice_l420) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l428) begin
                      allowPadding_0 <= 1'b0;
                    end
                    if(when_ArraySlice_l431) begin
                      selectReadFifo_0 <= 8'h0;
                      readAround_0 <= (! readAround_0);
                    end else begin
                      selectReadFifo_0 <= (_zz_selectReadFifo_0_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447) begin
              if(when_ArraySlice_l449) begin
                if(when_ArraySlice_l450) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_14 + 8'h01);
                end else begin
                  selectReadFifo_0 <= 8'h0;
                  readAround_0 <= (! readAround_0);
                  if(when_ArraySlice_l457) begin
                    holdReadOp_0 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461) begin
                  selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_1) begin
            if(when_ArraySlice_l382_1) begin
              if(when_ArraySlice_l383_1) begin
                if(when_ArraySlice_l384_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_1) begin
                if(when_ArraySlice_l393_1) begin
                  if(when_ArraySlice_l395_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_2 + _zz_selectReadFifo_1_4);
                  end else begin
                    if(when_ArraySlice_l400_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_1) begin
                      selectReadFifo_1 <= 8'h0;
                      readAround_1 <= (! readAround_1);
                    end else begin
                      selectReadFifo_1 <= (_zz_selectReadFifo_1_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_1) begin
                if(when_ArraySlice_l418_1) begin
                  if(when_ArraySlice_l420_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_1) begin
                      selectReadFifo_1 <= 8'h0;
                      readAround_1 <= (! readAround_1);
                    end else begin
                      selectReadFifo_1 <= (_zz_selectReadFifo_1_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_1) begin
              if(when_ArraySlice_l449_1) begin
                if(when_ArraySlice_l450_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_14 + 8'h01);
                end else begin
                  selectReadFifo_1 <= 8'h0;
                  readAround_1 <= (! readAround_1);
                  if(when_ArraySlice_l457_1) begin
                    holdReadOp_1 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_1) begin
                  selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_2) begin
            if(when_ArraySlice_l382_2) begin
              if(when_ArraySlice_l383_2) begin
                if(when_ArraySlice_l384_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_2) begin
                if(when_ArraySlice_l393_2) begin
                  if(when_ArraySlice_l395_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_2 + _zz_selectReadFifo_2_4);
                  end else begin
                    if(when_ArraySlice_l400_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_2) begin
                      selectReadFifo_2 <= 8'h0;
                      readAround_2 <= (! readAround_2);
                    end else begin
                      selectReadFifo_2 <= (_zz_selectReadFifo_2_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_2) begin
                if(when_ArraySlice_l418_2) begin
                  if(when_ArraySlice_l420_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_2) begin
                      selectReadFifo_2 <= 8'h0;
                      readAround_2 <= (! readAround_2);
                    end else begin
                      selectReadFifo_2 <= (_zz_selectReadFifo_2_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_2) begin
              if(when_ArraySlice_l449_2) begin
                if(when_ArraySlice_l450_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_14 + 8'h01);
                end else begin
                  selectReadFifo_2 <= 8'h0;
                  readAround_2 <= (! readAround_2);
                  if(when_ArraySlice_l457_2) begin
                    holdReadOp_2 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_2) begin
                  selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_3) begin
            if(when_ArraySlice_l382_3) begin
              if(when_ArraySlice_l383_3) begin
                if(when_ArraySlice_l384_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_3) begin
                if(when_ArraySlice_l393_3) begin
                  if(when_ArraySlice_l395_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_2 + _zz_selectReadFifo_3_4);
                  end else begin
                    if(when_ArraySlice_l400_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_3) begin
                      selectReadFifo_3 <= 8'h0;
                      readAround_3 <= (! readAround_3);
                    end else begin
                      selectReadFifo_3 <= (_zz_selectReadFifo_3_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_3) begin
                if(when_ArraySlice_l418_3) begin
                  if(when_ArraySlice_l420_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_3) begin
                      selectReadFifo_3 <= 8'h0;
                      readAround_3 <= (! readAround_3);
                    end else begin
                      selectReadFifo_3 <= (_zz_selectReadFifo_3_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_3) begin
              if(when_ArraySlice_l449_3) begin
                if(when_ArraySlice_l450_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_14 + 8'h01);
                end else begin
                  selectReadFifo_3 <= 8'h0;
                  readAround_3 <= (! readAround_3);
                  if(when_ArraySlice_l457_3) begin
                    holdReadOp_3 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_3) begin
                  selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_4) begin
            if(when_ArraySlice_l382_4) begin
              if(when_ArraySlice_l383_4) begin
                if(when_ArraySlice_l384_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_4) begin
                if(when_ArraySlice_l393_4) begin
                  if(when_ArraySlice_l395_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_2 + _zz_selectReadFifo_4_4);
                  end else begin
                    if(when_ArraySlice_l400_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_4) begin
                      selectReadFifo_4 <= 8'h0;
                      readAround_4 <= (! readAround_4);
                    end else begin
                      selectReadFifo_4 <= (_zz_selectReadFifo_4_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_4) begin
                if(when_ArraySlice_l418_4) begin
                  if(when_ArraySlice_l420_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_4) begin
                      selectReadFifo_4 <= 8'h0;
                      readAround_4 <= (! readAround_4);
                    end else begin
                      selectReadFifo_4 <= (_zz_selectReadFifo_4_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_4) begin
              if(when_ArraySlice_l449_4) begin
                if(when_ArraySlice_l450_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_14 + 8'h01);
                end else begin
                  selectReadFifo_4 <= 8'h0;
                  readAround_4 <= (! readAround_4);
                  if(when_ArraySlice_l457_4) begin
                    holdReadOp_4 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_4) begin
                  selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_5) begin
            if(when_ArraySlice_l382_5) begin
              if(when_ArraySlice_l383_5) begin
                if(when_ArraySlice_l384_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_5) begin
                if(when_ArraySlice_l393_5) begin
                  if(when_ArraySlice_l395_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_2 + _zz_selectReadFifo_5_4);
                  end else begin
                    if(when_ArraySlice_l400_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_5) begin
                      selectReadFifo_5 <= 8'h0;
                      readAround_5 <= (! readAround_5);
                    end else begin
                      selectReadFifo_5 <= (_zz_selectReadFifo_5_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_5) begin
                if(when_ArraySlice_l418_5) begin
                  if(when_ArraySlice_l420_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_5) begin
                      selectReadFifo_5 <= 8'h0;
                      readAround_5 <= (! readAround_5);
                    end else begin
                      selectReadFifo_5 <= (_zz_selectReadFifo_5_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_5) begin
              if(when_ArraySlice_l449_5) begin
                if(when_ArraySlice_l450_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_14 + 8'h01);
                end else begin
                  selectReadFifo_5 <= 8'h0;
                  readAround_5 <= (! readAround_5);
                  if(when_ArraySlice_l457_5) begin
                    holdReadOp_5 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_5) begin
                  selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_6) begin
            if(when_ArraySlice_l382_6) begin
              if(when_ArraySlice_l383_6) begin
                if(when_ArraySlice_l384_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_6) begin
                if(when_ArraySlice_l393_6) begin
                  if(when_ArraySlice_l395_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_2 + _zz_selectReadFifo_6_4);
                  end else begin
                    if(when_ArraySlice_l400_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_6) begin
                      selectReadFifo_6 <= 8'h0;
                      readAround_6 <= (! readAround_6);
                    end else begin
                      selectReadFifo_6 <= (_zz_selectReadFifo_6_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_6) begin
                if(when_ArraySlice_l418_6) begin
                  if(when_ArraySlice_l420_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_6) begin
                      selectReadFifo_6 <= 8'h0;
                      readAround_6 <= (! readAround_6);
                    end else begin
                      selectReadFifo_6 <= (_zz_selectReadFifo_6_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_6) begin
              if(when_ArraySlice_l449_6) begin
                if(when_ArraySlice_l450_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_14 + 8'h01);
                end else begin
                  selectReadFifo_6 <= 8'h0;
                  readAround_6 <= (! readAround_6);
                  if(when_ArraySlice_l457_6) begin
                    holdReadOp_6 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_6) begin
                  selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l376_7) begin
            if(when_ArraySlice_l382_7) begin
              if(when_ArraySlice_l383_7) begin
                if(when_ArraySlice_l384_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7 + 8'h01);
                end else begin
                  if(when_ArraySlice_l387_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l392_7) begin
                if(when_ArraySlice_l393_7) begin
                  if(when_ArraySlice_l395_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_2 + _zz_selectReadFifo_7_4);
                  end else begin
                    if(when_ArraySlice_l400_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l403_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                    if(when_ArraySlice_l406_7) begin
                      selectReadFifo_7 <= 8'h0;
                      readAround_7 <= (! readAround_7);
                    end else begin
                      selectReadFifo_7 <= (_zz_selectReadFifo_7_6 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l413_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l417_7) begin
                if(when_ArraySlice_l418_7) begin
                  if(when_ArraySlice_l420_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_9 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l425_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l428_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                    if(when_ArraySlice_l431_7) begin
                      selectReadFifo_7 <= 8'h0;
                      readAround_7 <= (! readAround_7);
                    end else begin
                      selectReadFifo_7 <= (_zz_selectReadFifo_7_11 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l438_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l447_7) begin
              if(when_ArraySlice_l449_7) begin
                if(when_ArraySlice_l450_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_14 + 8'h01);
                end else begin
                  selectReadFifo_7 <= 8'h0;
                  readAround_7 <= (! readAround_7);
                  if(when_ArraySlice_l457_7) begin
                    holdReadOp_7 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l461_7) begin
                  selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l478) begin
            holdReadOp_0 <= 1'b0;
            if(when_ArraySlice_l481) begin
              allowPadding_0 <= 1'b1;
            end
            holdReadOp_1 <= 1'b0;
            if(when_ArraySlice_l481_1) begin
              allowPadding_1 <= 1'b1;
            end
            holdReadOp_2 <= 1'b0;
            if(when_ArraySlice_l481_2) begin
              allowPadding_2 <= 1'b1;
            end
            holdReadOp_3 <= 1'b0;
            if(when_ArraySlice_l481_3) begin
              allowPadding_3 <= 1'b1;
            end
            holdReadOp_4 <= 1'b0;
            if(when_ArraySlice_l481_4) begin
              allowPadding_4 <= 1'b1;
            end
            holdReadOp_5 <= 1'b0;
            if(when_ArraySlice_l481_5) begin
              allowPadding_5 <= 1'b1;
            end
            holdReadOp_6 <= 1'b0;
            if(when_ArraySlice_l481_6) begin
              allowPadding_6 <= 1'b1;
            end
            holdReadOp_7 <= 1'b0;
            if(when_ArraySlice_l481_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        arraySliceStateMachine_enumDef_readWriteData : begin
          if(when_ArraySlice_l233) begin
            if(when_ArraySlice_l239) begin
              if(when_ArraySlice_l240) begin
                if(when_ArraySlice_l241) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249) begin
                if(when_ArraySlice_l250) begin
                  if(when_ArraySlice_l252) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_18 + _zz_selectReadFifo_0_20);
                  end else begin
                    if(when_ArraySlice_l257) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l260) begin
                      allowPadding_0 <= 1'b0;
                    end
                    if(when_ArraySlice_l263) begin
                      selectReadFifo_0 <= 8'h0;
                      readAround_0 <= (! readAround_0);
                    end else begin
                      selectReadFifo_0 <= (_zz_selectReadFifo_0_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274) begin
                if(when_ArraySlice_l275) begin
                  if(when_ArraySlice_l277) begin
                    selectReadFifo_0 <= (_zz_selectReadFifo_0_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282) begin
                      holdReadOp_0 <= 1'b1;
                    end
                    if(when_ArraySlice_l285) begin
                      allowPadding_0 <= 1'b0;
                    end
                    if(when_ArraySlice_l288) begin
                      selectReadFifo_0 <= 8'h0;
                      readAround_0 <= (! readAround_0);
                    end else begin
                      selectReadFifo_0 <= (_zz_selectReadFifo_0_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295) begin
                    selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304) begin
              if(when_ArraySlice_l306) begin
                if(when_ArraySlice_l307) begin
                  selectReadFifo_0 <= (_zz_selectReadFifo_0_30 + 8'h01);
                end else begin
                  selectReadFifo_0 <= 8'h0;
                  readAround_0 <= (! readAround_0);
                  if(when_ArraySlice_l314) begin
                    holdReadOp_0 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318) begin
                  selectReadFifo_0 <= (selectReadFifo_0 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_1) begin
            if(when_ArraySlice_l239_1) begin
              if(when_ArraySlice_l240_1) begin
                if(when_ArraySlice_l241_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_1) begin
                if(when_ArraySlice_l250_1) begin
                  if(when_ArraySlice_l252_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_18 + _zz_selectReadFifo_1_20);
                  end else begin
                    if(when_ArraySlice_l257_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_1) begin
                      selectReadFifo_1 <= 8'h0;
                      readAround_1 <= (! readAround_1);
                    end else begin
                      selectReadFifo_1 <= (_zz_selectReadFifo_1_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_1) begin
                if(when_ArraySlice_l275_1) begin
                  if(when_ArraySlice_l277_1) begin
                    selectReadFifo_1 <= (_zz_selectReadFifo_1_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_1) begin
                      holdReadOp_1 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_1) begin
                      allowPadding_1 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_1) begin
                      selectReadFifo_1 <= 8'h0;
                      readAround_1 <= (! readAround_1);
                    end else begin
                      selectReadFifo_1 <= (_zz_selectReadFifo_1_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_1) begin
                    selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_1) begin
              if(when_ArraySlice_l306_1) begin
                if(when_ArraySlice_l307_1) begin
                  selectReadFifo_1 <= (_zz_selectReadFifo_1_30 + 8'h01);
                end else begin
                  selectReadFifo_1 <= 8'h0;
                  readAround_1 <= (! readAround_1);
                  if(when_ArraySlice_l314_1) begin
                    holdReadOp_1 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_1) begin
                  selectReadFifo_1 <= (selectReadFifo_1 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_2) begin
            if(when_ArraySlice_l239_2) begin
              if(when_ArraySlice_l240_2) begin
                if(when_ArraySlice_l241_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_2) begin
                if(when_ArraySlice_l250_2) begin
                  if(when_ArraySlice_l252_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_18 + _zz_selectReadFifo_2_20);
                  end else begin
                    if(when_ArraySlice_l257_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_2) begin
                      selectReadFifo_2 <= 8'h0;
                      readAround_2 <= (! readAround_2);
                    end else begin
                      selectReadFifo_2 <= (_zz_selectReadFifo_2_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_2) begin
                if(when_ArraySlice_l275_2) begin
                  if(when_ArraySlice_l277_2) begin
                    selectReadFifo_2 <= (_zz_selectReadFifo_2_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_2) begin
                      holdReadOp_2 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_2) begin
                      allowPadding_2 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_2) begin
                      selectReadFifo_2 <= 8'h0;
                      readAround_2 <= (! readAround_2);
                    end else begin
                      selectReadFifo_2 <= (_zz_selectReadFifo_2_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_2) begin
                    selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_2) begin
              if(when_ArraySlice_l306_2) begin
                if(when_ArraySlice_l307_2) begin
                  selectReadFifo_2 <= (_zz_selectReadFifo_2_30 + 8'h01);
                end else begin
                  selectReadFifo_2 <= 8'h0;
                  readAround_2 <= (! readAround_2);
                  if(when_ArraySlice_l314_2) begin
                    holdReadOp_2 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_2) begin
                  selectReadFifo_2 <= (selectReadFifo_2 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_3) begin
            if(when_ArraySlice_l239_3) begin
              if(when_ArraySlice_l240_3) begin
                if(when_ArraySlice_l241_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_3) begin
                if(when_ArraySlice_l250_3) begin
                  if(when_ArraySlice_l252_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_18 + _zz_selectReadFifo_3_20);
                  end else begin
                    if(when_ArraySlice_l257_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_3) begin
                      selectReadFifo_3 <= 8'h0;
                      readAround_3 <= (! readAround_3);
                    end else begin
                      selectReadFifo_3 <= (_zz_selectReadFifo_3_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_3) begin
                if(when_ArraySlice_l275_3) begin
                  if(when_ArraySlice_l277_3) begin
                    selectReadFifo_3 <= (_zz_selectReadFifo_3_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_3) begin
                      holdReadOp_3 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_3) begin
                      allowPadding_3 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_3) begin
                      selectReadFifo_3 <= 8'h0;
                      readAround_3 <= (! readAround_3);
                    end else begin
                      selectReadFifo_3 <= (_zz_selectReadFifo_3_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_3) begin
                    selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_3) begin
              if(when_ArraySlice_l306_3) begin
                if(when_ArraySlice_l307_3) begin
                  selectReadFifo_3 <= (_zz_selectReadFifo_3_30 + 8'h01);
                end else begin
                  selectReadFifo_3 <= 8'h0;
                  readAround_3 <= (! readAround_3);
                  if(when_ArraySlice_l314_3) begin
                    holdReadOp_3 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_3) begin
                  selectReadFifo_3 <= (selectReadFifo_3 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_4) begin
            if(when_ArraySlice_l239_4) begin
              if(when_ArraySlice_l240_4) begin
                if(when_ArraySlice_l241_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_4) begin
                if(when_ArraySlice_l250_4) begin
                  if(when_ArraySlice_l252_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_18 + _zz_selectReadFifo_4_20);
                  end else begin
                    if(when_ArraySlice_l257_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_4) begin
                      selectReadFifo_4 <= 8'h0;
                      readAround_4 <= (! readAround_4);
                    end else begin
                      selectReadFifo_4 <= (_zz_selectReadFifo_4_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_4) begin
                if(when_ArraySlice_l275_4) begin
                  if(when_ArraySlice_l277_4) begin
                    selectReadFifo_4 <= (_zz_selectReadFifo_4_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_4) begin
                      holdReadOp_4 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_4) begin
                      allowPadding_4 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_4) begin
                      selectReadFifo_4 <= 8'h0;
                      readAround_4 <= (! readAround_4);
                    end else begin
                      selectReadFifo_4 <= (_zz_selectReadFifo_4_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_4) begin
                    selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_4) begin
              if(when_ArraySlice_l306_4) begin
                if(when_ArraySlice_l307_4) begin
                  selectReadFifo_4 <= (_zz_selectReadFifo_4_30 + 8'h01);
                end else begin
                  selectReadFifo_4 <= 8'h0;
                  readAround_4 <= (! readAround_4);
                  if(when_ArraySlice_l314_4) begin
                    holdReadOp_4 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_4) begin
                  selectReadFifo_4 <= (selectReadFifo_4 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_5) begin
            if(when_ArraySlice_l239_5) begin
              if(when_ArraySlice_l240_5) begin
                if(when_ArraySlice_l241_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_5) begin
                if(when_ArraySlice_l250_5) begin
                  if(when_ArraySlice_l252_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_18 + _zz_selectReadFifo_5_20);
                  end else begin
                    if(when_ArraySlice_l257_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_5) begin
                      selectReadFifo_5 <= 8'h0;
                      readAround_5 <= (! readAround_5);
                    end else begin
                      selectReadFifo_5 <= (_zz_selectReadFifo_5_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_5) begin
                if(when_ArraySlice_l275_5) begin
                  if(when_ArraySlice_l277_5) begin
                    selectReadFifo_5 <= (_zz_selectReadFifo_5_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_5) begin
                      holdReadOp_5 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_5) begin
                      allowPadding_5 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_5) begin
                      selectReadFifo_5 <= 8'h0;
                      readAround_5 <= (! readAround_5);
                    end else begin
                      selectReadFifo_5 <= (_zz_selectReadFifo_5_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_5) begin
                    selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_5) begin
              if(when_ArraySlice_l306_5) begin
                if(when_ArraySlice_l307_5) begin
                  selectReadFifo_5 <= (_zz_selectReadFifo_5_30 + 8'h01);
                end else begin
                  selectReadFifo_5 <= 8'h0;
                  readAround_5 <= (! readAround_5);
                  if(when_ArraySlice_l314_5) begin
                    holdReadOp_5 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_5) begin
                  selectReadFifo_5 <= (selectReadFifo_5 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_6) begin
            if(when_ArraySlice_l239_6) begin
              if(when_ArraySlice_l240_6) begin
                if(when_ArraySlice_l241_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_6) begin
                if(when_ArraySlice_l250_6) begin
                  if(when_ArraySlice_l252_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_18 + _zz_selectReadFifo_6_20);
                  end else begin
                    if(when_ArraySlice_l257_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_6) begin
                      selectReadFifo_6 <= 8'h0;
                      readAround_6 <= (! readAround_6);
                    end else begin
                      selectReadFifo_6 <= (_zz_selectReadFifo_6_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_6) begin
                if(when_ArraySlice_l275_6) begin
                  if(when_ArraySlice_l277_6) begin
                    selectReadFifo_6 <= (_zz_selectReadFifo_6_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_6) begin
                      holdReadOp_6 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_6) begin
                      allowPadding_6 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_6) begin
                      selectReadFifo_6 <= 8'h0;
                      readAround_6 <= (! readAround_6);
                    end else begin
                      selectReadFifo_6 <= (_zz_selectReadFifo_6_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_6) begin
                    selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_6) begin
              if(when_ArraySlice_l306_6) begin
                if(when_ArraySlice_l307_6) begin
                  selectReadFifo_6 <= (_zz_selectReadFifo_6_30 + 8'h01);
                end else begin
                  selectReadFifo_6 <= 8'h0;
                  readAround_6 <= (! readAround_6);
                  if(when_ArraySlice_l314_6) begin
                    holdReadOp_6 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_6) begin
                  selectReadFifo_6 <= (selectReadFifo_6 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l233_7) begin
            if(when_ArraySlice_l239_7) begin
              if(when_ArraySlice_l240_7) begin
                if(when_ArraySlice_l241_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_16 + 8'h01);
                end else begin
                  if(when_ArraySlice_l244_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l249_7) begin
                if(when_ArraySlice_l250_7) begin
                  if(when_ArraySlice_l252_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_18 + _zz_selectReadFifo_7_20);
                  end else begin
                    if(when_ArraySlice_l257_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l260_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                    if(when_ArraySlice_l263_7) begin
                      selectReadFifo_7 <= 8'h0;
                      readAround_7 <= (! readAround_7);
                    end else begin
                      selectReadFifo_7 <= (_zz_selectReadFifo_7_22 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l270_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
              if(when_ArraySlice_l274_7) begin
                if(when_ArraySlice_l275_7) begin
                  if(when_ArraySlice_l277_7) begin
                    selectReadFifo_7 <= (_zz_selectReadFifo_7_25 + 8'h01);
                  end else begin
                    if(when_ArraySlice_l282_7) begin
                      holdReadOp_7 <= 1'b1;
                    end
                    if(when_ArraySlice_l285_7) begin
                      allowPadding_7 <= 1'b0;
                    end
                    if(when_ArraySlice_l288_7) begin
                      selectReadFifo_7 <= 8'h0;
                      readAround_7 <= (! readAround_7);
                    end else begin
                      selectReadFifo_7 <= (_zz_selectReadFifo_7_27 + 8'h01);
                    end
                  end
                end else begin
                  if(when_ArraySlice_l295_7) begin
                    selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                  end
                end
              end
            end
          end else begin
            if(when_ArraySlice_l304_7) begin
              if(when_ArraySlice_l306_7) begin
                if(when_ArraySlice_l307_7) begin
                  selectReadFifo_7 <= (_zz_selectReadFifo_7_30 + 8'h01);
                end else begin
                  selectReadFifo_7 <= 8'h0;
                  readAround_7 <= (! readAround_7);
                  if(when_ArraySlice_l314_7) begin
                    holdReadOp_7 <= 1'b1;
                  end
                end
              end else begin
                if(when_ArraySlice_l318_7) begin
                  selectReadFifo_7 <= (selectReadFifo_7 + 8'h01);
                end
              end
            end
          end
          if(when_ArraySlice_l336) begin
            if(when_ArraySlice_l341) begin
              if(when_ArraySlice_l342) begin
                selectWriteFifo <= 7'h0;
                writeAround <= (! writeAround);
              end else begin
                selectWriteFifo <= (selectWriteFifo + 7'h01);
              end
            end
          end
          if(when_ArraySlice_l353) begin
            holdReadOp_0 <= 1'b0;
            holdReadOp_1 <= 1'b0;
            holdReadOp_2 <= 1'b0;
            holdReadOp_3 <= 1'b0;
            holdReadOp_4 <= 1'b0;
            holdReadOp_5 <= 1'b0;
            holdReadOp_6 <= 1'b0;
            holdReadOp_7 <= 1'b0;
          end
          if(when_ArraySlice_l361) begin
            if(when_ArraySlice_l364) begin
              allowPadding_0 <= 1'b1;
            end
            if(when_ArraySlice_l364_1) begin
              allowPadding_1 <= 1'b1;
            end
            if(when_ArraySlice_l364_2) begin
              allowPadding_2 <= 1'b1;
            end
            if(when_ArraySlice_l364_3) begin
              allowPadding_3 <= 1'b1;
            end
            if(when_ArraySlice_l364_4) begin
              allowPadding_4 <= 1'b1;
            end
            if(when_ArraySlice_l364_5) begin
              allowPadding_5 <= 1'b1;
            end
            if(when_ArraySlice_l364_6) begin
              allowPadding_6 <= 1'b1;
            end
            if(when_ArraySlice_l364_7) begin
              allowPadding_7 <= 1'b1;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end


endmodule

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

//StreamFifo replaced by StreamFifo

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [31:0]   io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [31:0]   io_pop_payload,
  input               io_flush,
  output reg [6:0]    io_occupancy,
  output reg [6:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [31:0]   _zz_logic_ram_port0;
  wire       [6:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [6:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [6:0]    _zz_io_occupancy;
  wire       [6:0]    _zz_io_availability;
  wire       [6:0]    _zz_io_availability_1;
  wire       [6:0]    _zz_io_availability_2;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [6:0]    logic_pushPtr_valueNext;
  reg        [6:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [6:0]    logic_popPtr_valueNext;
  reg        [6:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1021;
  wire       [6:0]    logic_ptrDif;
  reg [31:0] logic_ram [0:64];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {6'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {6'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_occupancy = (7'h41 + logic_ptrDif);
  assign _zz_io_availability = (7'h41 + _zz_io_availability_1);
  assign _zz_io_availability_1 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_availability_2 = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 7'h40);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    if(logic_pushPtr_willOverflow) begin
      logic_pushPtr_valueNext = 7'h0;
    end else begin
      logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    end
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 7'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 7'h40);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    if(logic_popPtr_willOverflow) begin
      logic_popPtr_valueNext = 7'h0;
    end else begin
      logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    end
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 7'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1021 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  always @(*) begin
    if(logic_ptrMatch) begin
      io_occupancy = (logic_risingOccupancy ? 7'h41 : 7'h0);
    end else begin
      io_occupancy = ((logic_popPtr_value < logic_pushPtr_value) ? logic_ptrDif : _zz_io_occupancy);
    end
  end

  always @(*) begin
    if(logic_ptrMatch) begin
      io_availability = (logic_risingOccupancy ? 7'h0 : 7'h41);
    end else begin
      io_availability = ((logic_popPtr_value < logic_pushPtr_value) ? _zz_io_availability : _zz_io_availability_2);
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      logic_pushPtr_value <= 7'h0;
      logic_popPtr_value <= 7'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1021) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule
