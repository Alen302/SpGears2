// Generator : SpinalHDL v1.6.1    git head : 3bf789d53b1b5a36974196e2d591342e15ddf28c
// Component : BitonicSortV2
// Git hash  : 8d6817b04a83e60e2277aeee5860ca026b136cda

`timescale 1ns/1ps 

module BitonicSortV2 (
  input               dataIn_valid,
  input      [7:0]    dataIn_payload_0,
  input      [7:0]    dataIn_payload_1,
  input      [7:0]    dataIn_payload_2,
  input      [7:0]    dataIn_payload_3,
  input      [7:0]    dataIn_payload_4,
  input      [7:0]    dataIn_payload_5,
  input      [7:0]    dataIn_payload_6,
  input      [7:0]    dataIn_payload_7,
  input      [7:0]    dataIn_payload_8,
  input      [7:0]    dataIn_payload_9,
  input      [7:0]    dataIn_payload_10,
  input      [7:0]    dataIn_payload_11,
  input      [7:0]    dataIn_payload_12,
  input      [7:0]    dataIn_payload_13,
  input      [7:0]    dataIn_payload_14,
  input      [7:0]    dataIn_payload_15,
  input      [7:0]    dataIn_payload_16,
  input      [7:0]    dataIn_payload_17,
  input      [7:0]    dataIn_payload_18,
  input      [7:0]    dataIn_payload_19,
  input      [7:0]    dataIn_payload_20,
  input      [7:0]    dataIn_payload_21,
  input      [7:0]    dataIn_payload_22,
  input      [7:0]    dataIn_payload_23,
  input      [7:0]    dataIn_payload_24,
  input      [7:0]    dataIn_payload_25,
  input      [7:0]    dataIn_payload_26,
  input      [7:0]    dataIn_payload_27,
  input      [7:0]    dataIn_payload_28,
  input      [7:0]    dataIn_payload_29,
  input      [7:0]    dataIn_payload_30,
  input      [7:0]    dataIn_payload_31,
  input      [7:0]    dataIn_payload_32,
  input      [7:0]    dataIn_payload_33,
  input      [7:0]    dataIn_payload_34,
  input      [7:0]    dataIn_payload_35,
  input      [7:0]    dataIn_payload_36,
  input      [7:0]    dataIn_payload_37,
  input      [7:0]    dataIn_payload_38,
  input      [7:0]    dataIn_payload_39,
  input      [7:0]    dataIn_payload_40,
  input      [7:0]    dataIn_payload_41,
  input      [7:0]    dataIn_payload_42,
  input      [7:0]    dataIn_payload_43,
  input      [7:0]    dataIn_payload_44,
  input      [7:0]    dataIn_payload_45,
  input      [7:0]    dataIn_payload_46,
  input      [7:0]    dataIn_payload_47,
  input      [7:0]    dataIn_payload_48,
  input      [7:0]    dataIn_payload_49,
  input      [7:0]    dataIn_payload_50,
  input      [7:0]    dataIn_payload_51,
  input      [7:0]    dataIn_payload_52,
  input      [7:0]    dataIn_payload_53,
  input      [7:0]    dataIn_payload_54,
  input      [7:0]    dataIn_payload_55,
  input      [7:0]    dataIn_payload_56,
  input      [7:0]    dataIn_payload_57,
  input      [7:0]    dataIn_payload_58,
  input      [7:0]    dataIn_payload_59,
  input      [7:0]    dataIn_payload_60,
  input      [7:0]    dataIn_payload_61,
  input      [7:0]    dataIn_payload_62,
  input      [7:0]    dataIn_payload_63,
  input      [7:0]    dataIn_payload_64,
  input      [7:0]    dataIn_payload_65,
  input      [7:0]    dataIn_payload_66,
  input      [7:0]    dataIn_payload_67,
  input      [7:0]    dataIn_payload_68,
  input      [7:0]    dataIn_payload_69,
  input      [7:0]    dataIn_payload_70,
  input      [7:0]    dataIn_payload_71,
  input      [7:0]    dataIn_payload_72,
  input      [7:0]    dataIn_payload_73,
  input      [7:0]    dataIn_payload_74,
  input      [7:0]    dataIn_payload_75,
  input      [7:0]    dataIn_payload_76,
  input      [7:0]    dataIn_payload_77,
  input      [7:0]    dataIn_payload_78,
  input      [7:0]    dataIn_payload_79,
  input      [7:0]    dataIn_payload_80,
  input      [7:0]    dataIn_payload_81,
  input      [7:0]    dataIn_payload_82,
  input      [7:0]    dataIn_payload_83,
  input      [7:0]    dataIn_payload_84,
  input      [7:0]    dataIn_payload_85,
  input      [7:0]    dataIn_payload_86,
  input      [7:0]    dataIn_payload_87,
  input      [7:0]    dataIn_payload_88,
  input      [7:0]    dataIn_payload_89,
  input      [7:0]    dataIn_payload_90,
  input      [7:0]    dataIn_payload_91,
  input      [7:0]    dataIn_payload_92,
  input      [7:0]    dataIn_payload_93,
  input      [7:0]    dataIn_payload_94,
  input      [7:0]    dataIn_payload_95,
  input      [7:0]    dataIn_payload_96,
  input      [7:0]    dataIn_payload_97,
  input      [7:0]    dataIn_payload_98,
  input      [7:0]    dataIn_payload_99,
  input      [7:0]    dataIn_payload_100,
  input      [7:0]    dataIn_payload_101,
  input      [7:0]    dataIn_payload_102,
  input      [7:0]    dataIn_payload_103,
  input      [7:0]    dataIn_payload_104,
  input      [7:0]    dataIn_payload_105,
  input      [7:0]    dataIn_payload_106,
  input      [7:0]    dataIn_payload_107,
  input      [7:0]    dataIn_payload_108,
  input      [7:0]    dataIn_payload_109,
  input      [7:0]    dataIn_payload_110,
  input      [7:0]    dataIn_payload_111,
  input      [7:0]    dataIn_payload_112,
  input      [7:0]    dataIn_payload_113,
  input      [7:0]    dataIn_payload_114,
  input      [7:0]    dataIn_payload_115,
  input      [7:0]    dataIn_payload_116,
  input      [7:0]    dataIn_payload_117,
  input      [7:0]    dataIn_payload_118,
  input      [7:0]    dataIn_payload_119,
  input      [7:0]    dataIn_payload_120,
  input      [7:0]    dataIn_payload_121,
  input      [7:0]    dataIn_payload_122,
  input      [7:0]    dataIn_payload_123,
  input      [7:0]    dataIn_payload_124,
  input      [7:0]    dataIn_payload_125,
  input      [7:0]    dataIn_payload_126,
  input      [7:0]    dataIn_payload_127,
  input      [7:0]    dataIn_payload_128,
  input      [7:0]    dataIn_payload_129,
  input      [7:0]    dataIn_payload_130,
  input      [7:0]    dataIn_payload_131,
  input      [7:0]    dataIn_payload_132,
  input      [7:0]    dataIn_payload_133,
  input      [7:0]    dataIn_payload_134,
  input      [7:0]    dataIn_payload_135,
  input      [7:0]    dataIn_payload_136,
  input      [7:0]    dataIn_payload_137,
  input      [7:0]    dataIn_payload_138,
  input      [7:0]    dataIn_payload_139,
  input      [7:0]    dataIn_payload_140,
  input      [7:0]    dataIn_payload_141,
  input      [7:0]    dataIn_payload_142,
  input      [7:0]    dataIn_payload_143,
  input      [7:0]    dataIn_payload_144,
  input      [7:0]    dataIn_payload_145,
  input      [7:0]    dataIn_payload_146,
  input      [7:0]    dataIn_payload_147,
  input      [7:0]    dataIn_payload_148,
  input      [7:0]    dataIn_payload_149,
  input      [7:0]    dataIn_payload_150,
  input      [7:0]    dataIn_payload_151,
  input      [7:0]    dataIn_payload_152,
  input      [7:0]    dataIn_payload_153,
  input      [7:0]    dataIn_payload_154,
  input      [7:0]    dataIn_payload_155,
  input      [7:0]    dataIn_payload_156,
  input      [7:0]    dataIn_payload_157,
  input      [7:0]    dataIn_payload_158,
  input      [7:0]    dataIn_payload_159,
  input      [7:0]    dataIn_payload_160,
  input      [7:0]    dataIn_payload_161,
  input      [7:0]    dataIn_payload_162,
  input      [7:0]    dataIn_payload_163,
  input      [7:0]    dataIn_payload_164,
  input      [7:0]    dataIn_payload_165,
  input      [7:0]    dataIn_payload_166,
  input      [7:0]    dataIn_payload_167,
  input      [7:0]    dataIn_payload_168,
  input      [7:0]    dataIn_payload_169,
  input      [7:0]    dataIn_payload_170,
  input      [7:0]    dataIn_payload_171,
  input      [7:0]    dataIn_payload_172,
  input      [7:0]    dataIn_payload_173,
  input      [7:0]    dataIn_payload_174,
  input      [7:0]    dataIn_payload_175,
  input      [7:0]    dataIn_payload_176,
  input      [7:0]    dataIn_payload_177,
  input      [7:0]    dataIn_payload_178,
  input      [7:0]    dataIn_payload_179,
  input      [7:0]    dataIn_payload_180,
  input      [7:0]    dataIn_payload_181,
  input      [7:0]    dataIn_payload_182,
  input      [7:0]    dataIn_payload_183,
  input      [7:0]    dataIn_payload_184,
  input      [7:0]    dataIn_payload_185,
  input      [7:0]    dataIn_payload_186,
  input      [7:0]    dataIn_payload_187,
  input      [7:0]    dataIn_payload_188,
  input      [7:0]    dataIn_payload_189,
  input      [7:0]    dataIn_payload_190,
  input      [7:0]    dataIn_payload_191,
  input      [7:0]    dataIn_payload_192,
  input      [7:0]    dataIn_payload_193,
  input      [7:0]    dataIn_payload_194,
  input      [7:0]    dataIn_payload_195,
  input      [7:0]    dataIn_payload_196,
  input      [7:0]    dataIn_payload_197,
  input      [7:0]    dataIn_payload_198,
  input      [7:0]    dataIn_payload_199,
  input      [7:0]    dataIn_payload_200,
  input      [7:0]    dataIn_payload_201,
  input      [7:0]    dataIn_payload_202,
  input      [7:0]    dataIn_payload_203,
  input      [7:0]    dataIn_payload_204,
  input      [7:0]    dataIn_payload_205,
  input      [7:0]    dataIn_payload_206,
  input      [7:0]    dataIn_payload_207,
  input      [7:0]    dataIn_payload_208,
  input      [7:0]    dataIn_payload_209,
  input      [7:0]    dataIn_payload_210,
  input      [7:0]    dataIn_payload_211,
  input      [7:0]    dataIn_payload_212,
  input      [7:0]    dataIn_payload_213,
  input      [7:0]    dataIn_payload_214,
  input      [7:0]    dataIn_payload_215,
  input      [7:0]    dataIn_payload_216,
  input      [7:0]    dataIn_payload_217,
  input      [7:0]    dataIn_payload_218,
  input      [7:0]    dataIn_payload_219,
  input      [7:0]    dataIn_payload_220,
  input      [7:0]    dataIn_payload_221,
  input      [7:0]    dataIn_payload_222,
  input      [7:0]    dataIn_payload_223,
  input      [7:0]    dataIn_payload_224,
  input      [7:0]    dataIn_payload_225,
  input      [7:0]    dataIn_payload_226,
  input      [7:0]    dataIn_payload_227,
  input      [7:0]    dataIn_payload_228,
  input      [7:0]    dataIn_payload_229,
  input      [7:0]    dataIn_payload_230,
  input      [7:0]    dataIn_payload_231,
  input      [7:0]    dataIn_payload_232,
  input      [7:0]    dataIn_payload_233,
  input      [7:0]    dataIn_payload_234,
  input      [7:0]    dataIn_payload_235,
  input      [7:0]    dataIn_payload_236,
  input      [7:0]    dataIn_payload_237,
  input      [7:0]    dataIn_payload_238,
  input      [7:0]    dataIn_payload_239,
  input      [7:0]    dataIn_payload_240,
  input      [7:0]    dataIn_payload_241,
  input      [7:0]    dataIn_payload_242,
  input      [7:0]    dataIn_payload_243,
  input      [7:0]    dataIn_payload_244,
  input      [7:0]    dataIn_payload_245,
  input      [7:0]    dataIn_payload_246,
  input      [7:0]    dataIn_payload_247,
  input      [7:0]    dataIn_payload_248,
  input      [7:0]    dataIn_payload_249,
  input      [7:0]    dataIn_payload_250,
  input      [7:0]    dataIn_payload_251,
  input      [7:0]    dataIn_payload_252,
  input      [7:0]    dataIn_payload_253,
  input      [7:0]    dataIn_payload_254,
  input      [7:0]    dataIn_payload_255,
  output              dataOut_valid,
  output     [7:0]    dataOut_payload_0,
  output     [7:0]    dataOut_payload_1,
  output     [7:0]    dataOut_payload_2,
  output     [7:0]    dataOut_payload_3,
  output     [7:0]    dataOut_payload_4,
  output     [7:0]    dataOut_payload_5,
  output     [7:0]    dataOut_payload_6,
  output     [7:0]    dataOut_payload_7,
  output     [7:0]    dataOut_payload_8,
  output     [7:0]    dataOut_payload_9,
  output     [7:0]    dataOut_payload_10,
  output     [7:0]    dataOut_payload_11,
  output     [7:0]    dataOut_payload_12,
  output     [7:0]    dataOut_payload_13,
  output     [7:0]    dataOut_payload_14,
  output     [7:0]    dataOut_payload_15,
  output     [7:0]    dataOut_payload_16,
  output     [7:0]    dataOut_payload_17,
  output     [7:0]    dataOut_payload_18,
  output     [7:0]    dataOut_payload_19,
  output     [7:0]    dataOut_payload_20,
  output     [7:0]    dataOut_payload_21,
  output     [7:0]    dataOut_payload_22,
  output     [7:0]    dataOut_payload_23,
  output     [7:0]    dataOut_payload_24,
  output     [7:0]    dataOut_payload_25,
  output     [7:0]    dataOut_payload_26,
  output     [7:0]    dataOut_payload_27,
  output     [7:0]    dataOut_payload_28,
  output     [7:0]    dataOut_payload_29,
  output     [7:0]    dataOut_payload_30,
  output     [7:0]    dataOut_payload_31,
  output     [7:0]    dataOut_payload_32,
  output     [7:0]    dataOut_payload_33,
  output     [7:0]    dataOut_payload_34,
  output     [7:0]    dataOut_payload_35,
  output     [7:0]    dataOut_payload_36,
  output     [7:0]    dataOut_payload_37,
  output     [7:0]    dataOut_payload_38,
  output     [7:0]    dataOut_payload_39,
  output     [7:0]    dataOut_payload_40,
  output     [7:0]    dataOut_payload_41,
  output     [7:0]    dataOut_payload_42,
  output     [7:0]    dataOut_payload_43,
  output     [7:0]    dataOut_payload_44,
  output     [7:0]    dataOut_payload_45,
  output     [7:0]    dataOut_payload_46,
  output     [7:0]    dataOut_payload_47,
  output     [7:0]    dataOut_payload_48,
  output     [7:0]    dataOut_payload_49,
  output     [7:0]    dataOut_payload_50,
  output     [7:0]    dataOut_payload_51,
  output     [7:0]    dataOut_payload_52,
  output     [7:0]    dataOut_payload_53,
  output     [7:0]    dataOut_payload_54,
  output     [7:0]    dataOut_payload_55,
  output     [7:0]    dataOut_payload_56,
  output     [7:0]    dataOut_payload_57,
  output     [7:0]    dataOut_payload_58,
  output     [7:0]    dataOut_payload_59,
  output     [7:0]    dataOut_payload_60,
  output     [7:0]    dataOut_payload_61,
  output     [7:0]    dataOut_payload_62,
  output     [7:0]    dataOut_payload_63,
  output     [7:0]    dataOut_payload_64,
  output     [7:0]    dataOut_payload_65,
  output     [7:0]    dataOut_payload_66,
  output     [7:0]    dataOut_payload_67,
  output     [7:0]    dataOut_payload_68,
  output     [7:0]    dataOut_payload_69,
  output     [7:0]    dataOut_payload_70,
  output     [7:0]    dataOut_payload_71,
  output     [7:0]    dataOut_payload_72,
  output     [7:0]    dataOut_payload_73,
  output     [7:0]    dataOut_payload_74,
  output     [7:0]    dataOut_payload_75,
  output     [7:0]    dataOut_payload_76,
  output     [7:0]    dataOut_payload_77,
  output     [7:0]    dataOut_payload_78,
  output     [7:0]    dataOut_payload_79,
  output     [7:0]    dataOut_payload_80,
  output     [7:0]    dataOut_payload_81,
  output     [7:0]    dataOut_payload_82,
  output     [7:0]    dataOut_payload_83,
  output     [7:0]    dataOut_payload_84,
  output     [7:0]    dataOut_payload_85,
  output     [7:0]    dataOut_payload_86,
  output     [7:0]    dataOut_payload_87,
  output     [7:0]    dataOut_payload_88,
  output     [7:0]    dataOut_payload_89,
  output     [7:0]    dataOut_payload_90,
  output     [7:0]    dataOut_payload_91,
  output     [7:0]    dataOut_payload_92,
  output     [7:0]    dataOut_payload_93,
  output     [7:0]    dataOut_payload_94,
  output     [7:0]    dataOut_payload_95,
  output     [7:0]    dataOut_payload_96,
  output     [7:0]    dataOut_payload_97,
  output     [7:0]    dataOut_payload_98,
  output     [7:0]    dataOut_payload_99,
  output     [7:0]    dataOut_payload_100,
  output     [7:0]    dataOut_payload_101,
  output     [7:0]    dataOut_payload_102,
  output     [7:0]    dataOut_payload_103,
  output     [7:0]    dataOut_payload_104,
  output     [7:0]    dataOut_payload_105,
  output     [7:0]    dataOut_payload_106,
  output     [7:0]    dataOut_payload_107,
  output     [7:0]    dataOut_payload_108,
  output     [7:0]    dataOut_payload_109,
  output     [7:0]    dataOut_payload_110,
  output     [7:0]    dataOut_payload_111,
  output     [7:0]    dataOut_payload_112,
  output     [7:0]    dataOut_payload_113,
  output     [7:0]    dataOut_payload_114,
  output     [7:0]    dataOut_payload_115,
  output     [7:0]    dataOut_payload_116,
  output     [7:0]    dataOut_payload_117,
  output     [7:0]    dataOut_payload_118,
  output     [7:0]    dataOut_payload_119,
  output     [7:0]    dataOut_payload_120,
  output     [7:0]    dataOut_payload_121,
  output     [7:0]    dataOut_payload_122,
  output     [7:0]    dataOut_payload_123,
  output     [7:0]    dataOut_payload_124,
  output     [7:0]    dataOut_payload_125,
  output     [7:0]    dataOut_payload_126,
  output     [7:0]    dataOut_payload_127,
  output     [7:0]    dataOut_payload_128,
  output     [7:0]    dataOut_payload_129,
  output     [7:0]    dataOut_payload_130,
  output     [7:0]    dataOut_payload_131,
  output     [7:0]    dataOut_payload_132,
  output     [7:0]    dataOut_payload_133,
  output     [7:0]    dataOut_payload_134,
  output     [7:0]    dataOut_payload_135,
  output     [7:0]    dataOut_payload_136,
  output     [7:0]    dataOut_payload_137,
  output     [7:0]    dataOut_payload_138,
  output     [7:0]    dataOut_payload_139,
  output     [7:0]    dataOut_payload_140,
  output     [7:0]    dataOut_payload_141,
  output     [7:0]    dataOut_payload_142,
  output     [7:0]    dataOut_payload_143,
  output     [7:0]    dataOut_payload_144,
  output     [7:0]    dataOut_payload_145,
  output     [7:0]    dataOut_payload_146,
  output     [7:0]    dataOut_payload_147,
  output     [7:0]    dataOut_payload_148,
  output     [7:0]    dataOut_payload_149,
  output     [7:0]    dataOut_payload_150,
  output     [7:0]    dataOut_payload_151,
  output     [7:0]    dataOut_payload_152,
  output     [7:0]    dataOut_payload_153,
  output     [7:0]    dataOut_payload_154,
  output     [7:0]    dataOut_payload_155,
  output     [7:0]    dataOut_payload_156,
  output     [7:0]    dataOut_payload_157,
  output     [7:0]    dataOut_payload_158,
  output     [7:0]    dataOut_payload_159,
  output     [7:0]    dataOut_payload_160,
  output     [7:0]    dataOut_payload_161,
  output     [7:0]    dataOut_payload_162,
  output     [7:0]    dataOut_payload_163,
  output     [7:0]    dataOut_payload_164,
  output     [7:0]    dataOut_payload_165,
  output     [7:0]    dataOut_payload_166,
  output     [7:0]    dataOut_payload_167,
  output     [7:0]    dataOut_payload_168,
  output     [7:0]    dataOut_payload_169,
  output     [7:0]    dataOut_payload_170,
  output     [7:0]    dataOut_payload_171,
  output     [7:0]    dataOut_payload_172,
  output     [7:0]    dataOut_payload_173,
  output     [7:0]    dataOut_payload_174,
  output     [7:0]    dataOut_payload_175,
  output     [7:0]    dataOut_payload_176,
  output     [7:0]    dataOut_payload_177,
  output     [7:0]    dataOut_payload_178,
  output     [7:0]    dataOut_payload_179,
  output     [7:0]    dataOut_payload_180,
  output     [7:0]    dataOut_payload_181,
  output     [7:0]    dataOut_payload_182,
  output     [7:0]    dataOut_payload_183,
  output     [7:0]    dataOut_payload_184,
  output     [7:0]    dataOut_payload_185,
  output     [7:0]    dataOut_payload_186,
  output     [7:0]    dataOut_payload_187,
  output     [7:0]    dataOut_payload_188,
  output     [7:0]    dataOut_payload_189,
  output     [7:0]    dataOut_payload_190,
  output     [7:0]    dataOut_payload_191,
  output     [7:0]    dataOut_payload_192,
  output     [7:0]    dataOut_payload_193,
  output     [7:0]    dataOut_payload_194,
  output     [7:0]    dataOut_payload_195,
  output     [7:0]    dataOut_payload_196,
  output     [7:0]    dataOut_payload_197,
  output     [7:0]    dataOut_payload_198,
  output     [7:0]    dataOut_payload_199,
  output     [7:0]    dataOut_payload_200,
  output     [7:0]    dataOut_payload_201,
  output     [7:0]    dataOut_payload_202,
  output     [7:0]    dataOut_payload_203,
  output     [7:0]    dataOut_payload_204,
  output     [7:0]    dataOut_payload_205,
  output     [7:0]    dataOut_payload_206,
  output     [7:0]    dataOut_payload_207,
  output     [7:0]    dataOut_payload_208,
  output     [7:0]    dataOut_payload_209,
  output     [7:0]    dataOut_payload_210,
  output     [7:0]    dataOut_payload_211,
  output     [7:0]    dataOut_payload_212,
  output     [7:0]    dataOut_payload_213,
  output     [7:0]    dataOut_payload_214,
  output     [7:0]    dataOut_payload_215,
  output     [7:0]    dataOut_payload_216,
  output     [7:0]    dataOut_payload_217,
  output     [7:0]    dataOut_payload_218,
  output     [7:0]    dataOut_payload_219,
  output     [7:0]    dataOut_payload_220,
  output     [7:0]    dataOut_payload_221,
  output     [7:0]    dataOut_payload_222,
  output     [7:0]    dataOut_payload_223,
  output     [7:0]    dataOut_payload_224,
  output     [7:0]    dataOut_payload_225,
  output     [7:0]    dataOut_payload_226,
  output     [7:0]    dataOut_payload_227,
  output     [7:0]    dataOut_payload_228,
  output     [7:0]    dataOut_payload_229,
  output     [7:0]    dataOut_payload_230,
  output     [7:0]    dataOut_payload_231,
  output     [7:0]    dataOut_payload_232,
  output     [7:0]    dataOut_payload_233,
  output     [7:0]    dataOut_payload_234,
  output     [7:0]    dataOut_payload_235,
  output     [7:0]    dataOut_payload_236,
  output     [7:0]    dataOut_payload_237,
  output     [7:0]    dataOut_payload_238,
  output     [7:0]    dataOut_payload_239,
  output     [7:0]    dataOut_payload_240,
  output     [7:0]    dataOut_payload_241,
  output     [7:0]    dataOut_payload_242,
  output     [7:0]    dataOut_payload_243,
  output     [7:0]    dataOut_payload_244,
  output     [7:0]    dataOut_payload_245,
  output     [7:0]    dataOut_payload_246,
  output     [7:0]    dataOut_payload_247,
  output     [7:0]    dataOut_payload_248,
  output     [7:0]    dataOut_payload_249,
  output     [7:0]    dataOut_payload_250,
  output     [7:0]    dataOut_payload_251,
  output     [7:0]    dataOut_payload_252,
  output     [7:0]    dataOut_payload_253,
  output     [7:0]    dataOut_payload_254,
  output     [7:0]    dataOut_payload_255,
  input               clk,
  input               reset
);

  wire                _zz_dataOut_payload_0;
  wire                _zz_dataOut_payload_0_1;
  wire                _zz_dataOut_payload_0_2;
  wire                _zz_dataOut_payload_0_3;
  wire                _zz_dataOut_payload_0_4;
  wire                _zz_dataOut_payload_0_5;
  wire                _zz_dataOut_payload_0_6;
  wire                _zz_dataOut_payload_0_7;
  wire                _zz_dataOut_payload_0_8;
  wire                _zz_dataOut_payload_0_9;
  wire                _zz_dataOut_payload_0_10;
  wire                _zz_dataOut_payload_0_11;
  wire                _zz_dataOut_payload_0_12;
  wire                _zz_dataOut_payload_0_13;
  wire                _zz_dataOut_payload_0_14;
  wire                _zz_dataOut_payload_0_15;
  wire                _zz_dataOut_payload_0_16;
  wire                _zz_dataOut_payload_0_17;
  wire                _zz_dataOut_payload_0_18;
  wire                _zz_dataOut_payload_0_19;
  wire                _zz_dataOut_payload_0_20;
  wire                _zz_dataOut_payload_0_21;
  wire                _zz_dataOut_payload_0_22;
  wire                _zz_dataOut_payload_0_23;
  wire                _zz_dataOut_payload_0_24;
  wire                _zz_dataOut_payload_0_25;
  wire                _zz_dataOut_payload_0_26;
  wire                _zz_dataOut_payload_0_27;
  wire                _zz_dataOut_payload_0_28;
  wire                _zz_dataOut_payload_0_29;
  wire                _zz_dataOut_payload_0_30;
  wire                _zz_dataOut_payload_0_31;
  wire                _zz_dataOut_payload_0_32;
  wire                _zz_dataOut_payload_0_33;
  wire                _zz_dataOut_payload_0_34;
  wire                _zz_dataOut_payload_0_35;
  wire                _zz_dataOut_payload_0_36;
  wire                _zz_dataOut_payload_0_37;
  wire                _zz_dataOut_payload_0_38;
  wire                _zz_dataOut_payload_0_39;
  wire                _zz_dataOut_payload_0_40;
  wire                _zz_dataOut_payload_0_41;
  wire                _zz_dataOut_payload_0_42;
  wire                _zz_dataOut_payload_0_43;
  wire                _zz_dataOut_payload_0_44;
  wire                _zz_dataOut_payload_0_45;
  wire                _zz_dataOut_payload_0_46;
  wire                _zz_dataOut_payload_0_47;
  wire                _zz_dataOut_payload_0_48;
  wire                _zz_dataOut_payload_0_49;
  wire                _zz_dataOut_payload_0_50;
  wire                _zz_dataOut_payload_0_51;
  wire                _zz_dataOut_payload_0_52;
  wire                _zz_dataOut_payload_0_53;
  wire                _zz_dataOut_payload_0_54;
  wire                _zz_dataOut_payload_0_55;
  wire                _zz_dataOut_payload_0_56;
  wire                _zz_dataOut_payload_0_57;
  wire                _zz_dataOut_payload_0_58;
  wire                _zz_dataOut_payload_0_59;
  wire                _zz_dataOut_payload_0_60;
  wire                _zz_dataOut_payload_0_61;
  wire                _zz_dataOut_payload_0_62;
  wire                _zz_dataOut_payload_0_63;
  wire                _zz_dataOut_payload_0_64;
  wire                _zz_dataOut_payload_0_65;
  wire                _zz_dataOut_payload_0_66;
  wire                _zz_dataOut_payload_0_67;
  wire                _zz_dataOut_payload_0_68;
  wire                _zz_dataOut_payload_0_69;
  wire                _zz_dataOut_payload_0_70;
  wire                _zz_dataOut_payload_0_71;
  wire                _zz_dataOut_payload_0_72;
  wire                _zz_dataOut_payload_0_73;
  wire                _zz_dataOut_payload_0_74;
  wire                _zz_dataOut_payload_0_75;
  wire                _zz_dataOut_payload_0_76;
  wire                _zz_dataOut_payload_0_77;
  wire                _zz_dataOut_payload_0_78;
  wire                _zz_dataOut_payload_0_79;
  wire                _zz_dataOut_payload_0_80;
  wire                _zz_dataOut_payload_0_81;
  wire                _zz_dataOut_payload_0_82;
  wire                _zz_dataOut_payload_0_83;
  wire                _zz_dataOut_payload_0_84;
  wire                _zz_dataOut_payload_0_85;
  wire                _zz_dataOut_payload_0_86;
  wire                _zz_dataOut_payload_0_87;
  wire                _zz_dataOut_payload_0_88;
  wire                _zz_dataOut_payload_0_89;
  wire                _zz_dataOut_payload_0_90;
  wire                _zz_dataOut_payload_0_91;
  wire                _zz_dataOut_payload_0_92;
  wire                _zz_dataOut_payload_0_93;
  wire                _zz_dataOut_payload_0_94;
  wire                _zz_dataOut_payload_0_95;
  wire                _zz_dataOut_payload_0_96;
  wire                _zz_dataOut_payload_0_97;
  wire                _zz_dataOut_payload_0_98;
  wire                _zz_dataOut_payload_0_99;
  wire                _zz_dataOut_payload_0_100;
  wire                _zz_dataOut_payload_0_101;
  wire                _zz_dataOut_payload_0_102;
  wire                _zz_dataOut_payload_0_103;
  wire                _zz_dataOut_payload_0_104;
  wire                _zz_dataOut_payload_0_105;
  wire                _zz_dataOut_payload_0_106;
  wire                _zz_dataOut_payload_0_107;
  wire                _zz_dataOut_payload_0_108;
  wire                _zz_dataOut_payload_0_109;
  wire                _zz_dataOut_payload_0_110;
  wire                _zz_dataOut_payload_0_111;
  wire                _zz_dataOut_payload_0_112;
  wire                _zz_dataOut_payload_0_113;
  wire                _zz_dataOut_payload_0_114;
  wire                _zz_dataOut_payload_0_115;
  wire                _zz_dataOut_payload_0_116;
  wire                _zz_dataOut_payload_0_117;
  wire                _zz_dataOut_payload_0_118;
  wire                _zz_dataOut_payload_0_119;
  wire                _zz_dataOut_payload_0_120;
  wire                _zz_dataOut_payload_0_121;
  wire                _zz_dataOut_payload_0_122;
  wire                _zz_dataOut_payload_0_123;
  wire                _zz_dataOut_payload_0_124;
  wire                _zz_dataOut_payload_0_125;
  wire                _zz_dataOut_payload_0_126;
  wire                _zz_dataOut_payload_0_127;
  reg        [7:0]    _zz_dataOut_payload_0_128;
  reg        [7:0]    _zz_dataOut_payload_0_129;
  reg        [7:0]    _zz_dataOut_payload_0_130;
  reg        [7:0]    _zz_dataOut_payload_0_131;
  reg        [7:0]    _zz_dataOut_payload_0_132;
  reg        [7:0]    _zz_dataOut_payload_0_133;
  reg        [7:0]    _zz_dataOut_payload_0_134;
  reg        [7:0]    _zz_dataOut_payload_0_135;
  reg        [7:0]    _zz_dataOut_payload_0_136;
  reg        [7:0]    _zz_dataOut_payload_0_137;
  reg        [7:0]    _zz_dataOut_payload_0_138;
  reg        [7:0]    _zz_dataOut_payload_0_139;
  reg        [7:0]    _zz_dataOut_payload_0_140;
  reg        [7:0]    _zz_dataOut_payload_0_141;
  reg        [7:0]    _zz_dataOut_payload_0_142;
  reg        [7:0]    _zz_dataOut_payload_0_143;
  reg        [7:0]    _zz_dataOut_payload_0_144;
  reg        [7:0]    _zz_dataOut_payload_0_145;
  reg        [7:0]    _zz_dataOut_payload_0_146;
  reg        [7:0]    _zz_dataOut_payload_0_147;
  reg        [7:0]    _zz_dataOut_payload_0_148;
  reg        [7:0]    _zz_dataOut_payload_0_149;
  reg        [7:0]    _zz_dataOut_payload_0_150;
  reg        [7:0]    _zz_dataOut_payload_0_151;
  reg        [7:0]    _zz_dataOut_payload_0_152;
  reg        [7:0]    _zz_dataOut_payload_0_153;
  reg        [7:0]    _zz_dataOut_payload_0_154;
  reg        [7:0]    _zz_dataOut_payload_0_155;
  reg        [7:0]    _zz_dataOut_payload_0_156;
  reg        [7:0]    _zz_dataOut_payload_0_157;
  reg        [7:0]    _zz_dataOut_payload_0_158;
  reg        [7:0]    _zz_dataOut_payload_0_159;
  reg        [7:0]    _zz_dataOut_payload_0_160;
  reg        [7:0]    _zz_dataOut_payload_0_161;
  reg        [7:0]    _zz_dataOut_payload_0_162;
  reg        [7:0]    _zz_dataOut_payload_0_163;
  reg        [7:0]    _zz_dataOut_payload_0_164;
  reg        [7:0]    _zz_dataOut_payload_0_165;
  reg        [7:0]    _zz_dataOut_payload_0_166;
  reg        [7:0]    _zz_dataOut_payload_0_167;
  reg        [7:0]    _zz_dataOut_payload_0_168;
  reg        [7:0]    _zz_dataOut_payload_0_169;
  reg        [7:0]    _zz_dataOut_payload_0_170;
  reg        [7:0]    _zz_dataOut_payload_0_171;
  reg        [7:0]    _zz_dataOut_payload_0_172;
  reg        [7:0]    _zz_dataOut_payload_0_173;
  reg        [7:0]    _zz_dataOut_payload_0_174;
  reg        [7:0]    _zz_dataOut_payload_0_175;
  reg        [7:0]    _zz_dataOut_payload_0_176;
  reg        [7:0]    _zz_dataOut_payload_0_177;
  reg        [7:0]    _zz_dataOut_payload_0_178;
  reg        [7:0]    _zz_dataOut_payload_0_179;
  reg        [7:0]    _zz_dataOut_payload_0_180;
  reg        [7:0]    _zz_dataOut_payload_0_181;
  reg        [7:0]    _zz_dataOut_payload_0_182;
  reg        [7:0]    _zz_dataOut_payload_0_183;
  reg        [7:0]    _zz_dataOut_payload_0_184;
  reg        [7:0]    _zz_dataOut_payload_0_185;
  reg        [7:0]    _zz_dataOut_payload_0_186;
  reg        [7:0]    _zz_dataOut_payload_0_187;
  reg        [7:0]    _zz_dataOut_payload_0_188;
  reg        [7:0]    _zz_dataOut_payload_0_189;
  reg        [7:0]    _zz_dataOut_payload_0_190;
  reg        [7:0]    _zz_dataOut_payload_0_191;
  reg        [7:0]    _zz_dataOut_payload_0_192;
  reg        [7:0]    _zz_dataOut_payload_0_193;
  reg        [7:0]    _zz_dataOut_payload_0_194;
  reg        [7:0]    _zz_dataOut_payload_0_195;
  reg        [7:0]    _zz_dataOut_payload_0_196;
  reg        [7:0]    _zz_dataOut_payload_0_197;
  reg        [7:0]    _zz_dataOut_payload_0_198;
  reg        [7:0]    _zz_dataOut_payload_0_199;
  reg        [7:0]    _zz_dataOut_payload_0_200;
  reg        [7:0]    _zz_dataOut_payload_0_201;
  reg        [7:0]    _zz_dataOut_payload_0_202;
  reg        [7:0]    _zz_dataOut_payload_0_203;
  reg        [7:0]    _zz_dataOut_payload_0_204;
  reg        [7:0]    _zz_dataOut_payload_0_205;
  reg        [7:0]    _zz_dataOut_payload_0_206;
  reg        [7:0]    _zz_dataOut_payload_0_207;
  reg        [7:0]    _zz_dataOut_payload_0_208;
  reg        [7:0]    _zz_dataOut_payload_0_209;
  reg        [7:0]    _zz_dataOut_payload_0_210;
  reg        [7:0]    _zz_dataOut_payload_0_211;
  reg        [7:0]    _zz_dataOut_payload_0_212;
  reg        [7:0]    _zz_dataOut_payload_0_213;
  reg        [7:0]    _zz_dataOut_payload_0_214;
  reg        [7:0]    _zz_dataOut_payload_0_215;
  reg        [7:0]    _zz_dataOut_payload_0_216;
  reg        [7:0]    _zz_dataOut_payload_0_217;
  reg        [7:0]    _zz_dataOut_payload_0_218;
  reg        [7:0]    _zz_dataOut_payload_0_219;
  reg        [7:0]    _zz_dataOut_payload_0_220;
  reg        [7:0]    _zz_dataOut_payload_0_221;
  reg        [7:0]    _zz_dataOut_payload_0_222;
  reg        [7:0]    _zz_dataOut_payload_0_223;
  reg        [7:0]    _zz_dataOut_payload_0_224;
  reg        [7:0]    _zz_dataOut_payload_0_225;
  reg        [7:0]    _zz_dataOut_payload_0_226;
  reg        [7:0]    _zz_dataOut_payload_0_227;
  reg        [7:0]    _zz_dataOut_payload_0_228;
  reg        [7:0]    _zz_dataOut_payload_0_229;
  reg        [7:0]    _zz_dataOut_payload_0_230;
  reg        [7:0]    _zz_dataOut_payload_0_231;
  reg        [7:0]    _zz_dataOut_payload_0_232;
  reg        [7:0]    _zz_dataOut_payload_0_233;
  reg        [7:0]    _zz_dataOut_payload_0_234;
  reg        [7:0]    _zz_dataOut_payload_0_235;
  reg        [7:0]    _zz_dataOut_payload_0_236;
  reg        [7:0]    _zz_dataOut_payload_0_237;
  reg        [7:0]    _zz_dataOut_payload_0_238;
  reg        [7:0]    _zz_dataOut_payload_0_239;
  reg        [7:0]    _zz_dataOut_payload_0_240;
  reg        [7:0]    _zz_dataOut_payload_0_241;
  reg        [7:0]    _zz_dataOut_payload_0_242;
  reg        [7:0]    _zz_dataOut_payload_0_243;
  reg        [7:0]    _zz_dataOut_payload_0_244;
  reg        [7:0]    _zz_dataOut_payload_0_245;
  reg        [7:0]    _zz_dataOut_payload_0_246;
  reg        [7:0]    _zz_dataOut_payload_0_247;
  reg        [7:0]    _zz_dataOut_payload_0_248;
  reg        [7:0]    _zz_dataOut_payload_0_249;
  reg        [7:0]    _zz_dataOut_payload_0_250;
  reg        [7:0]    _zz_dataOut_payload_0_251;
  reg        [7:0]    _zz_dataOut_payload_0_252;
  reg        [7:0]    _zz_dataOut_payload_0_253;
  reg        [7:0]    _zz_dataOut_payload_0_254;
  reg        [7:0]    _zz_dataOut_payload_0_255;
  reg        [7:0]    _zz_dataOut_payload_0_256;
  reg        [7:0]    _zz_dataOut_payload_0_257;
  reg        [7:0]    _zz_dataOut_payload_0_258;
  reg        [7:0]    _zz_dataOut_payload_0_259;
  reg        [7:0]    _zz_dataOut_payload_0_260;
  reg        [7:0]    _zz_dataOut_payload_0_261;
  reg        [7:0]    _zz_dataOut_payload_0_262;
  reg        [7:0]    _zz_dataOut_payload_0_263;
  reg        [7:0]    _zz_dataOut_payload_0_264;
  reg        [7:0]    _zz_dataOut_payload_0_265;
  reg        [7:0]    _zz_dataOut_payload_0_266;
  reg        [7:0]    _zz_dataOut_payload_0_267;
  reg        [7:0]    _zz_dataOut_payload_0_268;
  reg        [7:0]    _zz_dataOut_payload_0_269;
  reg        [7:0]    _zz_dataOut_payload_0_270;
  reg        [7:0]    _zz_dataOut_payload_0_271;
  reg        [7:0]    _zz_dataOut_payload_0_272;
  reg        [7:0]    _zz_dataOut_payload_0_273;
  reg        [7:0]    _zz_dataOut_payload_0_274;
  reg        [7:0]    _zz_dataOut_payload_0_275;
  reg        [7:0]    _zz_dataOut_payload_0_276;
  reg        [7:0]    _zz_dataOut_payload_0_277;
  reg        [7:0]    _zz_dataOut_payload_0_278;
  reg        [7:0]    _zz_dataOut_payload_0_279;
  reg        [7:0]    _zz_dataOut_payload_0_280;
  reg        [7:0]    _zz_dataOut_payload_0_281;
  reg        [7:0]    _zz_dataOut_payload_0_282;
  reg        [7:0]    _zz_dataOut_payload_0_283;
  reg        [7:0]    _zz_dataOut_payload_0_284;
  reg        [7:0]    _zz_dataOut_payload_0_285;
  reg        [7:0]    _zz_dataOut_payload_0_286;
  reg        [7:0]    _zz_dataOut_payload_0_287;
  reg        [7:0]    _zz_dataOut_payload_0_288;
  reg        [7:0]    _zz_dataOut_payload_0_289;
  reg        [7:0]    _zz_dataOut_payload_0_290;
  reg        [7:0]    _zz_dataOut_payload_0_291;
  reg        [7:0]    _zz_dataOut_payload_0_292;
  reg        [7:0]    _zz_dataOut_payload_0_293;
  reg        [7:0]    _zz_dataOut_payload_0_294;
  reg        [7:0]    _zz_dataOut_payload_0_295;
  reg        [7:0]    _zz_dataOut_payload_0_296;
  reg        [7:0]    _zz_dataOut_payload_0_297;
  reg        [7:0]    _zz_dataOut_payload_0_298;
  reg        [7:0]    _zz_dataOut_payload_0_299;
  reg        [7:0]    _zz_dataOut_payload_0_300;
  reg        [7:0]    _zz_dataOut_payload_0_301;
  reg        [7:0]    _zz_dataOut_payload_0_302;
  reg        [7:0]    _zz_dataOut_payload_0_303;
  reg        [7:0]    _zz_dataOut_payload_0_304;
  reg        [7:0]    _zz_dataOut_payload_0_305;
  reg        [7:0]    _zz_dataOut_payload_0_306;
  reg        [7:0]    _zz_dataOut_payload_0_307;
  reg        [7:0]    _zz_dataOut_payload_0_308;
  reg        [7:0]    _zz_dataOut_payload_0_309;
  reg        [7:0]    _zz_dataOut_payload_0_310;
  reg        [7:0]    _zz_dataOut_payload_0_311;
  reg        [7:0]    _zz_dataOut_payload_0_312;
  reg        [7:0]    _zz_dataOut_payload_0_313;
  reg        [7:0]    _zz_dataOut_payload_0_314;
  reg        [7:0]    _zz_dataOut_payload_0_315;
  reg        [7:0]    _zz_dataOut_payload_0_316;
  reg        [7:0]    _zz_dataOut_payload_0_317;
  reg        [7:0]    _zz_dataOut_payload_0_318;
  reg        [7:0]    _zz_dataOut_payload_0_319;
  reg        [7:0]    _zz_dataOut_payload_0_320;
  reg        [7:0]    _zz_dataOut_payload_0_321;
  reg        [7:0]    _zz_dataOut_payload_0_322;
  reg        [7:0]    _zz_dataOut_payload_0_323;
  reg        [7:0]    _zz_dataOut_payload_0_324;
  reg        [7:0]    _zz_dataOut_payload_0_325;
  reg        [7:0]    _zz_dataOut_payload_0_326;
  reg        [7:0]    _zz_dataOut_payload_0_327;
  reg        [7:0]    _zz_dataOut_payload_0_328;
  reg        [7:0]    _zz_dataOut_payload_0_329;
  reg        [7:0]    _zz_dataOut_payload_0_330;
  reg        [7:0]    _zz_dataOut_payload_0_331;
  reg        [7:0]    _zz_dataOut_payload_0_332;
  reg        [7:0]    _zz_dataOut_payload_0_333;
  reg        [7:0]    _zz_dataOut_payload_0_334;
  reg        [7:0]    _zz_dataOut_payload_0_335;
  reg        [7:0]    _zz_dataOut_payload_0_336;
  reg        [7:0]    _zz_dataOut_payload_0_337;
  reg        [7:0]    _zz_dataOut_payload_0_338;
  reg        [7:0]    _zz_dataOut_payload_0_339;
  reg        [7:0]    _zz_dataOut_payload_0_340;
  reg        [7:0]    _zz_dataOut_payload_0_341;
  reg        [7:0]    _zz_dataOut_payload_0_342;
  reg        [7:0]    _zz_dataOut_payload_0_343;
  reg        [7:0]    _zz_dataOut_payload_0_344;
  reg        [7:0]    _zz_dataOut_payload_0_345;
  reg        [7:0]    _zz_dataOut_payload_0_346;
  reg        [7:0]    _zz_dataOut_payload_0_347;
  reg        [7:0]    _zz_dataOut_payload_0_348;
  reg        [7:0]    _zz_dataOut_payload_0_349;
  reg        [7:0]    _zz_dataOut_payload_0_350;
  reg        [7:0]    _zz_dataOut_payload_0_351;
  reg        [7:0]    _zz_dataOut_payload_0_352;
  reg        [7:0]    _zz_dataOut_payload_0_353;
  reg        [7:0]    _zz_dataOut_payload_0_354;
  reg        [7:0]    _zz_dataOut_payload_0_355;
  reg        [7:0]    _zz_dataOut_payload_0_356;
  reg        [7:0]    _zz_dataOut_payload_0_357;
  reg        [7:0]    _zz_dataOut_payload_0_358;
  reg        [7:0]    _zz_dataOut_payload_0_359;
  reg        [7:0]    _zz_dataOut_payload_0_360;
  reg        [7:0]    _zz_dataOut_payload_0_361;
  reg        [7:0]    _zz_dataOut_payload_0_362;
  reg        [7:0]    _zz_dataOut_payload_0_363;
  reg        [7:0]    _zz_dataOut_payload_0_364;
  reg        [7:0]    _zz_dataOut_payload_0_365;
  reg        [7:0]    _zz_dataOut_payload_0_366;
  reg        [7:0]    _zz_dataOut_payload_0_367;
  reg        [7:0]    _zz_dataOut_payload_0_368;
  reg        [7:0]    _zz_dataOut_payload_0_369;
  reg        [7:0]    _zz_dataOut_payload_0_370;
  reg        [7:0]    _zz_dataOut_payload_0_371;
  reg        [7:0]    _zz_dataOut_payload_0_372;
  reg        [7:0]    _zz_dataOut_payload_0_373;
  reg        [7:0]    _zz_dataOut_payload_0_374;
  reg        [7:0]    _zz_dataOut_payload_0_375;
  reg        [7:0]    _zz_dataOut_payload_0_376;
  reg        [7:0]    _zz_dataOut_payload_0_377;
  reg        [7:0]    _zz_dataOut_payload_0_378;
  reg        [7:0]    _zz_dataOut_payload_0_379;
  reg        [7:0]    _zz_dataOut_payload_0_380;
  reg        [7:0]    _zz_dataOut_payload_0_381;
  reg        [7:0]    _zz_dataOut_payload_0_382;
  reg        [7:0]    _zz_dataOut_payload_0_383;
  wire                _zz_dataOut_payload_0_384;
  wire       [7:0]    _zz_dataOut_payload_0_385;
  wire       [7:0]    _zz_dataOut_payload_0_386;
  wire                _zz_dataOut_payload_0_387;
  wire       [7:0]    _zz_dataOut_payload_0_388;
  wire       [7:0]    _zz_dataOut_payload_0_389;
  wire                _zz_dataOut_payload_0_390;
  wire                _zz_dataOut_payload_0_391;
  reg        [7:0]    _zz_dataOut_payload_0_392;
  reg        [7:0]    _zz_dataOut_payload_0_393;
  reg        [7:0]    _zz_dataOut_payload_0_394;
  reg        [7:0]    _zz_dataOut_payload_0_395;
  wire                _zz_dataOut_payload_0_396;
  wire       [7:0]    _zz_dataOut_payload_0_397;
  wire       [7:0]    _zz_dataOut_payload_0_398;
  wire                _zz_dataOut_payload_0_399;
  wire       [7:0]    _zz_dataOut_payload_0_400;
  wire       [7:0]    _zz_dataOut_payload_0_401;
  wire                _zz_dataOut_payload_0_402;
  wire                _zz_dataOut_payload_0_403;
  reg        [7:0]    _zz_dataOut_payload_0_404;
  reg        [7:0]    _zz_dataOut_payload_0_405;
  reg        [7:0]    _zz_dataOut_payload_0_406;
  reg        [7:0]    _zz_dataOut_payload_0_407;
  wire                _zz_dataOut_payload_0_408;
  wire       [7:0]    _zz_dataOut_payload_0_409;
  wire       [7:0]    _zz_dataOut_payload_0_410;
  wire                _zz_dataOut_payload_0_411;
  wire       [7:0]    _zz_dataOut_payload_0_412;
  wire       [7:0]    _zz_dataOut_payload_0_413;
  wire                _zz_dataOut_payload_0_414;
  wire                _zz_dataOut_payload_0_415;
  reg        [7:0]    _zz_dataOut_payload_0_416;
  reg        [7:0]    _zz_dataOut_payload_0_417;
  reg        [7:0]    _zz_dataOut_payload_0_418;
  reg        [7:0]    _zz_dataOut_payload_0_419;
  wire                _zz_dataOut_payload_0_420;
  wire       [7:0]    _zz_dataOut_payload_0_421;
  wire       [7:0]    _zz_dataOut_payload_0_422;
  wire                _zz_dataOut_payload_0_423;
  wire       [7:0]    _zz_dataOut_payload_0_424;
  wire       [7:0]    _zz_dataOut_payload_0_425;
  wire                _zz_dataOut_payload_0_426;
  wire                _zz_dataOut_payload_0_427;
  reg        [7:0]    _zz_dataOut_payload_0_428;
  reg        [7:0]    _zz_dataOut_payload_0_429;
  reg        [7:0]    _zz_dataOut_payload_0_430;
  reg        [7:0]    _zz_dataOut_payload_0_431;
  wire                _zz_dataOut_payload_0_432;
  wire       [7:0]    _zz_dataOut_payload_0_433;
  wire       [7:0]    _zz_dataOut_payload_0_434;
  wire                _zz_dataOut_payload_0_435;
  wire       [7:0]    _zz_dataOut_payload_0_436;
  wire       [7:0]    _zz_dataOut_payload_0_437;
  wire                _zz_dataOut_payload_0_438;
  wire                _zz_dataOut_payload_0_439;
  reg        [7:0]    _zz_dataOut_payload_0_440;
  reg        [7:0]    _zz_dataOut_payload_0_441;
  reg        [7:0]    _zz_dataOut_payload_0_442;
  reg        [7:0]    _zz_dataOut_payload_0_443;
  wire                _zz_dataOut_payload_0_444;
  wire       [7:0]    _zz_dataOut_payload_0_445;
  wire       [7:0]    _zz_dataOut_payload_0_446;
  wire                _zz_dataOut_payload_0_447;
  wire       [7:0]    _zz_dataOut_payload_0_448;
  wire       [7:0]    _zz_dataOut_payload_0_449;
  wire                _zz_dataOut_payload_0_450;
  wire                _zz_dataOut_payload_0_451;
  reg        [7:0]    _zz_dataOut_payload_0_452;
  reg        [7:0]    _zz_dataOut_payload_0_453;
  reg        [7:0]    _zz_dataOut_payload_0_454;
  reg        [7:0]    _zz_dataOut_payload_0_455;
  wire                _zz_dataOut_payload_0_456;
  wire       [7:0]    _zz_dataOut_payload_0_457;
  wire       [7:0]    _zz_dataOut_payload_0_458;
  wire                _zz_dataOut_payload_0_459;
  wire       [7:0]    _zz_dataOut_payload_0_460;
  wire       [7:0]    _zz_dataOut_payload_0_461;
  wire                _zz_dataOut_payload_0_462;
  wire                _zz_dataOut_payload_0_463;
  reg        [7:0]    _zz_dataOut_payload_0_464;
  reg        [7:0]    _zz_dataOut_payload_0_465;
  reg        [7:0]    _zz_dataOut_payload_0_466;
  reg        [7:0]    _zz_dataOut_payload_0_467;
  wire                _zz_dataOut_payload_0_468;
  wire       [7:0]    _zz_dataOut_payload_0_469;
  wire       [7:0]    _zz_dataOut_payload_0_470;
  wire                _zz_dataOut_payload_0_471;
  wire       [7:0]    _zz_dataOut_payload_0_472;
  wire       [7:0]    _zz_dataOut_payload_0_473;
  wire                _zz_dataOut_payload_0_474;
  wire                _zz_dataOut_payload_0_475;
  reg        [7:0]    _zz_dataOut_payload_0_476;
  reg        [7:0]    _zz_dataOut_payload_0_477;
  reg        [7:0]    _zz_dataOut_payload_0_478;
  reg        [7:0]    _zz_dataOut_payload_0_479;
  wire                _zz_dataOut_payload_0_480;
  wire       [7:0]    _zz_dataOut_payload_0_481;
  wire       [7:0]    _zz_dataOut_payload_0_482;
  wire                _zz_dataOut_payload_0_483;
  wire       [7:0]    _zz_dataOut_payload_0_484;
  wire       [7:0]    _zz_dataOut_payload_0_485;
  wire                _zz_dataOut_payload_0_486;
  wire                _zz_dataOut_payload_0_487;
  reg        [7:0]    _zz_dataOut_payload_0_488;
  reg        [7:0]    _zz_dataOut_payload_0_489;
  reg        [7:0]    _zz_dataOut_payload_0_490;
  reg        [7:0]    _zz_dataOut_payload_0_491;
  wire                _zz_dataOut_payload_0_492;
  wire       [7:0]    _zz_dataOut_payload_0_493;
  wire       [7:0]    _zz_dataOut_payload_0_494;
  wire                _zz_dataOut_payload_0_495;
  wire       [7:0]    _zz_dataOut_payload_0_496;
  wire       [7:0]    _zz_dataOut_payload_0_497;
  wire                _zz_dataOut_payload_0_498;
  wire                _zz_dataOut_payload_0_499;
  reg        [7:0]    _zz_dataOut_payload_0_500;
  reg        [7:0]    _zz_dataOut_payload_0_501;
  reg        [7:0]    _zz_dataOut_payload_0_502;
  reg        [7:0]    _zz_dataOut_payload_0_503;
  wire                _zz_dataOut_payload_0_504;
  wire       [7:0]    _zz_dataOut_payload_0_505;
  wire       [7:0]    _zz_dataOut_payload_0_506;
  wire                _zz_dataOut_payload_0_507;
  wire       [7:0]    _zz_dataOut_payload_0_508;
  wire       [7:0]    _zz_dataOut_payload_0_509;
  wire                _zz_dataOut_payload_0_510;
  wire                _zz_dataOut_payload_0_511;
  reg        [7:0]    _zz_dataOut_payload_0_512;
  reg        [7:0]    _zz_dataOut_payload_0_513;
  reg        [7:0]    _zz_dataOut_payload_0_514;
  reg        [7:0]    _zz_dataOut_payload_0_515;
  wire                _zz_dataOut_payload_0_516;
  wire       [7:0]    _zz_dataOut_payload_0_517;
  wire       [7:0]    _zz_dataOut_payload_0_518;
  wire                _zz_dataOut_payload_0_519;
  wire       [7:0]    _zz_dataOut_payload_0_520;
  wire       [7:0]    _zz_dataOut_payload_0_521;
  wire                _zz_dataOut_payload_0_522;
  wire                _zz_dataOut_payload_0_523;
  reg        [7:0]    _zz_dataOut_payload_0_524;
  reg        [7:0]    _zz_dataOut_payload_0_525;
  reg        [7:0]    _zz_dataOut_payload_0_526;
  reg        [7:0]    _zz_dataOut_payload_0_527;
  wire                _zz_dataOut_payload_0_528;
  wire       [7:0]    _zz_dataOut_payload_0_529;
  wire       [7:0]    _zz_dataOut_payload_0_530;
  wire                _zz_dataOut_payload_0_531;
  wire       [7:0]    _zz_dataOut_payload_0_532;
  wire       [7:0]    _zz_dataOut_payload_0_533;
  wire                _zz_dataOut_payload_0_534;
  wire                _zz_dataOut_payload_0_535;
  reg        [7:0]    _zz_dataOut_payload_0_536;
  reg        [7:0]    _zz_dataOut_payload_0_537;
  reg        [7:0]    _zz_dataOut_payload_0_538;
  reg        [7:0]    _zz_dataOut_payload_0_539;
  wire                _zz_dataOut_payload_0_540;
  wire       [7:0]    _zz_dataOut_payload_0_541;
  wire       [7:0]    _zz_dataOut_payload_0_542;
  wire                _zz_dataOut_payload_0_543;
  wire       [7:0]    _zz_dataOut_payload_0_544;
  wire       [7:0]    _zz_dataOut_payload_0_545;
  wire                _zz_dataOut_payload_0_546;
  wire                _zz_dataOut_payload_0_547;
  reg        [7:0]    _zz_dataOut_payload_0_548;
  reg        [7:0]    _zz_dataOut_payload_0_549;
  reg        [7:0]    _zz_dataOut_payload_0_550;
  reg        [7:0]    _zz_dataOut_payload_0_551;
  wire                _zz_dataOut_payload_0_552;
  wire       [7:0]    _zz_dataOut_payload_0_553;
  wire       [7:0]    _zz_dataOut_payload_0_554;
  wire                _zz_dataOut_payload_0_555;
  wire       [7:0]    _zz_dataOut_payload_0_556;
  wire       [7:0]    _zz_dataOut_payload_0_557;
  wire                _zz_dataOut_payload_0_558;
  wire                _zz_dataOut_payload_0_559;
  reg        [7:0]    _zz_dataOut_payload_0_560;
  reg        [7:0]    _zz_dataOut_payload_0_561;
  reg        [7:0]    _zz_dataOut_payload_0_562;
  reg        [7:0]    _zz_dataOut_payload_0_563;
  wire                _zz_dataOut_payload_0_564;
  wire       [7:0]    _zz_dataOut_payload_0_565;
  wire       [7:0]    _zz_dataOut_payload_0_566;
  wire                _zz_dataOut_payload_0_567;
  wire       [7:0]    _zz_dataOut_payload_0_568;
  wire       [7:0]    _zz_dataOut_payload_0_569;
  wire                _zz_dataOut_payload_0_570;
  wire                _zz_dataOut_payload_0_571;
  reg        [7:0]    _zz_dataOut_payload_0_572;
  reg        [7:0]    _zz_dataOut_payload_0_573;
  reg        [7:0]    _zz_dataOut_payload_0_574;
  reg        [7:0]    _zz_dataOut_payload_0_575;
  wire                _zz_dataOut_payload_0_576;
  wire       [7:0]    _zz_dataOut_payload_0_577;
  wire       [7:0]    _zz_dataOut_payload_0_578;
  wire                _zz_dataOut_payload_0_579;
  wire       [7:0]    _zz_dataOut_payload_0_580;
  wire       [7:0]    _zz_dataOut_payload_0_581;
  wire                _zz_dataOut_payload_0_582;
  wire                _zz_dataOut_payload_0_583;
  reg        [7:0]    _zz_dataOut_payload_0_584;
  reg        [7:0]    _zz_dataOut_payload_0_585;
  reg        [7:0]    _zz_dataOut_payload_0_586;
  reg        [7:0]    _zz_dataOut_payload_0_587;
  wire                _zz_dataOut_payload_0_588;
  wire       [7:0]    _zz_dataOut_payload_0_589;
  wire       [7:0]    _zz_dataOut_payload_0_590;
  wire                _zz_dataOut_payload_0_591;
  wire       [7:0]    _zz_dataOut_payload_0_592;
  wire       [7:0]    _zz_dataOut_payload_0_593;
  wire                _zz_dataOut_payload_0_594;
  wire                _zz_dataOut_payload_0_595;
  reg        [7:0]    _zz_dataOut_payload_0_596;
  reg        [7:0]    _zz_dataOut_payload_0_597;
  reg        [7:0]    _zz_dataOut_payload_0_598;
  reg        [7:0]    _zz_dataOut_payload_0_599;
  wire                _zz_dataOut_payload_0_600;
  wire       [7:0]    _zz_dataOut_payload_0_601;
  wire       [7:0]    _zz_dataOut_payload_0_602;
  wire                _zz_dataOut_payload_0_603;
  wire       [7:0]    _zz_dataOut_payload_0_604;
  wire       [7:0]    _zz_dataOut_payload_0_605;
  wire                _zz_dataOut_payload_0_606;
  wire                _zz_dataOut_payload_0_607;
  reg        [7:0]    _zz_dataOut_payload_0_608;
  reg        [7:0]    _zz_dataOut_payload_0_609;
  reg        [7:0]    _zz_dataOut_payload_0_610;
  reg        [7:0]    _zz_dataOut_payload_0_611;
  wire                _zz_dataOut_payload_0_612;
  wire       [7:0]    _zz_dataOut_payload_0_613;
  wire       [7:0]    _zz_dataOut_payload_0_614;
  wire                _zz_dataOut_payload_0_615;
  wire       [7:0]    _zz_dataOut_payload_0_616;
  wire       [7:0]    _zz_dataOut_payload_0_617;
  wire                _zz_dataOut_payload_0_618;
  wire                _zz_dataOut_payload_0_619;
  reg        [7:0]    _zz_dataOut_payload_0_620;
  reg        [7:0]    _zz_dataOut_payload_0_621;
  reg        [7:0]    _zz_dataOut_payload_0_622;
  reg        [7:0]    _zz_dataOut_payload_0_623;
  wire                _zz_dataOut_payload_0_624;
  wire       [7:0]    _zz_dataOut_payload_0_625;
  wire       [7:0]    _zz_dataOut_payload_0_626;
  wire                _zz_dataOut_payload_0_627;
  wire       [7:0]    _zz_dataOut_payload_0_628;
  wire       [7:0]    _zz_dataOut_payload_0_629;
  wire                _zz_dataOut_payload_0_630;
  wire                _zz_dataOut_payload_0_631;
  reg        [7:0]    _zz_dataOut_payload_0_632;
  reg        [7:0]    _zz_dataOut_payload_0_633;
  reg        [7:0]    _zz_dataOut_payload_0_634;
  reg        [7:0]    _zz_dataOut_payload_0_635;
  wire                _zz_dataOut_payload_0_636;
  wire       [7:0]    _zz_dataOut_payload_0_637;
  wire       [7:0]    _zz_dataOut_payload_0_638;
  wire                _zz_dataOut_payload_0_639;
  wire       [7:0]    _zz_dataOut_payload_0_640;
  wire       [7:0]    _zz_dataOut_payload_0_641;
  wire                _zz_dataOut_payload_0_642;
  wire                _zz_dataOut_payload_0_643;
  reg        [7:0]    _zz_dataOut_payload_0_644;
  reg        [7:0]    _zz_dataOut_payload_0_645;
  reg        [7:0]    _zz_dataOut_payload_0_646;
  reg        [7:0]    _zz_dataOut_payload_0_647;
  wire                _zz_dataOut_payload_0_648;
  wire       [7:0]    _zz_dataOut_payload_0_649;
  wire       [7:0]    _zz_dataOut_payload_0_650;
  wire                _zz_dataOut_payload_0_651;
  wire       [7:0]    _zz_dataOut_payload_0_652;
  wire       [7:0]    _zz_dataOut_payload_0_653;
  wire                _zz_dataOut_payload_0_654;
  wire                _zz_dataOut_payload_0_655;
  reg        [7:0]    _zz_dataOut_payload_0_656;
  reg        [7:0]    _zz_dataOut_payload_0_657;
  reg        [7:0]    _zz_dataOut_payload_0_658;
  reg        [7:0]    _zz_dataOut_payload_0_659;
  wire                _zz_dataOut_payload_0_660;
  wire       [7:0]    _zz_dataOut_payload_0_661;
  wire       [7:0]    _zz_dataOut_payload_0_662;
  wire                _zz_dataOut_payload_0_663;
  wire       [7:0]    _zz_dataOut_payload_0_664;
  wire       [7:0]    _zz_dataOut_payload_0_665;
  wire                _zz_dataOut_payload_0_666;
  wire                _zz_dataOut_payload_0_667;
  reg        [7:0]    _zz_dataOut_payload_0_668;
  reg        [7:0]    _zz_dataOut_payload_0_669;
  reg        [7:0]    _zz_dataOut_payload_0_670;
  reg        [7:0]    _zz_dataOut_payload_0_671;
  wire                _zz_dataOut_payload_0_672;
  wire       [7:0]    _zz_dataOut_payload_0_673;
  wire       [7:0]    _zz_dataOut_payload_0_674;
  wire                _zz_dataOut_payload_0_675;
  wire       [7:0]    _zz_dataOut_payload_0_676;
  wire       [7:0]    _zz_dataOut_payload_0_677;
  wire                _zz_dataOut_payload_0_678;
  wire                _zz_dataOut_payload_0_679;
  reg        [7:0]    _zz_dataOut_payload_0_680;
  reg        [7:0]    _zz_dataOut_payload_0_681;
  reg        [7:0]    _zz_dataOut_payload_0_682;
  reg        [7:0]    _zz_dataOut_payload_0_683;
  wire                _zz_dataOut_payload_0_684;
  wire       [7:0]    _zz_dataOut_payload_0_685;
  wire       [7:0]    _zz_dataOut_payload_0_686;
  wire                _zz_dataOut_payload_0_687;
  wire       [7:0]    _zz_dataOut_payload_0_688;
  wire       [7:0]    _zz_dataOut_payload_0_689;
  wire                _zz_dataOut_payload_0_690;
  wire                _zz_dataOut_payload_0_691;
  reg        [7:0]    _zz_dataOut_payload_0_692;
  reg        [7:0]    _zz_dataOut_payload_0_693;
  reg        [7:0]    _zz_dataOut_payload_0_694;
  reg        [7:0]    _zz_dataOut_payload_0_695;
  wire                _zz_dataOut_payload_0_696;
  wire       [7:0]    _zz_dataOut_payload_0_697;
  wire       [7:0]    _zz_dataOut_payload_0_698;
  wire                _zz_dataOut_payload_0_699;
  wire       [7:0]    _zz_dataOut_payload_0_700;
  wire       [7:0]    _zz_dataOut_payload_0_701;
  wire                _zz_dataOut_payload_0_702;
  wire                _zz_dataOut_payload_0_703;
  reg        [7:0]    _zz_dataOut_payload_0_704;
  reg        [7:0]    _zz_dataOut_payload_0_705;
  reg        [7:0]    _zz_dataOut_payload_0_706;
  reg        [7:0]    _zz_dataOut_payload_0_707;
  wire                _zz_dataOut_payload_0_708;
  wire       [7:0]    _zz_dataOut_payload_0_709;
  wire       [7:0]    _zz_dataOut_payload_0_710;
  wire                _zz_dataOut_payload_0_711;
  wire       [7:0]    _zz_dataOut_payload_0_712;
  wire       [7:0]    _zz_dataOut_payload_0_713;
  wire                _zz_dataOut_payload_0_714;
  wire                _zz_dataOut_payload_0_715;
  reg        [7:0]    _zz_dataOut_payload_0_716;
  reg        [7:0]    _zz_dataOut_payload_0_717;
  reg        [7:0]    _zz_dataOut_payload_0_718;
  reg        [7:0]    _zz_dataOut_payload_0_719;
  wire                _zz_dataOut_payload_0_720;
  wire       [7:0]    _zz_dataOut_payload_0_721;
  wire       [7:0]    _zz_dataOut_payload_0_722;
  wire                _zz_dataOut_payload_0_723;
  wire       [7:0]    _zz_dataOut_payload_0_724;
  wire       [7:0]    _zz_dataOut_payload_0_725;
  wire                _zz_dataOut_payload_0_726;
  wire                _zz_dataOut_payload_0_727;
  reg        [7:0]    _zz_dataOut_payload_0_728;
  reg        [7:0]    _zz_dataOut_payload_0_729;
  reg        [7:0]    _zz_dataOut_payload_0_730;
  reg        [7:0]    _zz_dataOut_payload_0_731;
  wire                _zz_dataOut_payload_0_732;
  wire       [7:0]    _zz_dataOut_payload_0_733;
  wire       [7:0]    _zz_dataOut_payload_0_734;
  wire                _zz_dataOut_payload_0_735;
  wire       [7:0]    _zz_dataOut_payload_0_736;
  wire       [7:0]    _zz_dataOut_payload_0_737;
  wire                _zz_dataOut_payload_0_738;
  wire                _zz_dataOut_payload_0_739;
  reg        [7:0]    _zz_dataOut_payload_0_740;
  reg        [7:0]    _zz_dataOut_payload_0_741;
  reg        [7:0]    _zz_dataOut_payload_0_742;
  reg        [7:0]    _zz_dataOut_payload_0_743;
  wire                _zz_dataOut_payload_0_744;
  wire       [7:0]    _zz_dataOut_payload_0_745;
  wire       [7:0]    _zz_dataOut_payload_0_746;
  wire                _zz_dataOut_payload_0_747;
  wire       [7:0]    _zz_dataOut_payload_0_748;
  wire       [7:0]    _zz_dataOut_payload_0_749;
  wire                _zz_dataOut_payload_0_750;
  wire                _zz_dataOut_payload_0_751;
  reg        [7:0]    _zz_dataOut_payload_0_752;
  reg        [7:0]    _zz_dataOut_payload_0_753;
  reg        [7:0]    _zz_dataOut_payload_0_754;
  reg        [7:0]    _zz_dataOut_payload_0_755;
  wire                _zz_dataOut_payload_0_756;
  wire       [7:0]    _zz_dataOut_payload_0_757;
  wire       [7:0]    _zz_dataOut_payload_0_758;
  wire                _zz_dataOut_payload_0_759;
  wire       [7:0]    _zz_dataOut_payload_0_760;
  wire       [7:0]    _zz_dataOut_payload_0_761;
  wire                _zz_dataOut_payload_0_762;
  wire                _zz_dataOut_payload_0_763;
  reg        [7:0]    _zz_dataOut_payload_0_764;
  reg        [7:0]    _zz_dataOut_payload_0_765;
  reg        [7:0]    _zz_dataOut_payload_0_766;
  reg        [7:0]    _zz_dataOut_payload_0_767;
  wire                _zz_dataOut_payload_0_768;
  wire       [7:0]    _zz_dataOut_payload_0_769;
  wire       [7:0]    _zz_dataOut_payload_0_770;
  wire                _zz_dataOut_payload_0_771;
  wire       [7:0]    _zz_dataOut_payload_0_772;
  wire       [7:0]    _zz_dataOut_payload_0_773;
  wire                _zz_dataOut_payload_0_774;
  wire                _zz_dataOut_payload_0_775;
  reg        [7:0]    _zz_dataOut_payload_0_776;
  reg        [7:0]    _zz_dataOut_payload_0_777;
  reg        [7:0]    _zz_dataOut_payload_0_778;
  reg        [7:0]    _zz_dataOut_payload_0_779;
  wire                _zz_dataOut_payload_0_780;
  wire       [7:0]    _zz_dataOut_payload_0_781;
  wire       [7:0]    _zz_dataOut_payload_0_782;
  wire                _zz_dataOut_payload_0_783;
  wire       [7:0]    _zz_dataOut_payload_0_784;
  wire       [7:0]    _zz_dataOut_payload_0_785;
  wire                _zz_dataOut_payload_0_786;
  wire                _zz_dataOut_payload_0_787;
  reg        [7:0]    _zz_dataOut_payload_0_788;
  reg        [7:0]    _zz_dataOut_payload_0_789;
  reg        [7:0]    _zz_dataOut_payload_0_790;
  reg        [7:0]    _zz_dataOut_payload_0_791;
  wire                _zz_dataOut_payload_0_792;
  wire       [7:0]    _zz_dataOut_payload_0_793;
  wire       [7:0]    _zz_dataOut_payload_0_794;
  wire                _zz_dataOut_payload_0_795;
  wire       [7:0]    _zz_dataOut_payload_0_796;
  wire       [7:0]    _zz_dataOut_payload_0_797;
  wire                _zz_dataOut_payload_0_798;
  wire                _zz_dataOut_payload_0_799;
  reg        [7:0]    _zz_dataOut_payload_0_800;
  reg        [7:0]    _zz_dataOut_payload_0_801;
  reg        [7:0]    _zz_dataOut_payload_0_802;
  reg        [7:0]    _zz_dataOut_payload_0_803;
  wire                _zz_dataOut_payload_0_804;
  wire       [7:0]    _zz_dataOut_payload_0_805;
  wire       [7:0]    _zz_dataOut_payload_0_806;
  wire                _zz_dataOut_payload_0_807;
  wire       [7:0]    _zz_dataOut_payload_0_808;
  wire       [7:0]    _zz_dataOut_payload_0_809;
  wire                _zz_dataOut_payload_0_810;
  wire                _zz_dataOut_payload_0_811;
  reg        [7:0]    _zz_dataOut_payload_0_812;
  reg        [7:0]    _zz_dataOut_payload_0_813;
  reg        [7:0]    _zz_dataOut_payload_0_814;
  reg        [7:0]    _zz_dataOut_payload_0_815;
  wire                _zz_dataOut_payload_0_816;
  wire       [7:0]    _zz_dataOut_payload_0_817;
  wire       [7:0]    _zz_dataOut_payload_0_818;
  wire                _zz_dataOut_payload_0_819;
  wire       [7:0]    _zz_dataOut_payload_0_820;
  wire       [7:0]    _zz_dataOut_payload_0_821;
  wire                _zz_dataOut_payload_0_822;
  wire                _zz_dataOut_payload_0_823;
  reg        [7:0]    _zz_dataOut_payload_0_824;
  reg        [7:0]    _zz_dataOut_payload_0_825;
  reg        [7:0]    _zz_dataOut_payload_0_826;
  reg        [7:0]    _zz_dataOut_payload_0_827;
  wire                _zz_dataOut_payload_0_828;
  wire       [7:0]    _zz_dataOut_payload_0_829;
  wire       [7:0]    _zz_dataOut_payload_0_830;
  wire                _zz_dataOut_payload_0_831;
  wire       [7:0]    _zz_dataOut_payload_0_832;
  wire       [7:0]    _zz_dataOut_payload_0_833;
  wire                _zz_dataOut_payload_0_834;
  wire                _zz_dataOut_payload_0_835;
  reg        [7:0]    _zz_dataOut_payload_0_836;
  reg        [7:0]    _zz_dataOut_payload_0_837;
  reg        [7:0]    _zz_dataOut_payload_0_838;
  reg        [7:0]    _zz_dataOut_payload_0_839;
  wire                _zz_dataOut_payload_0_840;
  wire       [7:0]    _zz_dataOut_payload_0_841;
  wire       [7:0]    _zz_dataOut_payload_0_842;
  wire                _zz_dataOut_payload_0_843;
  wire       [7:0]    _zz_dataOut_payload_0_844;
  wire       [7:0]    _zz_dataOut_payload_0_845;
  wire                _zz_dataOut_payload_0_846;
  wire                _zz_dataOut_payload_0_847;
  reg        [7:0]    _zz_dataOut_payload_0_848;
  reg        [7:0]    _zz_dataOut_payload_0_849;
  reg        [7:0]    _zz_dataOut_payload_0_850;
  reg        [7:0]    _zz_dataOut_payload_0_851;
  wire                _zz_dataOut_payload_0_852;
  wire       [7:0]    _zz_dataOut_payload_0_853;
  wire       [7:0]    _zz_dataOut_payload_0_854;
  wire                _zz_dataOut_payload_0_855;
  wire       [7:0]    _zz_dataOut_payload_0_856;
  wire       [7:0]    _zz_dataOut_payload_0_857;
  wire                _zz_dataOut_payload_0_858;
  wire                _zz_dataOut_payload_0_859;
  reg        [7:0]    _zz_dataOut_payload_0_860;
  reg        [7:0]    _zz_dataOut_payload_0_861;
  reg        [7:0]    _zz_dataOut_payload_0_862;
  reg        [7:0]    _zz_dataOut_payload_0_863;
  wire                _zz_dataOut_payload_0_864;
  wire       [7:0]    _zz_dataOut_payload_0_865;
  wire       [7:0]    _zz_dataOut_payload_0_866;
  wire                _zz_dataOut_payload_0_867;
  wire       [7:0]    _zz_dataOut_payload_0_868;
  wire       [7:0]    _zz_dataOut_payload_0_869;
  wire                _zz_dataOut_payload_0_870;
  wire                _zz_dataOut_payload_0_871;
  reg        [7:0]    _zz_dataOut_payload_0_872;
  reg        [7:0]    _zz_dataOut_payload_0_873;
  reg        [7:0]    _zz_dataOut_payload_0_874;
  reg        [7:0]    _zz_dataOut_payload_0_875;
  wire                _zz_dataOut_payload_0_876;
  wire       [7:0]    _zz_dataOut_payload_0_877;
  wire       [7:0]    _zz_dataOut_payload_0_878;
  wire                _zz_dataOut_payload_0_879;
  wire       [7:0]    _zz_dataOut_payload_0_880;
  wire       [7:0]    _zz_dataOut_payload_0_881;
  wire                _zz_dataOut_payload_0_882;
  wire                _zz_dataOut_payload_0_883;
  reg        [7:0]    _zz_dataOut_payload_0_884;
  reg        [7:0]    _zz_dataOut_payload_0_885;
  reg        [7:0]    _zz_dataOut_payload_0_886;
  reg        [7:0]    _zz_dataOut_payload_0_887;
  wire                _zz_dataOut_payload_0_888;
  wire       [7:0]    _zz_dataOut_payload_0_889;
  wire       [7:0]    _zz_dataOut_payload_0_890;
  wire                _zz_dataOut_payload_0_891;
  wire       [7:0]    _zz_dataOut_payload_0_892;
  wire       [7:0]    _zz_dataOut_payload_0_893;
  wire                _zz_dataOut_payload_0_894;
  wire                _zz_dataOut_payload_0_895;
  reg        [7:0]    _zz_dataOut_payload_0_896;
  reg        [7:0]    _zz_dataOut_payload_0_897;
  reg        [7:0]    _zz_dataOut_payload_0_898;
  reg        [7:0]    _zz_dataOut_payload_0_899;
  wire                _zz_dataOut_payload_0_900;
  wire       [7:0]    _zz_dataOut_payload_0_901;
  wire       [7:0]    _zz_dataOut_payload_0_902;
  wire                _zz_dataOut_payload_0_903;
  wire       [7:0]    _zz_dataOut_payload_0_904;
  wire       [7:0]    _zz_dataOut_payload_0_905;
  wire                _zz_dataOut_payload_0_906;
  wire                _zz_dataOut_payload_0_907;
  reg        [7:0]    _zz_dataOut_payload_0_908;
  reg        [7:0]    _zz_dataOut_payload_0_909;
  reg        [7:0]    _zz_dataOut_payload_0_910;
  reg        [7:0]    _zz_dataOut_payload_0_911;
  wire                _zz_dataOut_payload_0_912;
  wire       [7:0]    _zz_dataOut_payload_0_913;
  wire       [7:0]    _zz_dataOut_payload_0_914;
  wire                _zz_dataOut_payload_0_915;
  wire       [7:0]    _zz_dataOut_payload_0_916;
  wire       [7:0]    _zz_dataOut_payload_0_917;
  wire                _zz_dataOut_payload_0_918;
  wire                _zz_dataOut_payload_0_919;
  reg        [7:0]    _zz_dataOut_payload_0_920;
  reg        [7:0]    _zz_dataOut_payload_0_921;
  reg        [7:0]    _zz_dataOut_payload_0_922;
  reg        [7:0]    _zz_dataOut_payload_0_923;
  wire                _zz_dataOut_payload_0_924;
  wire       [7:0]    _zz_dataOut_payload_0_925;
  wire       [7:0]    _zz_dataOut_payload_0_926;
  wire                _zz_dataOut_payload_0_927;
  wire       [7:0]    _zz_dataOut_payload_0_928;
  wire       [7:0]    _zz_dataOut_payload_0_929;
  wire                _zz_dataOut_payload_0_930;
  wire                _zz_dataOut_payload_0_931;
  reg        [7:0]    _zz_dataOut_payload_0_932;
  reg        [7:0]    _zz_dataOut_payload_0_933;
  reg        [7:0]    _zz_dataOut_payload_0_934;
  reg        [7:0]    _zz_dataOut_payload_0_935;
  wire                _zz_dataOut_payload_0_936;
  wire       [7:0]    _zz_dataOut_payload_0_937;
  wire       [7:0]    _zz_dataOut_payload_0_938;
  wire                _zz_dataOut_payload_0_939;
  wire       [7:0]    _zz_dataOut_payload_0_940;
  wire       [7:0]    _zz_dataOut_payload_0_941;
  wire                _zz_dataOut_payload_0_942;
  wire                _zz_dataOut_payload_0_943;
  reg        [7:0]    _zz_dataOut_payload_0_944;
  reg        [7:0]    _zz_dataOut_payload_0_945;
  reg        [7:0]    _zz_dataOut_payload_0_946;
  reg        [7:0]    _zz_dataOut_payload_0_947;
  wire                _zz_dataOut_payload_0_948;
  wire       [7:0]    _zz_dataOut_payload_0_949;
  wire       [7:0]    _zz_dataOut_payload_0_950;
  wire                _zz_dataOut_payload_0_951;
  wire       [7:0]    _zz_dataOut_payload_0_952;
  wire       [7:0]    _zz_dataOut_payload_0_953;
  wire                _zz_dataOut_payload_0_954;
  wire                _zz_dataOut_payload_0_955;
  reg        [7:0]    _zz_dataOut_payload_0_956;
  reg        [7:0]    _zz_dataOut_payload_0_957;
  reg        [7:0]    _zz_dataOut_payload_0_958;
  reg        [7:0]    _zz_dataOut_payload_0_959;
  wire                _zz_dataOut_payload_0_960;
  wire       [7:0]    _zz_dataOut_payload_0_961;
  wire       [7:0]    _zz_dataOut_payload_0_962;
  wire                _zz_dataOut_payload_0_963;
  wire       [7:0]    _zz_dataOut_payload_0_964;
  wire       [7:0]    _zz_dataOut_payload_0_965;
  wire                _zz_dataOut_payload_0_966;
  wire                _zz_dataOut_payload_0_967;
  reg        [7:0]    _zz_dataOut_payload_0_968;
  reg        [7:0]    _zz_dataOut_payload_0_969;
  reg        [7:0]    _zz_dataOut_payload_0_970;
  reg        [7:0]    _zz_dataOut_payload_0_971;
  wire                _zz_dataOut_payload_0_972;
  wire       [7:0]    _zz_dataOut_payload_0_973;
  wire       [7:0]    _zz_dataOut_payload_0_974;
  wire                _zz_dataOut_payload_0_975;
  wire       [7:0]    _zz_dataOut_payload_0_976;
  wire       [7:0]    _zz_dataOut_payload_0_977;
  wire                _zz_dataOut_payload_0_978;
  wire                _zz_dataOut_payload_0_979;
  reg        [7:0]    _zz_dataOut_payload_0_980;
  reg        [7:0]    _zz_dataOut_payload_0_981;
  reg        [7:0]    _zz_dataOut_payload_0_982;
  reg        [7:0]    _zz_dataOut_payload_0_983;
  wire                _zz_dataOut_payload_0_984;
  wire       [7:0]    _zz_dataOut_payload_0_985;
  wire       [7:0]    _zz_dataOut_payload_0_986;
  wire                _zz_dataOut_payload_0_987;
  wire       [7:0]    _zz_dataOut_payload_0_988;
  wire       [7:0]    _zz_dataOut_payload_0_989;
  wire                _zz_dataOut_payload_0_990;
  wire                _zz_dataOut_payload_0_991;
  reg        [7:0]    _zz_dataOut_payload_0_992;
  reg        [7:0]    _zz_dataOut_payload_0_993;
  reg        [7:0]    _zz_dataOut_payload_0_994;
  reg        [7:0]    _zz_dataOut_payload_0_995;
  wire                _zz_dataOut_payload_0_996;
  wire       [7:0]    _zz_dataOut_payload_0_997;
  wire       [7:0]    _zz_dataOut_payload_0_998;
  wire                _zz_dataOut_payload_0_999;
  wire       [7:0]    _zz_dataOut_payload_0_1000;
  wire       [7:0]    _zz_dataOut_payload_0_1001;
  wire                _zz_dataOut_payload_0_1002;
  wire                _zz_dataOut_payload_0_1003;
  reg        [7:0]    _zz_dataOut_payload_0_1004;
  reg        [7:0]    _zz_dataOut_payload_0_1005;
  reg        [7:0]    _zz_dataOut_payload_0_1006;
  reg        [7:0]    _zz_dataOut_payload_0_1007;
  wire                _zz_dataOut_payload_0_1008;
  wire       [7:0]    _zz_dataOut_payload_0_1009;
  wire       [7:0]    _zz_dataOut_payload_0_1010;
  wire                _zz_dataOut_payload_0_1011;
  wire       [7:0]    _zz_dataOut_payload_0_1012;
  wire       [7:0]    _zz_dataOut_payload_0_1013;
  wire                _zz_dataOut_payload_0_1014;
  wire                _zz_dataOut_payload_0_1015;
  reg        [7:0]    _zz_dataOut_payload_0_1016;
  reg        [7:0]    _zz_dataOut_payload_0_1017;
  reg        [7:0]    _zz_dataOut_payload_0_1018;
  reg        [7:0]    _zz_dataOut_payload_0_1019;
  wire                _zz_dataOut_payload_0_1020;
  wire       [7:0]    _zz_dataOut_payload_0_1021;
  wire       [7:0]    _zz_dataOut_payload_0_1022;
  wire                _zz_dataOut_payload_0_1023;
  wire       [7:0]    _zz_dataOut_payload_0_1024;
  wire       [7:0]    _zz_dataOut_payload_0_1025;
  wire                _zz_dataOut_payload_0_1026;
  wire                _zz_dataOut_payload_0_1027;
  reg        [7:0]    _zz_dataOut_payload_0_1028;
  reg        [7:0]    _zz_dataOut_payload_0_1029;
  reg        [7:0]    _zz_dataOut_payload_0_1030;
  reg        [7:0]    _zz_dataOut_payload_0_1031;
  wire                _zz_dataOut_payload_0_1032;
  wire       [7:0]    _zz_dataOut_payload_0_1033;
  wire       [7:0]    _zz_dataOut_payload_0_1034;
  wire                _zz_dataOut_payload_0_1035;
  wire       [7:0]    _zz_dataOut_payload_0_1036;
  wire       [7:0]    _zz_dataOut_payload_0_1037;
  wire                _zz_dataOut_payload_0_1038;
  wire                _zz_dataOut_payload_0_1039;
  reg        [7:0]    _zz_dataOut_payload_0_1040;
  reg        [7:0]    _zz_dataOut_payload_0_1041;
  reg        [7:0]    _zz_dataOut_payload_0_1042;
  reg        [7:0]    _zz_dataOut_payload_0_1043;
  wire                _zz_dataOut_payload_0_1044;
  wire       [7:0]    _zz_dataOut_payload_0_1045;
  wire       [7:0]    _zz_dataOut_payload_0_1046;
  wire                _zz_dataOut_payload_0_1047;
  wire       [7:0]    _zz_dataOut_payload_0_1048;
  wire       [7:0]    _zz_dataOut_payload_0_1049;
  wire                _zz_dataOut_payload_0_1050;
  wire                _zz_dataOut_payload_0_1051;
  reg        [7:0]    _zz_dataOut_payload_0_1052;
  reg        [7:0]    _zz_dataOut_payload_0_1053;
  reg        [7:0]    _zz_dataOut_payload_0_1054;
  reg        [7:0]    _zz_dataOut_payload_0_1055;
  wire                _zz_dataOut_payload_0_1056;
  wire       [7:0]    _zz_dataOut_payload_0_1057;
  wire       [7:0]    _zz_dataOut_payload_0_1058;
  wire                _zz_dataOut_payload_0_1059;
  wire       [7:0]    _zz_dataOut_payload_0_1060;
  wire       [7:0]    _zz_dataOut_payload_0_1061;
  wire                _zz_dataOut_payload_0_1062;
  wire                _zz_dataOut_payload_0_1063;
  reg        [7:0]    _zz_dataOut_payload_0_1064;
  reg        [7:0]    _zz_dataOut_payload_0_1065;
  reg        [7:0]    _zz_dataOut_payload_0_1066;
  reg        [7:0]    _zz_dataOut_payload_0_1067;
  wire                _zz_dataOut_payload_0_1068;
  wire       [7:0]    _zz_dataOut_payload_0_1069;
  wire       [7:0]    _zz_dataOut_payload_0_1070;
  wire                _zz_dataOut_payload_0_1071;
  wire       [7:0]    _zz_dataOut_payload_0_1072;
  wire       [7:0]    _zz_dataOut_payload_0_1073;
  wire                _zz_dataOut_payload_0_1074;
  wire                _zz_dataOut_payload_0_1075;
  reg        [7:0]    _zz_dataOut_payload_0_1076;
  reg        [7:0]    _zz_dataOut_payload_0_1077;
  reg        [7:0]    _zz_dataOut_payload_0_1078;
  reg        [7:0]    _zz_dataOut_payload_0_1079;
  wire                _zz_dataOut_payload_0_1080;
  wire       [7:0]    _zz_dataOut_payload_0_1081;
  wire       [7:0]    _zz_dataOut_payload_0_1082;
  wire                _zz_dataOut_payload_0_1083;
  wire       [7:0]    _zz_dataOut_payload_0_1084;
  wire       [7:0]    _zz_dataOut_payload_0_1085;
  wire                _zz_dataOut_payload_0_1086;
  wire                _zz_dataOut_payload_0_1087;
  reg        [7:0]    _zz_dataOut_payload_0_1088;
  reg        [7:0]    _zz_dataOut_payload_0_1089;
  reg        [7:0]    _zz_dataOut_payload_0_1090;
  reg        [7:0]    _zz_dataOut_payload_0_1091;
  wire                _zz_dataOut_payload_0_1092;
  wire       [7:0]    _zz_dataOut_payload_0_1093;
  wire       [7:0]    _zz_dataOut_payload_0_1094;
  wire                _zz_dataOut_payload_0_1095;
  wire       [7:0]    _zz_dataOut_payload_0_1096;
  wire       [7:0]    _zz_dataOut_payload_0_1097;
  wire                _zz_dataOut_payload_0_1098;
  wire                _zz_dataOut_payload_0_1099;
  reg        [7:0]    _zz_dataOut_payload_0_1100;
  reg        [7:0]    _zz_dataOut_payload_0_1101;
  reg        [7:0]    _zz_dataOut_payload_0_1102;
  reg        [7:0]    _zz_dataOut_payload_0_1103;
  wire                _zz_dataOut_payload_0_1104;
  wire       [7:0]    _zz_dataOut_payload_0_1105;
  wire       [7:0]    _zz_dataOut_payload_0_1106;
  wire                _zz_dataOut_payload_0_1107;
  wire       [7:0]    _zz_dataOut_payload_0_1108;
  wire       [7:0]    _zz_dataOut_payload_0_1109;
  wire                _zz_dataOut_payload_0_1110;
  wire                _zz_dataOut_payload_0_1111;
  reg        [7:0]    _zz_dataOut_payload_0_1112;
  reg        [7:0]    _zz_dataOut_payload_0_1113;
  reg        [7:0]    _zz_dataOut_payload_0_1114;
  reg        [7:0]    _zz_dataOut_payload_0_1115;
  wire                _zz_dataOut_payload_0_1116;
  wire       [7:0]    _zz_dataOut_payload_0_1117;
  wire       [7:0]    _zz_dataOut_payload_0_1118;
  wire                _zz_dataOut_payload_0_1119;
  wire       [7:0]    _zz_dataOut_payload_0_1120;
  wire       [7:0]    _zz_dataOut_payload_0_1121;
  wire                _zz_dataOut_payload_0_1122;
  wire                _zz_dataOut_payload_0_1123;
  reg        [7:0]    _zz_dataOut_payload_0_1124;
  reg        [7:0]    _zz_dataOut_payload_0_1125;
  reg        [7:0]    _zz_dataOut_payload_0_1126;
  reg        [7:0]    _zz_dataOut_payload_0_1127;
  wire                _zz_dataOut_payload_0_1128;
  wire       [7:0]    _zz_dataOut_payload_0_1129;
  wire       [7:0]    _zz_dataOut_payload_0_1130;
  wire                _zz_dataOut_payload_0_1131;
  wire       [7:0]    _zz_dataOut_payload_0_1132;
  wire       [7:0]    _zz_dataOut_payload_0_1133;
  wire                _zz_dataOut_payload_0_1134;
  wire                _zz_dataOut_payload_0_1135;
  reg        [7:0]    _zz_dataOut_payload_0_1136;
  reg        [7:0]    _zz_dataOut_payload_0_1137;
  reg        [7:0]    _zz_dataOut_payload_0_1138;
  reg        [7:0]    _zz_dataOut_payload_0_1139;
  wire                _zz_dataOut_payload_0_1140;
  wire       [7:0]    _zz_dataOut_payload_0_1141;
  wire       [7:0]    _zz_dataOut_payload_0_1142;
  wire                _zz_dataOut_payload_0_1143;
  wire       [7:0]    _zz_dataOut_payload_0_1144;
  wire       [7:0]    _zz_dataOut_payload_0_1145;
  wire                _zz_dataOut_payload_0_1146;
  wire                _zz_dataOut_payload_0_1147;
  reg        [7:0]    _zz_dataOut_payload_0_1148;
  reg        [7:0]    _zz_dataOut_payload_0_1149;
  reg        [7:0]    _zz_dataOut_payload_0_1150;
  reg        [7:0]    _zz_dataOut_payload_0_1151;
  reg        [7:0]    _zz_dataOut_payload_0_1152;
  reg        [7:0]    _zz_dataOut_payload_0_1153;
  reg        [7:0]    _zz_dataOut_payload_0_1154;
  reg        [7:0]    _zz_dataOut_payload_0_1155;
  reg        [7:0]    _zz_dataOut_payload_0_1156;
  reg        [7:0]    _zz_dataOut_payload_0_1157;
  reg        [7:0]    _zz_dataOut_payload_0_1158;
  reg        [7:0]    _zz_dataOut_payload_0_1159;
  reg        [7:0]    _zz_dataOut_payload_0_1160;
  reg        [7:0]    _zz_dataOut_payload_0_1161;
  reg        [7:0]    _zz_dataOut_payload_0_1162;
  reg        [7:0]    _zz_dataOut_payload_0_1163;
  reg        [7:0]    _zz_dataOut_payload_0_1164;
  reg        [7:0]    _zz_dataOut_payload_0_1165;
  reg        [7:0]    _zz_dataOut_payload_0_1166;
  reg        [7:0]    _zz_dataOut_payload_0_1167;
  reg        [7:0]    _zz_dataOut_payload_0_1168;
  reg        [7:0]    _zz_dataOut_payload_0_1169;
  reg        [7:0]    _zz_dataOut_payload_0_1170;
  reg        [7:0]    _zz_dataOut_payload_0_1171;
  reg        [7:0]    _zz_dataOut_payload_0_1172;
  reg        [7:0]    _zz_dataOut_payload_0_1173;
  reg        [7:0]    _zz_dataOut_payload_0_1174;
  reg        [7:0]    _zz_dataOut_payload_0_1175;
  reg        [7:0]    _zz_dataOut_payload_0_1176;
  reg        [7:0]    _zz_dataOut_payload_0_1177;
  reg        [7:0]    _zz_dataOut_payload_0_1178;
  reg        [7:0]    _zz_dataOut_payload_0_1179;
  reg        [7:0]    _zz_dataOut_payload_0_1180;
  reg        [7:0]    _zz_dataOut_payload_0_1181;
  reg        [7:0]    _zz_dataOut_payload_0_1182;
  reg        [7:0]    _zz_dataOut_payload_0_1183;
  reg        [7:0]    _zz_dataOut_payload_0_1184;
  reg        [7:0]    _zz_dataOut_payload_0_1185;
  reg        [7:0]    _zz_dataOut_payload_0_1186;
  reg        [7:0]    _zz_dataOut_payload_0_1187;
  reg        [7:0]    _zz_dataOut_payload_0_1188;
  reg        [7:0]    _zz_dataOut_payload_0_1189;
  reg        [7:0]    _zz_dataOut_payload_0_1190;
  reg        [7:0]    _zz_dataOut_payload_0_1191;
  reg        [7:0]    _zz_dataOut_payload_0_1192;
  reg        [7:0]    _zz_dataOut_payload_0_1193;
  reg        [7:0]    _zz_dataOut_payload_0_1194;
  reg        [7:0]    _zz_dataOut_payload_0_1195;
  reg        [7:0]    _zz_dataOut_payload_0_1196;
  reg        [7:0]    _zz_dataOut_payload_0_1197;
  reg        [7:0]    _zz_dataOut_payload_0_1198;
  reg        [7:0]    _zz_dataOut_payload_0_1199;
  reg        [7:0]    _zz_dataOut_payload_0_1200;
  reg        [7:0]    _zz_dataOut_payload_0_1201;
  reg        [7:0]    _zz_dataOut_payload_0_1202;
  reg        [7:0]    _zz_dataOut_payload_0_1203;
  reg        [7:0]    _zz_dataOut_payload_0_1204;
  reg        [7:0]    _zz_dataOut_payload_0_1205;
  reg        [7:0]    _zz_dataOut_payload_0_1206;
  reg        [7:0]    _zz_dataOut_payload_0_1207;
  reg        [7:0]    _zz_dataOut_payload_0_1208;
  reg        [7:0]    _zz_dataOut_payload_0_1209;
  reg        [7:0]    _zz_dataOut_payload_0_1210;
  reg        [7:0]    _zz_dataOut_payload_0_1211;
  reg        [7:0]    _zz_dataOut_payload_0_1212;
  reg        [7:0]    _zz_dataOut_payload_0_1213;
  reg        [7:0]    _zz_dataOut_payload_0_1214;
  reg        [7:0]    _zz_dataOut_payload_0_1215;
  reg        [7:0]    _zz_dataOut_payload_0_1216;
  reg        [7:0]    _zz_dataOut_payload_0_1217;
  reg        [7:0]    _zz_dataOut_payload_0_1218;
  reg        [7:0]    _zz_dataOut_payload_0_1219;
  reg        [7:0]    _zz_dataOut_payload_0_1220;
  reg        [7:0]    _zz_dataOut_payload_0_1221;
  reg        [7:0]    _zz_dataOut_payload_0_1222;
  reg        [7:0]    _zz_dataOut_payload_0_1223;
  reg        [7:0]    _zz_dataOut_payload_0_1224;
  reg        [7:0]    _zz_dataOut_payload_0_1225;
  reg        [7:0]    _zz_dataOut_payload_0_1226;
  reg        [7:0]    _zz_dataOut_payload_0_1227;
  reg        [7:0]    _zz_dataOut_payload_0_1228;
  reg        [7:0]    _zz_dataOut_payload_0_1229;
  reg        [7:0]    _zz_dataOut_payload_0_1230;
  reg        [7:0]    _zz_dataOut_payload_0_1231;
  reg        [7:0]    _zz_dataOut_payload_0_1232;
  reg        [7:0]    _zz_dataOut_payload_0_1233;
  reg        [7:0]    _zz_dataOut_payload_0_1234;
  reg        [7:0]    _zz_dataOut_payload_0_1235;
  reg        [7:0]    _zz_dataOut_payload_0_1236;
  reg        [7:0]    _zz_dataOut_payload_0_1237;
  reg        [7:0]    _zz_dataOut_payload_0_1238;
  reg        [7:0]    _zz_dataOut_payload_0_1239;
  reg        [7:0]    _zz_dataOut_payload_0_1240;
  reg        [7:0]    _zz_dataOut_payload_0_1241;
  reg        [7:0]    _zz_dataOut_payload_0_1242;
  reg        [7:0]    _zz_dataOut_payload_0_1243;
  reg        [7:0]    _zz_dataOut_payload_0_1244;
  reg        [7:0]    _zz_dataOut_payload_0_1245;
  reg        [7:0]    _zz_dataOut_payload_0_1246;
  reg        [7:0]    _zz_dataOut_payload_0_1247;
  reg        [7:0]    _zz_dataOut_payload_0_1248;
  reg        [7:0]    _zz_dataOut_payload_0_1249;
  reg        [7:0]    _zz_dataOut_payload_0_1250;
  reg        [7:0]    _zz_dataOut_payload_0_1251;
  reg        [7:0]    _zz_dataOut_payload_0_1252;
  reg        [7:0]    _zz_dataOut_payload_0_1253;
  reg        [7:0]    _zz_dataOut_payload_0_1254;
  reg        [7:0]    _zz_dataOut_payload_0_1255;
  reg        [7:0]    _zz_dataOut_payload_0_1256;
  reg        [7:0]    _zz_dataOut_payload_0_1257;
  reg        [7:0]    _zz_dataOut_payload_0_1258;
  reg        [7:0]    _zz_dataOut_payload_0_1259;
  reg        [7:0]    _zz_dataOut_payload_0_1260;
  reg        [7:0]    _zz_dataOut_payload_0_1261;
  reg        [7:0]    _zz_dataOut_payload_0_1262;
  reg        [7:0]    _zz_dataOut_payload_0_1263;
  reg        [7:0]    _zz_dataOut_payload_0_1264;
  reg        [7:0]    _zz_dataOut_payload_0_1265;
  reg        [7:0]    _zz_dataOut_payload_0_1266;
  reg        [7:0]    _zz_dataOut_payload_0_1267;
  reg        [7:0]    _zz_dataOut_payload_0_1268;
  reg        [7:0]    _zz_dataOut_payload_0_1269;
  reg        [7:0]    _zz_dataOut_payload_0_1270;
  reg        [7:0]    _zz_dataOut_payload_0_1271;
  reg        [7:0]    _zz_dataOut_payload_0_1272;
  reg        [7:0]    _zz_dataOut_payload_0_1273;
  reg        [7:0]    _zz_dataOut_payload_0_1274;
  reg        [7:0]    _zz_dataOut_payload_0_1275;
  reg        [7:0]    _zz_dataOut_payload_0_1276;
  reg        [7:0]    _zz_dataOut_payload_0_1277;
  reg        [7:0]    _zz_dataOut_payload_0_1278;
  reg        [7:0]    _zz_dataOut_payload_0_1279;
  reg        [7:0]    _zz_dataOut_payload_0_1280;
  reg        [7:0]    _zz_dataOut_payload_0_1281;
  reg        [7:0]    _zz_dataOut_payload_0_1282;
  reg        [7:0]    _zz_dataOut_payload_0_1283;
  reg        [7:0]    _zz_dataOut_payload_0_1284;
  reg        [7:0]    _zz_dataOut_payload_0_1285;
  reg        [7:0]    _zz_dataOut_payload_0_1286;
  reg        [7:0]    _zz_dataOut_payload_0_1287;
  reg        [7:0]    _zz_dataOut_payload_0_1288;
  reg        [7:0]    _zz_dataOut_payload_0_1289;
  reg        [7:0]    _zz_dataOut_payload_0_1290;
  reg        [7:0]    _zz_dataOut_payload_0_1291;
  reg        [7:0]    _zz_dataOut_payload_0_1292;
  reg        [7:0]    _zz_dataOut_payload_0_1293;
  reg        [7:0]    _zz_dataOut_payload_0_1294;
  reg        [7:0]    _zz_dataOut_payload_0_1295;
  reg        [7:0]    _zz_dataOut_payload_0_1296;
  reg        [7:0]    _zz_dataOut_payload_0_1297;
  reg        [7:0]    _zz_dataOut_payload_0_1298;
  reg        [7:0]    _zz_dataOut_payload_0_1299;
  reg        [7:0]    _zz_dataOut_payload_0_1300;
  reg        [7:0]    _zz_dataOut_payload_0_1301;
  reg        [7:0]    _zz_dataOut_payload_0_1302;
  reg        [7:0]    _zz_dataOut_payload_0_1303;
  reg        [7:0]    _zz_dataOut_payload_0_1304;
  reg        [7:0]    _zz_dataOut_payload_0_1305;
  reg        [7:0]    _zz_dataOut_payload_0_1306;
  reg        [7:0]    _zz_dataOut_payload_0_1307;
  reg        [7:0]    _zz_dataOut_payload_0_1308;
  reg        [7:0]    _zz_dataOut_payload_0_1309;
  reg        [7:0]    _zz_dataOut_payload_0_1310;
  reg        [7:0]    _zz_dataOut_payload_0_1311;
  reg        [7:0]    _zz_dataOut_payload_0_1312;
  reg        [7:0]    _zz_dataOut_payload_0_1313;
  reg        [7:0]    _zz_dataOut_payload_0_1314;
  reg        [7:0]    _zz_dataOut_payload_0_1315;
  reg        [7:0]    _zz_dataOut_payload_0_1316;
  reg        [7:0]    _zz_dataOut_payload_0_1317;
  reg        [7:0]    _zz_dataOut_payload_0_1318;
  reg        [7:0]    _zz_dataOut_payload_0_1319;
  reg        [7:0]    _zz_dataOut_payload_0_1320;
  reg        [7:0]    _zz_dataOut_payload_0_1321;
  reg        [7:0]    _zz_dataOut_payload_0_1322;
  reg        [7:0]    _zz_dataOut_payload_0_1323;
  reg        [7:0]    _zz_dataOut_payload_0_1324;
  reg        [7:0]    _zz_dataOut_payload_0_1325;
  reg        [7:0]    _zz_dataOut_payload_0_1326;
  reg        [7:0]    _zz_dataOut_payload_0_1327;
  reg        [7:0]    _zz_dataOut_payload_0_1328;
  reg        [7:0]    _zz_dataOut_payload_0_1329;
  reg        [7:0]    _zz_dataOut_payload_0_1330;
  reg        [7:0]    _zz_dataOut_payload_0_1331;
  reg        [7:0]    _zz_dataOut_payload_0_1332;
  reg        [7:0]    _zz_dataOut_payload_0_1333;
  reg        [7:0]    _zz_dataOut_payload_0_1334;
  reg        [7:0]    _zz_dataOut_payload_0_1335;
  reg        [7:0]    _zz_dataOut_payload_0_1336;
  reg        [7:0]    _zz_dataOut_payload_0_1337;
  reg        [7:0]    _zz_dataOut_payload_0_1338;
  reg        [7:0]    _zz_dataOut_payload_0_1339;
  reg        [7:0]    _zz_dataOut_payload_0_1340;
  reg        [7:0]    _zz_dataOut_payload_0_1341;
  reg        [7:0]    _zz_dataOut_payload_0_1342;
  reg        [7:0]    _zz_dataOut_payload_0_1343;
  reg        [7:0]    _zz_dataOut_payload_0_1344;
  reg        [7:0]    _zz_dataOut_payload_0_1345;
  reg        [7:0]    _zz_dataOut_payload_0_1346;
  reg        [7:0]    _zz_dataOut_payload_0_1347;
  reg        [7:0]    _zz_dataOut_payload_0_1348;
  reg        [7:0]    _zz_dataOut_payload_0_1349;
  reg        [7:0]    _zz_dataOut_payload_0_1350;
  reg        [7:0]    _zz_dataOut_payload_0_1351;
  reg        [7:0]    _zz_dataOut_payload_0_1352;
  reg        [7:0]    _zz_dataOut_payload_0_1353;
  reg        [7:0]    _zz_dataOut_payload_0_1354;
  reg        [7:0]    _zz_dataOut_payload_0_1355;
  reg        [7:0]    _zz_dataOut_payload_0_1356;
  reg        [7:0]    _zz_dataOut_payload_0_1357;
  reg        [7:0]    _zz_dataOut_payload_0_1358;
  reg        [7:0]    _zz_dataOut_payload_0_1359;
  reg        [7:0]    _zz_dataOut_payload_0_1360;
  reg        [7:0]    _zz_dataOut_payload_0_1361;
  reg        [7:0]    _zz_dataOut_payload_0_1362;
  reg        [7:0]    _zz_dataOut_payload_0_1363;
  reg        [7:0]    _zz_dataOut_payload_0_1364;
  reg        [7:0]    _zz_dataOut_payload_0_1365;
  reg        [7:0]    _zz_dataOut_payload_0_1366;
  reg        [7:0]    _zz_dataOut_payload_0_1367;
  reg        [7:0]    _zz_dataOut_payload_0_1368;
  reg        [7:0]    _zz_dataOut_payload_0_1369;
  reg        [7:0]    _zz_dataOut_payload_0_1370;
  reg        [7:0]    _zz_dataOut_payload_0_1371;
  reg        [7:0]    _zz_dataOut_payload_0_1372;
  reg        [7:0]    _zz_dataOut_payload_0_1373;
  reg        [7:0]    _zz_dataOut_payload_0_1374;
  reg        [7:0]    _zz_dataOut_payload_0_1375;
  reg        [7:0]    _zz_dataOut_payload_0_1376;
  reg        [7:0]    _zz_dataOut_payload_0_1377;
  reg        [7:0]    _zz_dataOut_payload_0_1378;
  reg        [7:0]    _zz_dataOut_payload_0_1379;
  reg        [7:0]    _zz_dataOut_payload_0_1380;
  reg        [7:0]    _zz_dataOut_payload_0_1381;
  reg        [7:0]    _zz_dataOut_payload_0_1382;
  reg        [7:0]    _zz_dataOut_payload_0_1383;
  reg        [7:0]    _zz_dataOut_payload_0_1384;
  reg        [7:0]    _zz_dataOut_payload_0_1385;
  reg        [7:0]    _zz_dataOut_payload_0_1386;
  reg        [7:0]    _zz_dataOut_payload_0_1387;
  reg        [7:0]    _zz_dataOut_payload_0_1388;
  reg        [7:0]    _zz_dataOut_payload_0_1389;
  reg        [7:0]    _zz_dataOut_payload_0_1390;
  reg        [7:0]    _zz_dataOut_payload_0_1391;
  reg        [7:0]    _zz_dataOut_payload_0_1392;
  reg        [7:0]    _zz_dataOut_payload_0_1393;
  reg        [7:0]    _zz_dataOut_payload_0_1394;
  reg        [7:0]    _zz_dataOut_payload_0_1395;
  reg        [7:0]    _zz_dataOut_payload_0_1396;
  reg        [7:0]    _zz_dataOut_payload_0_1397;
  reg        [7:0]    _zz_dataOut_payload_0_1398;
  reg        [7:0]    _zz_dataOut_payload_0_1399;
  reg        [7:0]    _zz_dataOut_payload_0_1400;
  reg        [7:0]    _zz_dataOut_payload_0_1401;
  reg        [7:0]    _zz_dataOut_payload_0_1402;
  reg        [7:0]    _zz_dataOut_payload_0_1403;
  reg        [7:0]    _zz_dataOut_payload_0_1404;
  reg        [7:0]    _zz_dataOut_payload_0_1405;
  reg        [7:0]    _zz_dataOut_payload_0_1406;
  reg        [7:0]    _zz_dataOut_payload_0_1407;
  wire                _zz_dataOut_payload_0_1408;
  wire       [7:0]    _zz_dataOut_payload_0_1409;
  wire       [7:0]    _zz_dataOut_payload_0_1410;
  wire                _zz_dataOut_payload_0_1411;
  wire       [7:0]    _zz_dataOut_payload_0_1412;
  wire       [7:0]    _zz_dataOut_payload_0_1413;
  wire                _zz_dataOut_payload_0_1414;
  wire       [7:0]    _zz_dataOut_payload_0_1415;
  wire       [7:0]    _zz_dataOut_payload_0_1416;
  wire                _zz_dataOut_payload_0_1417;
  wire       [7:0]    _zz_dataOut_payload_0_1418;
  wire       [7:0]    _zz_dataOut_payload_0_1419;
  wire                _zz_dataOut_payload_0_1420;
  wire       [7:0]    _zz_dataOut_payload_0_1421;
  wire       [7:0]    _zz_dataOut_payload_0_1422;
  wire                _zz_dataOut_payload_0_1423;
  wire       [7:0]    _zz_dataOut_payload_0_1424;
  wire       [7:0]    _zz_dataOut_payload_0_1425;
  wire                _zz_dataOut_payload_0_1426;
  wire                _zz_dataOut_payload_0_1427;
  reg        [7:0]    _zz_dataOut_payload_0_1428;
  reg        [7:0]    _zz_dataOut_payload_0_1429;
  reg        [7:0]    _zz_dataOut_payload_0_1430;
  reg        [7:0]    _zz_dataOut_payload_0_1431;
  wire                _zz_dataOut_payload_0_1432;
  wire       [7:0]    _zz_dataOut_payload_0_1433;
  wire       [7:0]    _zz_dataOut_payload_0_1434;
  wire                _zz_dataOut_payload_0_1435;
  wire       [7:0]    _zz_dataOut_payload_0_1436;
  wire       [7:0]    _zz_dataOut_payload_0_1437;
  wire                _zz_dataOut_payload_0_1438;
  wire                _zz_dataOut_payload_0_1439;
  reg        [7:0]    _zz_dataOut_payload_0_1440;
  reg        [7:0]    _zz_dataOut_payload_0_1441;
  reg        [7:0]    _zz_dataOut_payload_0_1442;
  reg        [7:0]    _zz_dataOut_payload_0_1443;
  reg        [7:0]    _zz_dataOut_payload_0_1444;
  reg        [7:0]    _zz_dataOut_payload_0_1445;
  reg        [7:0]    _zz_dataOut_payload_0_1446;
  reg        [7:0]    _zz_dataOut_payload_0_1447;
  reg        [7:0]    _zz_dataOut_payload_0_1448;
  reg        [7:0]    _zz_dataOut_payload_0_1449;
  reg        [7:0]    _zz_dataOut_payload_0_1450;
  reg        [7:0]    _zz_dataOut_payload_0_1451;
  wire                _zz_dataOut_payload_0_1452;
  wire       [7:0]    _zz_dataOut_payload_0_1453;
  wire       [7:0]    _zz_dataOut_payload_0_1454;
  wire                _zz_dataOut_payload_0_1455;
  wire       [7:0]    _zz_dataOut_payload_0_1456;
  wire       [7:0]    _zz_dataOut_payload_0_1457;
  wire                _zz_dataOut_payload_0_1458;
  wire       [7:0]    _zz_dataOut_payload_0_1459;
  wire       [7:0]    _zz_dataOut_payload_0_1460;
  wire                _zz_dataOut_payload_0_1461;
  wire       [7:0]    _zz_dataOut_payload_0_1462;
  wire       [7:0]    _zz_dataOut_payload_0_1463;
  wire                _zz_dataOut_payload_0_1464;
  wire       [7:0]    _zz_dataOut_payload_0_1465;
  wire       [7:0]    _zz_dataOut_payload_0_1466;
  wire                _zz_dataOut_payload_0_1467;
  wire       [7:0]    _zz_dataOut_payload_0_1468;
  wire       [7:0]    _zz_dataOut_payload_0_1469;
  wire                _zz_dataOut_payload_0_1470;
  wire                _zz_dataOut_payload_0_1471;
  reg        [7:0]    _zz_dataOut_payload_0_1472;
  reg        [7:0]    _zz_dataOut_payload_0_1473;
  reg        [7:0]    _zz_dataOut_payload_0_1474;
  reg        [7:0]    _zz_dataOut_payload_0_1475;
  wire                _zz_dataOut_payload_0_1476;
  wire       [7:0]    _zz_dataOut_payload_0_1477;
  wire       [7:0]    _zz_dataOut_payload_0_1478;
  wire                _zz_dataOut_payload_0_1479;
  wire       [7:0]    _zz_dataOut_payload_0_1480;
  wire       [7:0]    _zz_dataOut_payload_0_1481;
  wire                _zz_dataOut_payload_0_1482;
  wire                _zz_dataOut_payload_0_1483;
  reg        [7:0]    _zz_dataOut_payload_0_1484;
  reg        [7:0]    _zz_dataOut_payload_0_1485;
  reg        [7:0]    _zz_dataOut_payload_0_1486;
  reg        [7:0]    _zz_dataOut_payload_0_1487;
  reg        [7:0]    _zz_dataOut_payload_0_1488;
  reg        [7:0]    _zz_dataOut_payload_0_1489;
  reg        [7:0]    _zz_dataOut_payload_0_1490;
  reg        [7:0]    _zz_dataOut_payload_0_1491;
  reg        [7:0]    _zz_dataOut_payload_0_1492;
  reg        [7:0]    _zz_dataOut_payload_0_1493;
  reg        [7:0]    _zz_dataOut_payload_0_1494;
  reg        [7:0]    _zz_dataOut_payload_0_1495;
  wire                _zz_dataOut_payload_0_1496;
  wire       [7:0]    _zz_dataOut_payload_0_1497;
  wire       [7:0]    _zz_dataOut_payload_0_1498;
  wire                _zz_dataOut_payload_0_1499;
  wire       [7:0]    _zz_dataOut_payload_0_1500;
  wire       [7:0]    _zz_dataOut_payload_0_1501;
  wire                _zz_dataOut_payload_0_1502;
  wire       [7:0]    _zz_dataOut_payload_0_1503;
  wire       [7:0]    _zz_dataOut_payload_0_1504;
  wire                _zz_dataOut_payload_0_1505;
  wire       [7:0]    _zz_dataOut_payload_0_1506;
  wire       [7:0]    _zz_dataOut_payload_0_1507;
  wire                _zz_dataOut_payload_0_1508;
  wire       [7:0]    _zz_dataOut_payload_0_1509;
  wire       [7:0]    _zz_dataOut_payload_0_1510;
  wire                _zz_dataOut_payload_0_1511;
  wire       [7:0]    _zz_dataOut_payload_0_1512;
  wire       [7:0]    _zz_dataOut_payload_0_1513;
  wire                _zz_dataOut_payload_0_1514;
  wire                _zz_dataOut_payload_0_1515;
  reg        [7:0]    _zz_dataOut_payload_0_1516;
  reg        [7:0]    _zz_dataOut_payload_0_1517;
  reg        [7:0]    _zz_dataOut_payload_0_1518;
  reg        [7:0]    _zz_dataOut_payload_0_1519;
  wire                _zz_dataOut_payload_0_1520;
  wire       [7:0]    _zz_dataOut_payload_0_1521;
  wire       [7:0]    _zz_dataOut_payload_0_1522;
  wire                _zz_dataOut_payload_0_1523;
  wire       [7:0]    _zz_dataOut_payload_0_1524;
  wire       [7:0]    _zz_dataOut_payload_0_1525;
  wire                _zz_dataOut_payload_0_1526;
  wire                _zz_dataOut_payload_0_1527;
  reg        [7:0]    _zz_dataOut_payload_0_1528;
  reg        [7:0]    _zz_dataOut_payload_0_1529;
  reg        [7:0]    _zz_dataOut_payload_0_1530;
  reg        [7:0]    _zz_dataOut_payload_0_1531;
  reg        [7:0]    _zz_dataOut_payload_0_1532;
  reg        [7:0]    _zz_dataOut_payload_0_1533;
  reg        [7:0]    _zz_dataOut_payload_0_1534;
  reg        [7:0]    _zz_dataOut_payload_0_1535;
  reg        [7:0]    _zz_dataOut_payload_0_1536;
  reg        [7:0]    _zz_dataOut_payload_0_1537;
  reg        [7:0]    _zz_dataOut_payload_0_1538;
  reg        [7:0]    _zz_dataOut_payload_0_1539;
  wire                _zz_dataOut_payload_0_1540;
  wire       [7:0]    _zz_dataOut_payload_0_1541;
  wire       [7:0]    _zz_dataOut_payload_0_1542;
  wire                _zz_dataOut_payload_0_1543;
  wire       [7:0]    _zz_dataOut_payload_0_1544;
  wire       [7:0]    _zz_dataOut_payload_0_1545;
  wire                _zz_dataOut_payload_0_1546;
  wire       [7:0]    _zz_dataOut_payload_0_1547;
  wire       [7:0]    _zz_dataOut_payload_0_1548;
  wire                _zz_dataOut_payload_0_1549;
  wire       [7:0]    _zz_dataOut_payload_0_1550;
  wire       [7:0]    _zz_dataOut_payload_0_1551;
  wire                _zz_dataOut_payload_0_1552;
  wire       [7:0]    _zz_dataOut_payload_0_1553;
  wire       [7:0]    _zz_dataOut_payload_0_1554;
  wire                _zz_dataOut_payload_0_1555;
  wire       [7:0]    _zz_dataOut_payload_0_1556;
  wire       [7:0]    _zz_dataOut_payload_0_1557;
  wire                _zz_dataOut_payload_0_1558;
  wire                _zz_dataOut_payload_0_1559;
  reg        [7:0]    _zz_dataOut_payload_0_1560;
  reg        [7:0]    _zz_dataOut_payload_0_1561;
  reg        [7:0]    _zz_dataOut_payload_0_1562;
  reg        [7:0]    _zz_dataOut_payload_0_1563;
  wire                _zz_dataOut_payload_0_1564;
  wire       [7:0]    _zz_dataOut_payload_0_1565;
  wire       [7:0]    _zz_dataOut_payload_0_1566;
  wire                _zz_dataOut_payload_0_1567;
  wire       [7:0]    _zz_dataOut_payload_0_1568;
  wire       [7:0]    _zz_dataOut_payload_0_1569;
  wire                _zz_dataOut_payload_0_1570;
  wire                _zz_dataOut_payload_0_1571;
  reg        [7:0]    _zz_dataOut_payload_0_1572;
  reg        [7:0]    _zz_dataOut_payload_0_1573;
  reg        [7:0]    _zz_dataOut_payload_0_1574;
  reg        [7:0]    _zz_dataOut_payload_0_1575;
  reg        [7:0]    _zz_dataOut_payload_0_1576;
  reg        [7:0]    _zz_dataOut_payload_0_1577;
  reg        [7:0]    _zz_dataOut_payload_0_1578;
  reg        [7:0]    _zz_dataOut_payload_0_1579;
  reg        [7:0]    _zz_dataOut_payload_0_1580;
  reg        [7:0]    _zz_dataOut_payload_0_1581;
  reg        [7:0]    _zz_dataOut_payload_0_1582;
  reg        [7:0]    _zz_dataOut_payload_0_1583;
  wire                _zz_dataOut_payload_0_1584;
  wire       [7:0]    _zz_dataOut_payload_0_1585;
  wire       [7:0]    _zz_dataOut_payload_0_1586;
  wire                _zz_dataOut_payload_0_1587;
  wire       [7:0]    _zz_dataOut_payload_0_1588;
  wire       [7:0]    _zz_dataOut_payload_0_1589;
  wire                _zz_dataOut_payload_0_1590;
  wire       [7:0]    _zz_dataOut_payload_0_1591;
  wire       [7:0]    _zz_dataOut_payload_0_1592;
  wire                _zz_dataOut_payload_0_1593;
  wire       [7:0]    _zz_dataOut_payload_0_1594;
  wire       [7:0]    _zz_dataOut_payload_0_1595;
  wire                _zz_dataOut_payload_0_1596;
  wire       [7:0]    _zz_dataOut_payload_0_1597;
  wire       [7:0]    _zz_dataOut_payload_0_1598;
  wire                _zz_dataOut_payload_0_1599;
  wire       [7:0]    _zz_dataOut_payload_0_1600;
  wire       [7:0]    _zz_dataOut_payload_0_1601;
  wire                _zz_dataOut_payload_0_1602;
  wire                _zz_dataOut_payload_0_1603;
  reg        [7:0]    _zz_dataOut_payload_0_1604;
  reg        [7:0]    _zz_dataOut_payload_0_1605;
  reg        [7:0]    _zz_dataOut_payload_0_1606;
  reg        [7:0]    _zz_dataOut_payload_0_1607;
  wire                _zz_dataOut_payload_0_1608;
  wire       [7:0]    _zz_dataOut_payload_0_1609;
  wire       [7:0]    _zz_dataOut_payload_0_1610;
  wire                _zz_dataOut_payload_0_1611;
  wire       [7:0]    _zz_dataOut_payload_0_1612;
  wire       [7:0]    _zz_dataOut_payload_0_1613;
  wire                _zz_dataOut_payload_0_1614;
  wire                _zz_dataOut_payload_0_1615;
  reg        [7:0]    _zz_dataOut_payload_0_1616;
  reg        [7:0]    _zz_dataOut_payload_0_1617;
  reg        [7:0]    _zz_dataOut_payload_0_1618;
  reg        [7:0]    _zz_dataOut_payload_0_1619;
  reg        [7:0]    _zz_dataOut_payload_0_1620;
  reg        [7:0]    _zz_dataOut_payload_0_1621;
  reg        [7:0]    _zz_dataOut_payload_0_1622;
  reg        [7:0]    _zz_dataOut_payload_0_1623;
  reg        [7:0]    _zz_dataOut_payload_0_1624;
  reg        [7:0]    _zz_dataOut_payload_0_1625;
  reg        [7:0]    _zz_dataOut_payload_0_1626;
  reg        [7:0]    _zz_dataOut_payload_0_1627;
  wire                _zz_dataOut_payload_0_1628;
  wire       [7:0]    _zz_dataOut_payload_0_1629;
  wire       [7:0]    _zz_dataOut_payload_0_1630;
  wire                _zz_dataOut_payload_0_1631;
  wire       [7:0]    _zz_dataOut_payload_0_1632;
  wire       [7:0]    _zz_dataOut_payload_0_1633;
  wire                _zz_dataOut_payload_0_1634;
  wire       [7:0]    _zz_dataOut_payload_0_1635;
  wire       [7:0]    _zz_dataOut_payload_0_1636;
  wire                _zz_dataOut_payload_0_1637;
  wire       [7:0]    _zz_dataOut_payload_0_1638;
  wire       [7:0]    _zz_dataOut_payload_0_1639;
  wire                _zz_dataOut_payload_0_1640;
  wire       [7:0]    _zz_dataOut_payload_0_1641;
  wire       [7:0]    _zz_dataOut_payload_0_1642;
  wire                _zz_dataOut_payload_0_1643;
  wire       [7:0]    _zz_dataOut_payload_0_1644;
  wire       [7:0]    _zz_dataOut_payload_0_1645;
  wire                _zz_dataOut_payload_0_1646;
  wire                _zz_dataOut_payload_0_1647;
  reg        [7:0]    _zz_dataOut_payload_0_1648;
  reg        [7:0]    _zz_dataOut_payload_0_1649;
  reg        [7:0]    _zz_dataOut_payload_0_1650;
  reg        [7:0]    _zz_dataOut_payload_0_1651;
  wire                _zz_dataOut_payload_0_1652;
  wire       [7:0]    _zz_dataOut_payload_0_1653;
  wire       [7:0]    _zz_dataOut_payload_0_1654;
  wire                _zz_dataOut_payload_0_1655;
  wire       [7:0]    _zz_dataOut_payload_0_1656;
  wire       [7:0]    _zz_dataOut_payload_0_1657;
  wire                _zz_dataOut_payload_0_1658;
  wire                _zz_dataOut_payload_0_1659;
  reg        [7:0]    _zz_dataOut_payload_0_1660;
  reg        [7:0]    _zz_dataOut_payload_0_1661;
  reg        [7:0]    _zz_dataOut_payload_0_1662;
  reg        [7:0]    _zz_dataOut_payload_0_1663;
  reg        [7:0]    _zz_dataOut_payload_0_1664;
  reg        [7:0]    _zz_dataOut_payload_0_1665;
  reg        [7:0]    _zz_dataOut_payload_0_1666;
  reg        [7:0]    _zz_dataOut_payload_0_1667;
  reg        [7:0]    _zz_dataOut_payload_0_1668;
  reg        [7:0]    _zz_dataOut_payload_0_1669;
  reg        [7:0]    _zz_dataOut_payload_0_1670;
  reg        [7:0]    _zz_dataOut_payload_0_1671;
  wire                _zz_dataOut_payload_0_1672;
  wire       [7:0]    _zz_dataOut_payload_0_1673;
  wire       [7:0]    _zz_dataOut_payload_0_1674;
  wire                _zz_dataOut_payload_0_1675;
  wire       [7:0]    _zz_dataOut_payload_0_1676;
  wire       [7:0]    _zz_dataOut_payload_0_1677;
  wire                _zz_dataOut_payload_0_1678;
  wire       [7:0]    _zz_dataOut_payload_0_1679;
  wire       [7:0]    _zz_dataOut_payload_0_1680;
  wire                _zz_dataOut_payload_0_1681;
  wire       [7:0]    _zz_dataOut_payload_0_1682;
  wire       [7:0]    _zz_dataOut_payload_0_1683;
  wire                _zz_dataOut_payload_0_1684;
  wire       [7:0]    _zz_dataOut_payload_0_1685;
  wire       [7:0]    _zz_dataOut_payload_0_1686;
  wire                _zz_dataOut_payload_0_1687;
  wire       [7:0]    _zz_dataOut_payload_0_1688;
  wire       [7:0]    _zz_dataOut_payload_0_1689;
  wire                _zz_dataOut_payload_0_1690;
  wire                _zz_dataOut_payload_0_1691;
  reg        [7:0]    _zz_dataOut_payload_0_1692;
  reg        [7:0]    _zz_dataOut_payload_0_1693;
  reg        [7:0]    _zz_dataOut_payload_0_1694;
  reg        [7:0]    _zz_dataOut_payload_0_1695;
  wire                _zz_dataOut_payload_0_1696;
  wire       [7:0]    _zz_dataOut_payload_0_1697;
  wire       [7:0]    _zz_dataOut_payload_0_1698;
  wire                _zz_dataOut_payload_0_1699;
  wire       [7:0]    _zz_dataOut_payload_0_1700;
  wire       [7:0]    _zz_dataOut_payload_0_1701;
  wire                _zz_dataOut_payload_0_1702;
  wire                _zz_dataOut_payload_0_1703;
  reg        [7:0]    _zz_dataOut_payload_0_1704;
  reg        [7:0]    _zz_dataOut_payload_0_1705;
  reg        [7:0]    _zz_dataOut_payload_0_1706;
  reg        [7:0]    _zz_dataOut_payload_0_1707;
  reg        [7:0]    _zz_dataOut_payload_0_1708;
  reg        [7:0]    _zz_dataOut_payload_0_1709;
  reg        [7:0]    _zz_dataOut_payload_0_1710;
  reg        [7:0]    _zz_dataOut_payload_0_1711;
  reg        [7:0]    _zz_dataOut_payload_0_1712;
  reg        [7:0]    _zz_dataOut_payload_0_1713;
  reg        [7:0]    _zz_dataOut_payload_0_1714;
  reg        [7:0]    _zz_dataOut_payload_0_1715;
  wire                _zz_dataOut_payload_0_1716;
  wire       [7:0]    _zz_dataOut_payload_0_1717;
  wire       [7:0]    _zz_dataOut_payload_0_1718;
  wire                _zz_dataOut_payload_0_1719;
  wire       [7:0]    _zz_dataOut_payload_0_1720;
  wire       [7:0]    _zz_dataOut_payload_0_1721;
  wire                _zz_dataOut_payload_0_1722;
  wire       [7:0]    _zz_dataOut_payload_0_1723;
  wire       [7:0]    _zz_dataOut_payload_0_1724;
  wire                _zz_dataOut_payload_0_1725;
  wire       [7:0]    _zz_dataOut_payload_0_1726;
  wire       [7:0]    _zz_dataOut_payload_0_1727;
  wire                _zz_dataOut_payload_0_1728;
  wire       [7:0]    _zz_dataOut_payload_0_1729;
  wire       [7:0]    _zz_dataOut_payload_0_1730;
  wire                _zz_dataOut_payload_0_1731;
  wire       [7:0]    _zz_dataOut_payload_0_1732;
  wire       [7:0]    _zz_dataOut_payload_0_1733;
  wire                _zz_dataOut_payload_0_1734;
  wire                _zz_dataOut_payload_0_1735;
  reg        [7:0]    _zz_dataOut_payload_0_1736;
  reg        [7:0]    _zz_dataOut_payload_0_1737;
  reg        [7:0]    _zz_dataOut_payload_0_1738;
  reg        [7:0]    _zz_dataOut_payload_0_1739;
  wire                _zz_dataOut_payload_0_1740;
  wire       [7:0]    _zz_dataOut_payload_0_1741;
  wire       [7:0]    _zz_dataOut_payload_0_1742;
  wire                _zz_dataOut_payload_0_1743;
  wire       [7:0]    _zz_dataOut_payload_0_1744;
  wire       [7:0]    _zz_dataOut_payload_0_1745;
  wire                _zz_dataOut_payload_0_1746;
  wire                _zz_dataOut_payload_0_1747;
  reg        [7:0]    _zz_dataOut_payload_0_1748;
  reg        [7:0]    _zz_dataOut_payload_0_1749;
  reg        [7:0]    _zz_dataOut_payload_0_1750;
  reg        [7:0]    _zz_dataOut_payload_0_1751;
  reg        [7:0]    _zz_dataOut_payload_0_1752;
  reg        [7:0]    _zz_dataOut_payload_0_1753;
  reg        [7:0]    _zz_dataOut_payload_0_1754;
  reg        [7:0]    _zz_dataOut_payload_0_1755;
  reg        [7:0]    _zz_dataOut_payload_0_1756;
  reg        [7:0]    _zz_dataOut_payload_0_1757;
  reg        [7:0]    _zz_dataOut_payload_0_1758;
  reg        [7:0]    _zz_dataOut_payload_0_1759;
  wire                _zz_dataOut_payload_0_1760;
  wire       [7:0]    _zz_dataOut_payload_0_1761;
  wire       [7:0]    _zz_dataOut_payload_0_1762;
  wire                _zz_dataOut_payload_0_1763;
  wire       [7:0]    _zz_dataOut_payload_0_1764;
  wire       [7:0]    _zz_dataOut_payload_0_1765;
  wire                _zz_dataOut_payload_0_1766;
  wire       [7:0]    _zz_dataOut_payload_0_1767;
  wire       [7:0]    _zz_dataOut_payload_0_1768;
  wire                _zz_dataOut_payload_0_1769;
  wire       [7:0]    _zz_dataOut_payload_0_1770;
  wire       [7:0]    _zz_dataOut_payload_0_1771;
  wire                _zz_dataOut_payload_0_1772;
  wire       [7:0]    _zz_dataOut_payload_0_1773;
  wire       [7:0]    _zz_dataOut_payload_0_1774;
  wire                _zz_dataOut_payload_0_1775;
  wire       [7:0]    _zz_dataOut_payload_0_1776;
  wire       [7:0]    _zz_dataOut_payload_0_1777;
  wire                _zz_dataOut_payload_0_1778;
  wire                _zz_dataOut_payload_0_1779;
  reg        [7:0]    _zz_dataOut_payload_0_1780;
  reg        [7:0]    _zz_dataOut_payload_0_1781;
  reg        [7:0]    _zz_dataOut_payload_0_1782;
  reg        [7:0]    _zz_dataOut_payload_0_1783;
  wire                _zz_dataOut_payload_0_1784;
  wire       [7:0]    _zz_dataOut_payload_0_1785;
  wire       [7:0]    _zz_dataOut_payload_0_1786;
  wire                _zz_dataOut_payload_0_1787;
  wire       [7:0]    _zz_dataOut_payload_0_1788;
  wire       [7:0]    _zz_dataOut_payload_0_1789;
  wire                _zz_dataOut_payload_0_1790;
  wire                _zz_dataOut_payload_0_1791;
  reg        [7:0]    _zz_dataOut_payload_0_1792;
  reg        [7:0]    _zz_dataOut_payload_0_1793;
  reg        [7:0]    _zz_dataOut_payload_0_1794;
  reg        [7:0]    _zz_dataOut_payload_0_1795;
  reg        [7:0]    _zz_dataOut_payload_0_1796;
  reg        [7:0]    _zz_dataOut_payload_0_1797;
  reg        [7:0]    _zz_dataOut_payload_0_1798;
  reg        [7:0]    _zz_dataOut_payload_0_1799;
  reg        [7:0]    _zz_dataOut_payload_0_1800;
  reg        [7:0]    _zz_dataOut_payload_0_1801;
  reg        [7:0]    _zz_dataOut_payload_0_1802;
  reg        [7:0]    _zz_dataOut_payload_0_1803;
  wire                _zz_dataOut_payload_0_1804;
  wire       [7:0]    _zz_dataOut_payload_0_1805;
  wire       [7:0]    _zz_dataOut_payload_0_1806;
  wire                _zz_dataOut_payload_0_1807;
  wire       [7:0]    _zz_dataOut_payload_0_1808;
  wire       [7:0]    _zz_dataOut_payload_0_1809;
  wire                _zz_dataOut_payload_0_1810;
  wire       [7:0]    _zz_dataOut_payload_0_1811;
  wire       [7:0]    _zz_dataOut_payload_0_1812;
  wire                _zz_dataOut_payload_0_1813;
  wire       [7:0]    _zz_dataOut_payload_0_1814;
  wire       [7:0]    _zz_dataOut_payload_0_1815;
  wire                _zz_dataOut_payload_0_1816;
  wire       [7:0]    _zz_dataOut_payload_0_1817;
  wire       [7:0]    _zz_dataOut_payload_0_1818;
  wire                _zz_dataOut_payload_0_1819;
  wire       [7:0]    _zz_dataOut_payload_0_1820;
  wire       [7:0]    _zz_dataOut_payload_0_1821;
  wire                _zz_dataOut_payload_0_1822;
  wire                _zz_dataOut_payload_0_1823;
  reg        [7:0]    _zz_dataOut_payload_0_1824;
  reg        [7:0]    _zz_dataOut_payload_0_1825;
  reg        [7:0]    _zz_dataOut_payload_0_1826;
  reg        [7:0]    _zz_dataOut_payload_0_1827;
  wire                _zz_dataOut_payload_0_1828;
  wire       [7:0]    _zz_dataOut_payload_0_1829;
  wire       [7:0]    _zz_dataOut_payload_0_1830;
  wire                _zz_dataOut_payload_0_1831;
  wire       [7:0]    _zz_dataOut_payload_0_1832;
  wire       [7:0]    _zz_dataOut_payload_0_1833;
  wire                _zz_dataOut_payload_0_1834;
  wire                _zz_dataOut_payload_0_1835;
  reg        [7:0]    _zz_dataOut_payload_0_1836;
  reg        [7:0]    _zz_dataOut_payload_0_1837;
  reg        [7:0]    _zz_dataOut_payload_0_1838;
  reg        [7:0]    _zz_dataOut_payload_0_1839;
  reg        [7:0]    _zz_dataOut_payload_0_1840;
  reg        [7:0]    _zz_dataOut_payload_0_1841;
  reg        [7:0]    _zz_dataOut_payload_0_1842;
  reg        [7:0]    _zz_dataOut_payload_0_1843;
  reg        [7:0]    _zz_dataOut_payload_0_1844;
  reg        [7:0]    _zz_dataOut_payload_0_1845;
  reg        [7:0]    _zz_dataOut_payload_0_1846;
  reg        [7:0]    _zz_dataOut_payload_0_1847;
  wire                _zz_dataOut_payload_0_1848;
  wire       [7:0]    _zz_dataOut_payload_0_1849;
  wire       [7:0]    _zz_dataOut_payload_0_1850;
  wire                _zz_dataOut_payload_0_1851;
  wire       [7:0]    _zz_dataOut_payload_0_1852;
  wire       [7:0]    _zz_dataOut_payload_0_1853;
  wire                _zz_dataOut_payload_0_1854;
  wire       [7:0]    _zz_dataOut_payload_0_1855;
  wire       [7:0]    _zz_dataOut_payload_0_1856;
  wire                _zz_dataOut_payload_0_1857;
  wire       [7:0]    _zz_dataOut_payload_0_1858;
  wire       [7:0]    _zz_dataOut_payload_0_1859;
  wire                _zz_dataOut_payload_0_1860;
  wire       [7:0]    _zz_dataOut_payload_0_1861;
  wire       [7:0]    _zz_dataOut_payload_0_1862;
  wire                _zz_dataOut_payload_0_1863;
  wire       [7:0]    _zz_dataOut_payload_0_1864;
  wire       [7:0]    _zz_dataOut_payload_0_1865;
  wire                _zz_dataOut_payload_0_1866;
  wire                _zz_dataOut_payload_0_1867;
  reg        [7:0]    _zz_dataOut_payload_0_1868;
  reg        [7:0]    _zz_dataOut_payload_0_1869;
  reg        [7:0]    _zz_dataOut_payload_0_1870;
  reg        [7:0]    _zz_dataOut_payload_0_1871;
  wire                _zz_dataOut_payload_0_1872;
  wire       [7:0]    _zz_dataOut_payload_0_1873;
  wire       [7:0]    _zz_dataOut_payload_0_1874;
  wire                _zz_dataOut_payload_0_1875;
  wire       [7:0]    _zz_dataOut_payload_0_1876;
  wire       [7:0]    _zz_dataOut_payload_0_1877;
  wire                _zz_dataOut_payload_0_1878;
  wire                _zz_dataOut_payload_0_1879;
  reg        [7:0]    _zz_dataOut_payload_0_1880;
  reg        [7:0]    _zz_dataOut_payload_0_1881;
  reg        [7:0]    _zz_dataOut_payload_0_1882;
  reg        [7:0]    _zz_dataOut_payload_0_1883;
  reg        [7:0]    _zz_dataOut_payload_0_1884;
  reg        [7:0]    _zz_dataOut_payload_0_1885;
  reg        [7:0]    _zz_dataOut_payload_0_1886;
  reg        [7:0]    _zz_dataOut_payload_0_1887;
  reg        [7:0]    _zz_dataOut_payload_0_1888;
  reg        [7:0]    _zz_dataOut_payload_0_1889;
  reg        [7:0]    _zz_dataOut_payload_0_1890;
  reg        [7:0]    _zz_dataOut_payload_0_1891;
  wire                _zz_dataOut_payload_0_1892;
  wire       [7:0]    _zz_dataOut_payload_0_1893;
  wire       [7:0]    _zz_dataOut_payload_0_1894;
  wire                _zz_dataOut_payload_0_1895;
  wire       [7:0]    _zz_dataOut_payload_0_1896;
  wire       [7:0]    _zz_dataOut_payload_0_1897;
  wire                _zz_dataOut_payload_0_1898;
  wire       [7:0]    _zz_dataOut_payload_0_1899;
  wire       [7:0]    _zz_dataOut_payload_0_1900;
  wire                _zz_dataOut_payload_0_1901;
  wire       [7:0]    _zz_dataOut_payload_0_1902;
  wire       [7:0]    _zz_dataOut_payload_0_1903;
  wire                _zz_dataOut_payload_0_1904;
  wire       [7:0]    _zz_dataOut_payload_0_1905;
  wire       [7:0]    _zz_dataOut_payload_0_1906;
  wire                _zz_dataOut_payload_0_1907;
  wire       [7:0]    _zz_dataOut_payload_0_1908;
  wire       [7:0]    _zz_dataOut_payload_0_1909;
  wire                _zz_dataOut_payload_0_1910;
  wire                _zz_dataOut_payload_0_1911;
  reg        [7:0]    _zz_dataOut_payload_0_1912;
  reg        [7:0]    _zz_dataOut_payload_0_1913;
  reg        [7:0]    _zz_dataOut_payload_0_1914;
  reg        [7:0]    _zz_dataOut_payload_0_1915;
  wire                _zz_dataOut_payload_0_1916;
  wire       [7:0]    _zz_dataOut_payload_0_1917;
  wire       [7:0]    _zz_dataOut_payload_0_1918;
  wire                _zz_dataOut_payload_0_1919;
  wire       [7:0]    _zz_dataOut_payload_0_1920;
  wire       [7:0]    _zz_dataOut_payload_0_1921;
  wire                _zz_dataOut_payload_0_1922;
  wire                _zz_dataOut_payload_0_1923;
  reg        [7:0]    _zz_dataOut_payload_0_1924;
  reg        [7:0]    _zz_dataOut_payload_0_1925;
  reg        [7:0]    _zz_dataOut_payload_0_1926;
  reg        [7:0]    _zz_dataOut_payload_0_1927;
  reg        [7:0]    _zz_dataOut_payload_0_1928;
  reg        [7:0]    _zz_dataOut_payload_0_1929;
  reg        [7:0]    _zz_dataOut_payload_0_1930;
  reg        [7:0]    _zz_dataOut_payload_0_1931;
  reg        [7:0]    _zz_dataOut_payload_0_1932;
  reg        [7:0]    _zz_dataOut_payload_0_1933;
  reg        [7:0]    _zz_dataOut_payload_0_1934;
  reg        [7:0]    _zz_dataOut_payload_0_1935;
  wire                _zz_dataOut_payload_0_1936;
  wire       [7:0]    _zz_dataOut_payload_0_1937;
  wire       [7:0]    _zz_dataOut_payload_0_1938;
  wire                _zz_dataOut_payload_0_1939;
  wire       [7:0]    _zz_dataOut_payload_0_1940;
  wire       [7:0]    _zz_dataOut_payload_0_1941;
  wire                _zz_dataOut_payload_0_1942;
  wire       [7:0]    _zz_dataOut_payload_0_1943;
  wire       [7:0]    _zz_dataOut_payload_0_1944;
  wire                _zz_dataOut_payload_0_1945;
  wire       [7:0]    _zz_dataOut_payload_0_1946;
  wire       [7:0]    _zz_dataOut_payload_0_1947;
  wire                _zz_dataOut_payload_0_1948;
  wire       [7:0]    _zz_dataOut_payload_0_1949;
  wire       [7:0]    _zz_dataOut_payload_0_1950;
  wire                _zz_dataOut_payload_0_1951;
  wire       [7:0]    _zz_dataOut_payload_0_1952;
  wire       [7:0]    _zz_dataOut_payload_0_1953;
  wire                _zz_dataOut_payload_0_1954;
  wire                _zz_dataOut_payload_0_1955;
  reg        [7:0]    _zz_dataOut_payload_0_1956;
  reg        [7:0]    _zz_dataOut_payload_0_1957;
  reg        [7:0]    _zz_dataOut_payload_0_1958;
  reg        [7:0]    _zz_dataOut_payload_0_1959;
  wire                _zz_dataOut_payload_0_1960;
  wire       [7:0]    _zz_dataOut_payload_0_1961;
  wire       [7:0]    _zz_dataOut_payload_0_1962;
  wire                _zz_dataOut_payload_0_1963;
  wire       [7:0]    _zz_dataOut_payload_0_1964;
  wire       [7:0]    _zz_dataOut_payload_0_1965;
  wire                _zz_dataOut_payload_0_1966;
  wire                _zz_dataOut_payload_0_1967;
  reg        [7:0]    _zz_dataOut_payload_0_1968;
  reg        [7:0]    _zz_dataOut_payload_0_1969;
  reg        [7:0]    _zz_dataOut_payload_0_1970;
  reg        [7:0]    _zz_dataOut_payload_0_1971;
  reg        [7:0]    _zz_dataOut_payload_0_1972;
  reg        [7:0]    _zz_dataOut_payload_0_1973;
  reg        [7:0]    _zz_dataOut_payload_0_1974;
  reg        [7:0]    _zz_dataOut_payload_0_1975;
  reg        [7:0]    _zz_dataOut_payload_0_1976;
  reg        [7:0]    _zz_dataOut_payload_0_1977;
  reg        [7:0]    _zz_dataOut_payload_0_1978;
  reg        [7:0]    _zz_dataOut_payload_0_1979;
  wire                _zz_dataOut_payload_0_1980;
  wire       [7:0]    _zz_dataOut_payload_0_1981;
  wire       [7:0]    _zz_dataOut_payload_0_1982;
  wire                _zz_dataOut_payload_0_1983;
  wire       [7:0]    _zz_dataOut_payload_0_1984;
  wire       [7:0]    _zz_dataOut_payload_0_1985;
  wire                _zz_dataOut_payload_0_1986;
  wire       [7:0]    _zz_dataOut_payload_0_1987;
  wire       [7:0]    _zz_dataOut_payload_0_1988;
  wire                _zz_dataOut_payload_0_1989;
  wire       [7:0]    _zz_dataOut_payload_0_1990;
  wire       [7:0]    _zz_dataOut_payload_0_1991;
  wire                _zz_dataOut_payload_0_1992;
  wire       [7:0]    _zz_dataOut_payload_0_1993;
  wire       [7:0]    _zz_dataOut_payload_0_1994;
  wire                _zz_dataOut_payload_0_1995;
  wire       [7:0]    _zz_dataOut_payload_0_1996;
  wire       [7:0]    _zz_dataOut_payload_0_1997;
  wire                _zz_dataOut_payload_0_1998;
  wire                _zz_dataOut_payload_0_1999;
  reg        [7:0]    _zz_dataOut_payload_0_2000;
  reg        [7:0]    _zz_dataOut_payload_0_2001;
  reg        [7:0]    _zz_dataOut_payload_0_2002;
  reg        [7:0]    _zz_dataOut_payload_0_2003;
  wire                _zz_dataOut_payload_0_2004;
  wire       [7:0]    _zz_dataOut_payload_0_2005;
  wire       [7:0]    _zz_dataOut_payload_0_2006;
  wire                _zz_dataOut_payload_0_2007;
  wire       [7:0]    _zz_dataOut_payload_0_2008;
  wire       [7:0]    _zz_dataOut_payload_0_2009;
  wire                _zz_dataOut_payload_0_2010;
  wire                _zz_dataOut_payload_0_2011;
  reg        [7:0]    _zz_dataOut_payload_0_2012;
  reg        [7:0]    _zz_dataOut_payload_0_2013;
  reg        [7:0]    _zz_dataOut_payload_0_2014;
  reg        [7:0]    _zz_dataOut_payload_0_2015;
  reg        [7:0]    _zz_dataOut_payload_0_2016;
  reg        [7:0]    _zz_dataOut_payload_0_2017;
  reg        [7:0]    _zz_dataOut_payload_0_2018;
  reg        [7:0]    _zz_dataOut_payload_0_2019;
  reg        [7:0]    _zz_dataOut_payload_0_2020;
  reg        [7:0]    _zz_dataOut_payload_0_2021;
  reg        [7:0]    _zz_dataOut_payload_0_2022;
  reg        [7:0]    _zz_dataOut_payload_0_2023;
  wire                _zz_dataOut_payload_0_2024;
  wire       [7:0]    _zz_dataOut_payload_0_2025;
  wire       [7:0]    _zz_dataOut_payload_0_2026;
  wire                _zz_dataOut_payload_0_2027;
  wire       [7:0]    _zz_dataOut_payload_0_2028;
  wire       [7:0]    _zz_dataOut_payload_0_2029;
  wire                _zz_dataOut_payload_0_2030;
  wire       [7:0]    _zz_dataOut_payload_0_2031;
  wire       [7:0]    _zz_dataOut_payload_0_2032;
  wire                _zz_dataOut_payload_0_2033;
  wire       [7:0]    _zz_dataOut_payload_0_2034;
  wire       [7:0]    _zz_dataOut_payload_0_2035;
  wire                _zz_dataOut_payload_0_2036;
  wire       [7:0]    _zz_dataOut_payload_0_2037;
  wire       [7:0]    _zz_dataOut_payload_0_2038;
  wire                _zz_dataOut_payload_0_2039;
  wire       [7:0]    _zz_dataOut_payload_0_2040;
  wire       [7:0]    _zz_dataOut_payload_0_2041;
  wire                _zz_dataOut_payload_0_2042;
  wire                _zz_dataOut_payload_0_2043;
  reg        [7:0]    _zz_dataOut_payload_0_2044;
  reg        [7:0]    _zz_dataOut_payload_0_2045;
  reg        [7:0]    _zz_dataOut_payload_0_2046;
  reg        [7:0]    _zz_dataOut_payload_0_2047;
  wire                _zz_dataOut_payload_0_2048;
  wire       [7:0]    _zz_dataOut_payload_0_2049;
  wire       [7:0]    _zz_dataOut_payload_0_2050;
  wire                _zz_dataOut_payload_0_2051;
  wire       [7:0]    _zz_dataOut_payload_0_2052;
  wire       [7:0]    _zz_dataOut_payload_0_2053;
  wire                _zz_dataOut_payload_0_2054;
  wire                _zz_dataOut_payload_0_2055;
  reg        [7:0]    _zz_dataOut_payload_0_2056;
  reg        [7:0]    _zz_dataOut_payload_0_2057;
  reg        [7:0]    _zz_dataOut_payload_0_2058;
  reg        [7:0]    _zz_dataOut_payload_0_2059;
  reg        [7:0]    _zz_dataOut_payload_0_2060;
  reg        [7:0]    _zz_dataOut_payload_0_2061;
  reg        [7:0]    _zz_dataOut_payload_0_2062;
  reg        [7:0]    _zz_dataOut_payload_0_2063;
  reg        [7:0]    _zz_dataOut_payload_0_2064;
  reg        [7:0]    _zz_dataOut_payload_0_2065;
  reg        [7:0]    _zz_dataOut_payload_0_2066;
  reg        [7:0]    _zz_dataOut_payload_0_2067;
  wire                _zz_dataOut_payload_0_2068;
  wire       [7:0]    _zz_dataOut_payload_0_2069;
  wire       [7:0]    _zz_dataOut_payload_0_2070;
  wire                _zz_dataOut_payload_0_2071;
  wire       [7:0]    _zz_dataOut_payload_0_2072;
  wire       [7:0]    _zz_dataOut_payload_0_2073;
  wire                _zz_dataOut_payload_0_2074;
  wire       [7:0]    _zz_dataOut_payload_0_2075;
  wire       [7:0]    _zz_dataOut_payload_0_2076;
  wire                _zz_dataOut_payload_0_2077;
  wire       [7:0]    _zz_dataOut_payload_0_2078;
  wire       [7:0]    _zz_dataOut_payload_0_2079;
  wire                _zz_dataOut_payload_0_2080;
  wire       [7:0]    _zz_dataOut_payload_0_2081;
  wire       [7:0]    _zz_dataOut_payload_0_2082;
  wire                _zz_dataOut_payload_0_2083;
  wire       [7:0]    _zz_dataOut_payload_0_2084;
  wire       [7:0]    _zz_dataOut_payload_0_2085;
  wire                _zz_dataOut_payload_0_2086;
  wire                _zz_dataOut_payload_0_2087;
  reg        [7:0]    _zz_dataOut_payload_0_2088;
  reg        [7:0]    _zz_dataOut_payload_0_2089;
  reg        [7:0]    _zz_dataOut_payload_0_2090;
  reg        [7:0]    _zz_dataOut_payload_0_2091;
  wire                _zz_dataOut_payload_0_2092;
  wire       [7:0]    _zz_dataOut_payload_0_2093;
  wire       [7:0]    _zz_dataOut_payload_0_2094;
  wire                _zz_dataOut_payload_0_2095;
  wire       [7:0]    _zz_dataOut_payload_0_2096;
  wire       [7:0]    _zz_dataOut_payload_0_2097;
  wire                _zz_dataOut_payload_0_2098;
  wire                _zz_dataOut_payload_0_2099;
  reg        [7:0]    _zz_dataOut_payload_0_2100;
  reg        [7:0]    _zz_dataOut_payload_0_2101;
  reg        [7:0]    _zz_dataOut_payload_0_2102;
  reg        [7:0]    _zz_dataOut_payload_0_2103;
  reg        [7:0]    _zz_dataOut_payload_0_2104;
  reg        [7:0]    _zz_dataOut_payload_0_2105;
  reg        [7:0]    _zz_dataOut_payload_0_2106;
  reg        [7:0]    _zz_dataOut_payload_0_2107;
  reg        [7:0]    _zz_dataOut_payload_0_2108;
  reg        [7:0]    _zz_dataOut_payload_0_2109;
  reg        [7:0]    _zz_dataOut_payload_0_2110;
  reg        [7:0]    _zz_dataOut_payload_0_2111;
  wire                _zz_dataOut_payload_0_2112;
  wire       [7:0]    _zz_dataOut_payload_0_2113;
  wire       [7:0]    _zz_dataOut_payload_0_2114;
  wire                _zz_dataOut_payload_0_2115;
  wire       [7:0]    _zz_dataOut_payload_0_2116;
  wire       [7:0]    _zz_dataOut_payload_0_2117;
  wire                _zz_dataOut_payload_0_2118;
  wire       [7:0]    _zz_dataOut_payload_0_2119;
  wire       [7:0]    _zz_dataOut_payload_0_2120;
  wire                _zz_dataOut_payload_0_2121;
  wire       [7:0]    _zz_dataOut_payload_0_2122;
  wire       [7:0]    _zz_dataOut_payload_0_2123;
  wire                _zz_dataOut_payload_0_2124;
  wire       [7:0]    _zz_dataOut_payload_0_2125;
  wire       [7:0]    _zz_dataOut_payload_0_2126;
  wire                _zz_dataOut_payload_0_2127;
  wire       [7:0]    _zz_dataOut_payload_0_2128;
  wire       [7:0]    _zz_dataOut_payload_0_2129;
  wire                _zz_dataOut_payload_0_2130;
  wire                _zz_dataOut_payload_0_2131;
  reg        [7:0]    _zz_dataOut_payload_0_2132;
  reg        [7:0]    _zz_dataOut_payload_0_2133;
  reg        [7:0]    _zz_dataOut_payload_0_2134;
  reg        [7:0]    _zz_dataOut_payload_0_2135;
  wire                _zz_dataOut_payload_0_2136;
  wire       [7:0]    _zz_dataOut_payload_0_2137;
  wire       [7:0]    _zz_dataOut_payload_0_2138;
  wire                _zz_dataOut_payload_0_2139;
  wire       [7:0]    _zz_dataOut_payload_0_2140;
  wire       [7:0]    _zz_dataOut_payload_0_2141;
  wire                _zz_dataOut_payload_0_2142;
  wire                _zz_dataOut_payload_0_2143;
  reg        [7:0]    _zz_dataOut_payload_0_2144;
  reg        [7:0]    _zz_dataOut_payload_0_2145;
  reg        [7:0]    _zz_dataOut_payload_0_2146;
  reg        [7:0]    _zz_dataOut_payload_0_2147;
  reg        [7:0]    _zz_dataOut_payload_0_2148;
  reg        [7:0]    _zz_dataOut_payload_0_2149;
  reg        [7:0]    _zz_dataOut_payload_0_2150;
  reg        [7:0]    _zz_dataOut_payload_0_2151;
  reg        [7:0]    _zz_dataOut_payload_0_2152;
  reg        [7:0]    _zz_dataOut_payload_0_2153;
  reg        [7:0]    _zz_dataOut_payload_0_2154;
  reg        [7:0]    _zz_dataOut_payload_0_2155;
  wire                _zz_dataOut_payload_0_2156;
  wire       [7:0]    _zz_dataOut_payload_0_2157;
  wire       [7:0]    _zz_dataOut_payload_0_2158;
  wire                _zz_dataOut_payload_0_2159;
  wire       [7:0]    _zz_dataOut_payload_0_2160;
  wire       [7:0]    _zz_dataOut_payload_0_2161;
  wire                _zz_dataOut_payload_0_2162;
  wire       [7:0]    _zz_dataOut_payload_0_2163;
  wire       [7:0]    _zz_dataOut_payload_0_2164;
  wire                _zz_dataOut_payload_0_2165;
  wire       [7:0]    _zz_dataOut_payload_0_2166;
  wire       [7:0]    _zz_dataOut_payload_0_2167;
  wire                _zz_dataOut_payload_0_2168;
  wire       [7:0]    _zz_dataOut_payload_0_2169;
  wire       [7:0]    _zz_dataOut_payload_0_2170;
  wire                _zz_dataOut_payload_0_2171;
  wire       [7:0]    _zz_dataOut_payload_0_2172;
  wire       [7:0]    _zz_dataOut_payload_0_2173;
  wire                _zz_dataOut_payload_0_2174;
  wire                _zz_dataOut_payload_0_2175;
  reg        [7:0]    _zz_dataOut_payload_0_2176;
  reg        [7:0]    _zz_dataOut_payload_0_2177;
  reg        [7:0]    _zz_dataOut_payload_0_2178;
  reg        [7:0]    _zz_dataOut_payload_0_2179;
  wire                _zz_dataOut_payload_0_2180;
  wire       [7:0]    _zz_dataOut_payload_0_2181;
  wire       [7:0]    _zz_dataOut_payload_0_2182;
  wire                _zz_dataOut_payload_0_2183;
  wire       [7:0]    _zz_dataOut_payload_0_2184;
  wire       [7:0]    _zz_dataOut_payload_0_2185;
  wire                _zz_dataOut_payload_0_2186;
  wire                _zz_dataOut_payload_0_2187;
  reg        [7:0]    _zz_dataOut_payload_0_2188;
  reg        [7:0]    _zz_dataOut_payload_0_2189;
  reg        [7:0]    _zz_dataOut_payload_0_2190;
  reg        [7:0]    _zz_dataOut_payload_0_2191;
  reg        [7:0]    _zz_dataOut_payload_0_2192;
  reg        [7:0]    _zz_dataOut_payload_0_2193;
  reg        [7:0]    _zz_dataOut_payload_0_2194;
  reg        [7:0]    _zz_dataOut_payload_0_2195;
  reg        [7:0]    _zz_dataOut_payload_0_2196;
  reg        [7:0]    _zz_dataOut_payload_0_2197;
  reg        [7:0]    _zz_dataOut_payload_0_2198;
  reg        [7:0]    _zz_dataOut_payload_0_2199;
  wire                _zz_dataOut_payload_0_2200;
  wire       [7:0]    _zz_dataOut_payload_0_2201;
  wire       [7:0]    _zz_dataOut_payload_0_2202;
  wire                _zz_dataOut_payload_0_2203;
  wire       [7:0]    _zz_dataOut_payload_0_2204;
  wire       [7:0]    _zz_dataOut_payload_0_2205;
  wire                _zz_dataOut_payload_0_2206;
  wire       [7:0]    _zz_dataOut_payload_0_2207;
  wire       [7:0]    _zz_dataOut_payload_0_2208;
  wire                _zz_dataOut_payload_0_2209;
  wire       [7:0]    _zz_dataOut_payload_0_2210;
  wire       [7:0]    _zz_dataOut_payload_0_2211;
  wire                _zz_dataOut_payload_0_2212;
  wire       [7:0]    _zz_dataOut_payload_0_2213;
  wire       [7:0]    _zz_dataOut_payload_0_2214;
  wire                _zz_dataOut_payload_0_2215;
  wire       [7:0]    _zz_dataOut_payload_0_2216;
  wire       [7:0]    _zz_dataOut_payload_0_2217;
  wire                _zz_dataOut_payload_0_2218;
  wire                _zz_dataOut_payload_0_2219;
  reg        [7:0]    _zz_dataOut_payload_0_2220;
  reg        [7:0]    _zz_dataOut_payload_0_2221;
  reg        [7:0]    _zz_dataOut_payload_0_2222;
  reg        [7:0]    _zz_dataOut_payload_0_2223;
  wire                _zz_dataOut_payload_0_2224;
  wire       [7:0]    _zz_dataOut_payload_0_2225;
  wire       [7:0]    _zz_dataOut_payload_0_2226;
  wire                _zz_dataOut_payload_0_2227;
  wire       [7:0]    _zz_dataOut_payload_0_2228;
  wire       [7:0]    _zz_dataOut_payload_0_2229;
  wire                _zz_dataOut_payload_0_2230;
  wire                _zz_dataOut_payload_0_2231;
  reg        [7:0]    _zz_dataOut_payload_0_2232;
  reg        [7:0]    _zz_dataOut_payload_0_2233;
  reg        [7:0]    _zz_dataOut_payload_0_2234;
  reg        [7:0]    _zz_dataOut_payload_0_2235;
  reg        [7:0]    _zz_dataOut_payload_0_2236;
  reg        [7:0]    _zz_dataOut_payload_0_2237;
  reg        [7:0]    _zz_dataOut_payload_0_2238;
  reg        [7:0]    _zz_dataOut_payload_0_2239;
  reg        [7:0]    _zz_dataOut_payload_0_2240;
  reg        [7:0]    _zz_dataOut_payload_0_2241;
  reg        [7:0]    _zz_dataOut_payload_0_2242;
  reg        [7:0]    _zz_dataOut_payload_0_2243;
  wire                _zz_dataOut_payload_0_2244;
  wire       [7:0]    _zz_dataOut_payload_0_2245;
  wire       [7:0]    _zz_dataOut_payload_0_2246;
  wire                _zz_dataOut_payload_0_2247;
  wire       [7:0]    _zz_dataOut_payload_0_2248;
  wire       [7:0]    _zz_dataOut_payload_0_2249;
  wire                _zz_dataOut_payload_0_2250;
  wire       [7:0]    _zz_dataOut_payload_0_2251;
  wire       [7:0]    _zz_dataOut_payload_0_2252;
  wire                _zz_dataOut_payload_0_2253;
  wire       [7:0]    _zz_dataOut_payload_0_2254;
  wire       [7:0]    _zz_dataOut_payload_0_2255;
  wire                _zz_dataOut_payload_0_2256;
  wire       [7:0]    _zz_dataOut_payload_0_2257;
  wire       [7:0]    _zz_dataOut_payload_0_2258;
  wire                _zz_dataOut_payload_0_2259;
  wire       [7:0]    _zz_dataOut_payload_0_2260;
  wire       [7:0]    _zz_dataOut_payload_0_2261;
  wire                _zz_dataOut_payload_0_2262;
  wire                _zz_dataOut_payload_0_2263;
  reg        [7:0]    _zz_dataOut_payload_0_2264;
  reg        [7:0]    _zz_dataOut_payload_0_2265;
  reg        [7:0]    _zz_dataOut_payload_0_2266;
  reg        [7:0]    _zz_dataOut_payload_0_2267;
  wire                _zz_dataOut_payload_0_2268;
  wire       [7:0]    _zz_dataOut_payload_0_2269;
  wire       [7:0]    _zz_dataOut_payload_0_2270;
  wire                _zz_dataOut_payload_0_2271;
  wire       [7:0]    _zz_dataOut_payload_0_2272;
  wire       [7:0]    _zz_dataOut_payload_0_2273;
  wire                _zz_dataOut_payload_0_2274;
  wire                _zz_dataOut_payload_0_2275;
  reg        [7:0]    _zz_dataOut_payload_0_2276;
  reg        [7:0]    _zz_dataOut_payload_0_2277;
  reg        [7:0]    _zz_dataOut_payload_0_2278;
  reg        [7:0]    _zz_dataOut_payload_0_2279;
  reg        [7:0]    _zz_dataOut_payload_0_2280;
  reg        [7:0]    _zz_dataOut_payload_0_2281;
  reg        [7:0]    _zz_dataOut_payload_0_2282;
  reg        [7:0]    _zz_dataOut_payload_0_2283;
  reg        [7:0]    _zz_dataOut_payload_0_2284;
  reg        [7:0]    _zz_dataOut_payload_0_2285;
  reg        [7:0]    _zz_dataOut_payload_0_2286;
  reg        [7:0]    _zz_dataOut_payload_0_2287;
  wire                _zz_dataOut_payload_0_2288;
  wire       [7:0]    _zz_dataOut_payload_0_2289;
  wire       [7:0]    _zz_dataOut_payload_0_2290;
  wire                _zz_dataOut_payload_0_2291;
  wire       [7:0]    _zz_dataOut_payload_0_2292;
  wire       [7:0]    _zz_dataOut_payload_0_2293;
  wire                _zz_dataOut_payload_0_2294;
  wire       [7:0]    _zz_dataOut_payload_0_2295;
  wire       [7:0]    _zz_dataOut_payload_0_2296;
  wire                _zz_dataOut_payload_0_2297;
  wire       [7:0]    _zz_dataOut_payload_0_2298;
  wire       [7:0]    _zz_dataOut_payload_0_2299;
  wire                _zz_dataOut_payload_0_2300;
  wire       [7:0]    _zz_dataOut_payload_0_2301;
  wire       [7:0]    _zz_dataOut_payload_0_2302;
  wire                _zz_dataOut_payload_0_2303;
  wire       [7:0]    _zz_dataOut_payload_0_2304;
  wire       [7:0]    _zz_dataOut_payload_0_2305;
  wire                _zz_dataOut_payload_0_2306;
  wire                _zz_dataOut_payload_0_2307;
  reg        [7:0]    _zz_dataOut_payload_0_2308;
  reg        [7:0]    _zz_dataOut_payload_0_2309;
  reg        [7:0]    _zz_dataOut_payload_0_2310;
  reg        [7:0]    _zz_dataOut_payload_0_2311;
  wire                _zz_dataOut_payload_0_2312;
  wire       [7:0]    _zz_dataOut_payload_0_2313;
  wire       [7:0]    _zz_dataOut_payload_0_2314;
  wire                _zz_dataOut_payload_0_2315;
  wire       [7:0]    _zz_dataOut_payload_0_2316;
  wire       [7:0]    _zz_dataOut_payload_0_2317;
  wire                _zz_dataOut_payload_0_2318;
  wire                _zz_dataOut_payload_0_2319;
  reg        [7:0]    _zz_dataOut_payload_0_2320;
  reg        [7:0]    _zz_dataOut_payload_0_2321;
  reg        [7:0]    _zz_dataOut_payload_0_2322;
  reg        [7:0]    _zz_dataOut_payload_0_2323;
  reg        [7:0]    _zz_dataOut_payload_0_2324;
  reg        [7:0]    _zz_dataOut_payload_0_2325;
  reg        [7:0]    _zz_dataOut_payload_0_2326;
  reg        [7:0]    _zz_dataOut_payload_0_2327;
  reg        [7:0]    _zz_dataOut_payload_0_2328;
  reg        [7:0]    _zz_dataOut_payload_0_2329;
  reg        [7:0]    _zz_dataOut_payload_0_2330;
  reg        [7:0]    _zz_dataOut_payload_0_2331;
  wire                _zz_dataOut_payload_0_2332;
  wire       [7:0]    _zz_dataOut_payload_0_2333;
  wire       [7:0]    _zz_dataOut_payload_0_2334;
  wire                _zz_dataOut_payload_0_2335;
  wire       [7:0]    _zz_dataOut_payload_0_2336;
  wire       [7:0]    _zz_dataOut_payload_0_2337;
  wire                _zz_dataOut_payload_0_2338;
  wire       [7:0]    _zz_dataOut_payload_0_2339;
  wire       [7:0]    _zz_dataOut_payload_0_2340;
  wire                _zz_dataOut_payload_0_2341;
  wire       [7:0]    _zz_dataOut_payload_0_2342;
  wire       [7:0]    _zz_dataOut_payload_0_2343;
  wire                _zz_dataOut_payload_0_2344;
  wire       [7:0]    _zz_dataOut_payload_0_2345;
  wire       [7:0]    _zz_dataOut_payload_0_2346;
  wire                _zz_dataOut_payload_0_2347;
  wire       [7:0]    _zz_dataOut_payload_0_2348;
  wire       [7:0]    _zz_dataOut_payload_0_2349;
  wire                _zz_dataOut_payload_0_2350;
  wire                _zz_dataOut_payload_0_2351;
  reg        [7:0]    _zz_dataOut_payload_0_2352;
  reg        [7:0]    _zz_dataOut_payload_0_2353;
  reg        [7:0]    _zz_dataOut_payload_0_2354;
  reg        [7:0]    _zz_dataOut_payload_0_2355;
  wire                _zz_dataOut_payload_0_2356;
  wire       [7:0]    _zz_dataOut_payload_0_2357;
  wire       [7:0]    _zz_dataOut_payload_0_2358;
  wire                _zz_dataOut_payload_0_2359;
  wire       [7:0]    _zz_dataOut_payload_0_2360;
  wire       [7:0]    _zz_dataOut_payload_0_2361;
  wire                _zz_dataOut_payload_0_2362;
  wire                _zz_dataOut_payload_0_2363;
  reg        [7:0]    _zz_dataOut_payload_0_2364;
  reg        [7:0]    _zz_dataOut_payload_0_2365;
  reg        [7:0]    _zz_dataOut_payload_0_2366;
  reg        [7:0]    _zz_dataOut_payload_0_2367;
  reg        [7:0]    _zz_dataOut_payload_0_2368;
  reg        [7:0]    _zz_dataOut_payload_0_2369;
  reg        [7:0]    _zz_dataOut_payload_0_2370;
  reg        [7:0]    _zz_dataOut_payload_0_2371;
  reg        [7:0]    _zz_dataOut_payload_0_2372;
  reg        [7:0]    _zz_dataOut_payload_0_2373;
  reg        [7:0]    _zz_dataOut_payload_0_2374;
  reg        [7:0]    _zz_dataOut_payload_0_2375;
  wire                _zz_dataOut_payload_0_2376;
  wire       [7:0]    _zz_dataOut_payload_0_2377;
  wire       [7:0]    _zz_dataOut_payload_0_2378;
  wire                _zz_dataOut_payload_0_2379;
  wire       [7:0]    _zz_dataOut_payload_0_2380;
  wire       [7:0]    _zz_dataOut_payload_0_2381;
  wire                _zz_dataOut_payload_0_2382;
  wire       [7:0]    _zz_dataOut_payload_0_2383;
  wire       [7:0]    _zz_dataOut_payload_0_2384;
  wire                _zz_dataOut_payload_0_2385;
  wire       [7:0]    _zz_dataOut_payload_0_2386;
  wire       [7:0]    _zz_dataOut_payload_0_2387;
  wire                _zz_dataOut_payload_0_2388;
  wire       [7:0]    _zz_dataOut_payload_0_2389;
  wire       [7:0]    _zz_dataOut_payload_0_2390;
  wire                _zz_dataOut_payload_0_2391;
  wire       [7:0]    _zz_dataOut_payload_0_2392;
  wire       [7:0]    _zz_dataOut_payload_0_2393;
  wire                _zz_dataOut_payload_0_2394;
  wire                _zz_dataOut_payload_0_2395;
  reg        [7:0]    _zz_dataOut_payload_0_2396;
  reg        [7:0]    _zz_dataOut_payload_0_2397;
  reg        [7:0]    _zz_dataOut_payload_0_2398;
  reg        [7:0]    _zz_dataOut_payload_0_2399;
  wire                _zz_dataOut_payload_0_2400;
  wire       [7:0]    _zz_dataOut_payload_0_2401;
  wire       [7:0]    _zz_dataOut_payload_0_2402;
  wire                _zz_dataOut_payload_0_2403;
  wire       [7:0]    _zz_dataOut_payload_0_2404;
  wire       [7:0]    _zz_dataOut_payload_0_2405;
  wire                _zz_dataOut_payload_0_2406;
  wire                _zz_dataOut_payload_0_2407;
  reg        [7:0]    _zz_dataOut_payload_0_2408;
  reg        [7:0]    _zz_dataOut_payload_0_2409;
  reg        [7:0]    _zz_dataOut_payload_0_2410;
  reg        [7:0]    _zz_dataOut_payload_0_2411;
  reg        [7:0]    _zz_dataOut_payload_0_2412;
  reg        [7:0]    _zz_dataOut_payload_0_2413;
  reg        [7:0]    _zz_dataOut_payload_0_2414;
  reg        [7:0]    _zz_dataOut_payload_0_2415;
  reg        [7:0]    _zz_dataOut_payload_0_2416;
  reg        [7:0]    _zz_dataOut_payload_0_2417;
  reg        [7:0]    _zz_dataOut_payload_0_2418;
  reg        [7:0]    _zz_dataOut_payload_0_2419;
  wire                _zz_dataOut_payload_0_2420;
  wire       [7:0]    _zz_dataOut_payload_0_2421;
  wire       [7:0]    _zz_dataOut_payload_0_2422;
  wire                _zz_dataOut_payload_0_2423;
  wire       [7:0]    _zz_dataOut_payload_0_2424;
  wire       [7:0]    _zz_dataOut_payload_0_2425;
  wire                _zz_dataOut_payload_0_2426;
  wire       [7:0]    _zz_dataOut_payload_0_2427;
  wire       [7:0]    _zz_dataOut_payload_0_2428;
  wire                _zz_dataOut_payload_0_2429;
  wire       [7:0]    _zz_dataOut_payload_0_2430;
  wire       [7:0]    _zz_dataOut_payload_0_2431;
  wire                _zz_dataOut_payload_0_2432;
  wire       [7:0]    _zz_dataOut_payload_0_2433;
  wire       [7:0]    _zz_dataOut_payload_0_2434;
  wire                _zz_dataOut_payload_0_2435;
  wire       [7:0]    _zz_dataOut_payload_0_2436;
  wire       [7:0]    _zz_dataOut_payload_0_2437;
  wire                _zz_dataOut_payload_0_2438;
  wire                _zz_dataOut_payload_0_2439;
  reg        [7:0]    _zz_dataOut_payload_0_2440;
  reg        [7:0]    _zz_dataOut_payload_0_2441;
  reg        [7:0]    _zz_dataOut_payload_0_2442;
  reg        [7:0]    _zz_dataOut_payload_0_2443;
  wire                _zz_dataOut_payload_0_2444;
  wire       [7:0]    _zz_dataOut_payload_0_2445;
  wire       [7:0]    _zz_dataOut_payload_0_2446;
  wire                _zz_dataOut_payload_0_2447;
  wire       [7:0]    _zz_dataOut_payload_0_2448;
  wire       [7:0]    _zz_dataOut_payload_0_2449;
  wire                _zz_dataOut_payload_0_2450;
  wire                _zz_dataOut_payload_0_2451;
  reg        [7:0]    _zz_dataOut_payload_0_2452;
  reg        [7:0]    _zz_dataOut_payload_0_2453;
  reg        [7:0]    _zz_dataOut_payload_0_2454;
  reg        [7:0]    _zz_dataOut_payload_0_2455;
  reg        [7:0]    _zz_dataOut_payload_0_2456;
  reg        [7:0]    _zz_dataOut_payload_0_2457;
  reg        [7:0]    _zz_dataOut_payload_0_2458;
  reg        [7:0]    _zz_dataOut_payload_0_2459;
  reg        [7:0]    _zz_dataOut_payload_0_2460;
  reg        [7:0]    _zz_dataOut_payload_0_2461;
  reg        [7:0]    _zz_dataOut_payload_0_2462;
  reg        [7:0]    _zz_dataOut_payload_0_2463;
  wire                _zz_dataOut_payload_0_2464;
  wire       [7:0]    _zz_dataOut_payload_0_2465;
  wire       [7:0]    _zz_dataOut_payload_0_2466;
  wire                _zz_dataOut_payload_0_2467;
  wire       [7:0]    _zz_dataOut_payload_0_2468;
  wire       [7:0]    _zz_dataOut_payload_0_2469;
  wire                _zz_dataOut_payload_0_2470;
  wire       [7:0]    _zz_dataOut_payload_0_2471;
  wire       [7:0]    _zz_dataOut_payload_0_2472;
  wire                _zz_dataOut_payload_0_2473;
  wire       [7:0]    _zz_dataOut_payload_0_2474;
  wire       [7:0]    _zz_dataOut_payload_0_2475;
  wire                _zz_dataOut_payload_0_2476;
  wire       [7:0]    _zz_dataOut_payload_0_2477;
  wire       [7:0]    _zz_dataOut_payload_0_2478;
  wire                _zz_dataOut_payload_0_2479;
  wire       [7:0]    _zz_dataOut_payload_0_2480;
  wire       [7:0]    _zz_dataOut_payload_0_2481;
  wire                _zz_dataOut_payload_0_2482;
  wire                _zz_dataOut_payload_0_2483;
  reg        [7:0]    _zz_dataOut_payload_0_2484;
  reg        [7:0]    _zz_dataOut_payload_0_2485;
  reg        [7:0]    _zz_dataOut_payload_0_2486;
  reg        [7:0]    _zz_dataOut_payload_0_2487;
  wire                _zz_dataOut_payload_0_2488;
  wire       [7:0]    _zz_dataOut_payload_0_2489;
  wire       [7:0]    _zz_dataOut_payload_0_2490;
  wire                _zz_dataOut_payload_0_2491;
  wire       [7:0]    _zz_dataOut_payload_0_2492;
  wire       [7:0]    _zz_dataOut_payload_0_2493;
  wire                _zz_dataOut_payload_0_2494;
  wire                _zz_dataOut_payload_0_2495;
  reg        [7:0]    _zz_dataOut_payload_0_2496;
  reg        [7:0]    _zz_dataOut_payload_0_2497;
  reg        [7:0]    _zz_dataOut_payload_0_2498;
  reg        [7:0]    _zz_dataOut_payload_0_2499;
  reg        [7:0]    _zz_dataOut_payload_0_2500;
  reg        [7:0]    _zz_dataOut_payload_0_2501;
  reg        [7:0]    _zz_dataOut_payload_0_2502;
  reg        [7:0]    _zz_dataOut_payload_0_2503;
  reg        [7:0]    _zz_dataOut_payload_0_2504;
  reg        [7:0]    _zz_dataOut_payload_0_2505;
  reg        [7:0]    _zz_dataOut_payload_0_2506;
  reg        [7:0]    _zz_dataOut_payload_0_2507;
  wire                _zz_dataOut_payload_0_2508;
  wire       [7:0]    _zz_dataOut_payload_0_2509;
  wire       [7:0]    _zz_dataOut_payload_0_2510;
  wire                _zz_dataOut_payload_0_2511;
  wire       [7:0]    _zz_dataOut_payload_0_2512;
  wire       [7:0]    _zz_dataOut_payload_0_2513;
  wire                _zz_dataOut_payload_0_2514;
  wire       [7:0]    _zz_dataOut_payload_0_2515;
  wire       [7:0]    _zz_dataOut_payload_0_2516;
  wire                _zz_dataOut_payload_0_2517;
  wire       [7:0]    _zz_dataOut_payload_0_2518;
  wire       [7:0]    _zz_dataOut_payload_0_2519;
  wire                _zz_dataOut_payload_0_2520;
  wire       [7:0]    _zz_dataOut_payload_0_2521;
  wire       [7:0]    _zz_dataOut_payload_0_2522;
  wire                _zz_dataOut_payload_0_2523;
  wire       [7:0]    _zz_dataOut_payload_0_2524;
  wire       [7:0]    _zz_dataOut_payload_0_2525;
  wire                _zz_dataOut_payload_0_2526;
  wire                _zz_dataOut_payload_0_2527;
  reg        [7:0]    _zz_dataOut_payload_0_2528;
  reg        [7:0]    _zz_dataOut_payload_0_2529;
  reg        [7:0]    _zz_dataOut_payload_0_2530;
  reg        [7:0]    _zz_dataOut_payload_0_2531;
  wire                _zz_dataOut_payload_0_2532;
  wire       [7:0]    _zz_dataOut_payload_0_2533;
  wire       [7:0]    _zz_dataOut_payload_0_2534;
  wire                _zz_dataOut_payload_0_2535;
  wire       [7:0]    _zz_dataOut_payload_0_2536;
  wire       [7:0]    _zz_dataOut_payload_0_2537;
  wire                _zz_dataOut_payload_0_2538;
  wire                _zz_dataOut_payload_0_2539;
  reg        [7:0]    _zz_dataOut_payload_0_2540;
  reg        [7:0]    _zz_dataOut_payload_0_2541;
  reg        [7:0]    _zz_dataOut_payload_0_2542;
  reg        [7:0]    _zz_dataOut_payload_0_2543;
  reg        [7:0]    _zz_dataOut_payload_0_2544;
  reg        [7:0]    _zz_dataOut_payload_0_2545;
  reg        [7:0]    _zz_dataOut_payload_0_2546;
  reg        [7:0]    _zz_dataOut_payload_0_2547;
  reg        [7:0]    _zz_dataOut_payload_0_2548;
  reg        [7:0]    _zz_dataOut_payload_0_2549;
  reg        [7:0]    _zz_dataOut_payload_0_2550;
  reg        [7:0]    _zz_dataOut_payload_0_2551;
  wire                _zz_dataOut_payload_0_2552;
  wire       [7:0]    _zz_dataOut_payload_0_2553;
  wire       [7:0]    _zz_dataOut_payload_0_2554;
  wire                _zz_dataOut_payload_0_2555;
  wire       [7:0]    _zz_dataOut_payload_0_2556;
  wire       [7:0]    _zz_dataOut_payload_0_2557;
  wire                _zz_dataOut_payload_0_2558;
  wire       [7:0]    _zz_dataOut_payload_0_2559;
  wire       [7:0]    _zz_dataOut_payload_0_2560;
  wire                _zz_dataOut_payload_0_2561;
  wire       [7:0]    _zz_dataOut_payload_0_2562;
  wire       [7:0]    _zz_dataOut_payload_0_2563;
  wire                _zz_dataOut_payload_0_2564;
  wire       [7:0]    _zz_dataOut_payload_0_2565;
  wire       [7:0]    _zz_dataOut_payload_0_2566;
  wire                _zz_dataOut_payload_0_2567;
  wire       [7:0]    _zz_dataOut_payload_0_2568;
  wire       [7:0]    _zz_dataOut_payload_0_2569;
  wire                _zz_dataOut_payload_0_2570;
  wire                _zz_dataOut_payload_0_2571;
  reg        [7:0]    _zz_dataOut_payload_0_2572;
  reg        [7:0]    _zz_dataOut_payload_0_2573;
  reg        [7:0]    _zz_dataOut_payload_0_2574;
  reg        [7:0]    _zz_dataOut_payload_0_2575;
  wire                _zz_dataOut_payload_0_2576;
  wire       [7:0]    _zz_dataOut_payload_0_2577;
  wire       [7:0]    _zz_dataOut_payload_0_2578;
  wire                _zz_dataOut_payload_0_2579;
  wire       [7:0]    _zz_dataOut_payload_0_2580;
  wire       [7:0]    _zz_dataOut_payload_0_2581;
  wire                _zz_dataOut_payload_0_2582;
  wire                _zz_dataOut_payload_0_2583;
  reg        [7:0]    _zz_dataOut_payload_0_2584;
  reg        [7:0]    _zz_dataOut_payload_0_2585;
  reg        [7:0]    _zz_dataOut_payload_0_2586;
  reg        [7:0]    _zz_dataOut_payload_0_2587;
  reg        [7:0]    _zz_dataOut_payload_0_2588;
  reg        [7:0]    _zz_dataOut_payload_0_2589;
  reg        [7:0]    _zz_dataOut_payload_0_2590;
  reg        [7:0]    _zz_dataOut_payload_0_2591;
  reg        [7:0]    _zz_dataOut_payload_0_2592;
  reg        [7:0]    _zz_dataOut_payload_0_2593;
  reg        [7:0]    _zz_dataOut_payload_0_2594;
  reg        [7:0]    _zz_dataOut_payload_0_2595;
  wire                _zz_dataOut_payload_0_2596;
  wire       [7:0]    _zz_dataOut_payload_0_2597;
  wire       [7:0]    _zz_dataOut_payload_0_2598;
  wire                _zz_dataOut_payload_0_2599;
  wire       [7:0]    _zz_dataOut_payload_0_2600;
  wire       [7:0]    _zz_dataOut_payload_0_2601;
  wire                _zz_dataOut_payload_0_2602;
  wire       [7:0]    _zz_dataOut_payload_0_2603;
  wire       [7:0]    _zz_dataOut_payload_0_2604;
  wire                _zz_dataOut_payload_0_2605;
  wire       [7:0]    _zz_dataOut_payload_0_2606;
  wire       [7:0]    _zz_dataOut_payload_0_2607;
  wire                _zz_dataOut_payload_0_2608;
  wire       [7:0]    _zz_dataOut_payload_0_2609;
  wire       [7:0]    _zz_dataOut_payload_0_2610;
  wire                _zz_dataOut_payload_0_2611;
  wire       [7:0]    _zz_dataOut_payload_0_2612;
  wire       [7:0]    _zz_dataOut_payload_0_2613;
  wire                _zz_dataOut_payload_0_2614;
  wire                _zz_dataOut_payload_0_2615;
  reg        [7:0]    _zz_dataOut_payload_0_2616;
  reg        [7:0]    _zz_dataOut_payload_0_2617;
  reg        [7:0]    _zz_dataOut_payload_0_2618;
  reg        [7:0]    _zz_dataOut_payload_0_2619;
  wire                _zz_dataOut_payload_0_2620;
  wire       [7:0]    _zz_dataOut_payload_0_2621;
  wire       [7:0]    _zz_dataOut_payload_0_2622;
  wire                _zz_dataOut_payload_0_2623;
  wire       [7:0]    _zz_dataOut_payload_0_2624;
  wire       [7:0]    _zz_dataOut_payload_0_2625;
  wire                _zz_dataOut_payload_0_2626;
  wire                _zz_dataOut_payload_0_2627;
  reg        [7:0]    _zz_dataOut_payload_0_2628;
  reg        [7:0]    _zz_dataOut_payload_0_2629;
  reg        [7:0]    _zz_dataOut_payload_0_2630;
  reg        [7:0]    _zz_dataOut_payload_0_2631;
  reg        [7:0]    _zz_dataOut_payload_0_2632;
  reg        [7:0]    _zz_dataOut_payload_0_2633;
  reg        [7:0]    _zz_dataOut_payload_0_2634;
  reg        [7:0]    _zz_dataOut_payload_0_2635;
  reg        [7:0]    _zz_dataOut_payload_0_2636;
  reg        [7:0]    _zz_dataOut_payload_0_2637;
  reg        [7:0]    _zz_dataOut_payload_0_2638;
  reg        [7:0]    _zz_dataOut_payload_0_2639;
  wire                _zz_dataOut_payload_0_2640;
  wire       [7:0]    _zz_dataOut_payload_0_2641;
  wire       [7:0]    _zz_dataOut_payload_0_2642;
  wire                _zz_dataOut_payload_0_2643;
  wire       [7:0]    _zz_dataOut_payload_0_2644;
  wire       [7:0]    _zz_dataOut_payload_0_2645;
  wire                _zz_dataOut_payload_0_2646;
  wire       [7:0]    _zz_dataOut_payload_0_2647;
  wire       [7:0]    _zz_dataOut_payload_0_2648;
  wire                _zz_dataOut_payload_0_2649;
  wire       [7:0]    _zz_dataOut_payload_0_2650;
  wire       [7:0]    _zz_dataOut_payload_0_2651;
  wire                _zz_dataOut_payload_0_2652;
  wire       [7:0]    _zz_dataOut_payload_0_2653;
  wire       [7:0]    _zz_dataOut_payload_0_2654;
  wire                _zz_dataOut_payload_0_2655;
  wire       [7:0]    _zz_dataOut_payload_0_2656;
  wire       [7:0]    _zz_dataOut_payload_0_2657;
  wire                _zz_dataOut_payload_0_2658;
  wire                _zz_dataOut_payload_0_2659;
  reg        [7:0]    _zz_dataOut_payload_0_2660;
  reg        [7:0]    _zz_dataOut_payload_0_2661;
  reg        [7:0]    _zz_dataOut_payload_0_2662;
  reg        [7:0]    _zz_dataOut_payload_0_2663;
  wire                _zz_dataOut_payload_0_2664;
  wire       [7:0]    _zz_dataOut_payload_0_2665;
  wire       [7:0]    _zz_dataOut_payload_0_2666;
  wire                _zz_dataOut_payload_0_2667;
  wire       [7:0]    _zz_dataOut_payload_0_2668;
  wire       [7:0]    _zz_dataOut_payload_0_2669;
  wire                _zz_dataOut_payload_0_2670;
  wire                _zz_dataOut_payload_0_2671;
  reg        [7:0]    _zz_dataOut_payload_0_2672;
  reg        [7:0]    _zz_dataOut_payload_0_2673;
  reg        [7:0]    _zz_dataOut_payload_0_2674;
  reg        [7:0]    _zz_dataOut_payload_0_2675;
  reg        [7:0]    _zz_dataOut_payload_0_2676;
  reg        [7:0]    _zz_dataOut_payload_0_2677;
  reg        [7:0]    _zz_dataOut_payload_0_2678;
  reg        [7:0]    _zz_dataOut_payload_0_2679;
  reg        [7:0]    _zz_dataOut_payload_0_2680;
  reg        [7:0]    _zz_dataOut_payload_0_2681;
  reg        [7:0]    _zz_dataOut_payload_0_2682;
  reg        [7:0]    _zz_dataOut_payload_0_2683;
  wire                _zz_dataOut_payload_0_2684;
  wire       [7:0]    _zz_dataOut_payload_0_2685;
  wire       [7:0]    _zz_dataOut_payload_0_2686;
  wire                _zz_dataOut_payload_0_2687;
  wire       [7:0]    _zz_dataOut_payload_0_2688;
  wire       [7:0]    _zz_dataOut_payload_0_2689;
  wire                _zz_dataOut_payload_0_2690;
  wire       [7:0]    _zz_dataOut_payload_0_2691;
  wire       [7:0]    _zz_dataOut_payload_0_2692;
  wire                _zz_dataOut_payload_0_2693;
  wire       [7:0]    _zz_dataOut_payload_0_2694;
  wire       [7:0]    _zz_dataOut_payload_0_2695;
  wire                _zz_dataOut_payload_0_2696;
  wire       [7:0]    _zz_dataOut_payload_0_2697;
  wire       [7:0]    _zz_dataOut_payload_0_2698;
  wire                _zz_dataOut_payload_0_2699;
  wire       [7:0]    _zz_dataOut_payload_0_2700;
  wire       [7:0]    _zz_dataOut_payload_0_2701;
  wire                _zz_dataOut_payload_0_2702;
  wire                _zz_dataOut_payload_0_2703;
  reg        [7:0]    _zz_dataOut_payload_0_2704;
  reg        [7:0]    _zz_dataOut_payload_0_2705;
  reg        [7:0]    _zz_dataOut_payload_0_2706;
  reg        [7:0]    _zz_dataOut_payload_0_2707;
  wire                _zz_dataOut_payload_0_2708;
  wire       [7:0]    _zz_dataOut_payload_0_2709;
  wire       [7:0]    _zz_dataOut_payload_0_2710;
  wire                _zz_dataOut_payload_0_2711;
  wire       [7:0]    _zz_dataOut_payload_0_2712;
  wire       [7:0]    _zz_dataOut_payload_0_2713;
  wire                _zz_dataOut_payload_0_2714;
  wire                _zz_dataOut_payload_0_2715;
  reg        [7:0]    _zz_dataOut_payload_0_2716;
  reg        [7:0]    _zz_dataOut_payload_0_2717;
  reg        [7:0]    _zz_dataOut_payload_0_2718;
  reg        [7:0]    _zz_dataOut_payload_0_2719;
  reg        [7:0]    _zz_dataOut_payload_0_2720;
  reg        [7:0]    _zz_dataOut_payload_0_2721;
  reg        [7:0]    _zz_dataOut_payload_0_2722;
  reg        [7:0]    _zz_dataOut_payload_0_2723;
  reg        [7:0]    _zz_dataOut_payload_0_2724;
  reg        [7:0]    _zz_dataOut_payload_0_2725;
  reg        [7:0]    _zz_dataOut_payload_0_2726;
  reg        [7:0]    _zz_dataOut_payload_0_2727;
  wire                _zz_dataOut_payload_0_2728;
  wire       [7:0]    _zz_dataOut_payload_0_2729;
  wire       [7:0]    _zz_dataOut_payload_0_2730;
  wire                _zz_dataOut_payload_0_2731;
  wire       [7:0]    _zz_dataOut_payload_0_2732;
  wire       [7:0]    _zz_dataOut_payload_0_2733;
  wire                _zz_dataOut_payload_0_2734;
  wire       [7:0]    _zz_dataOut_payload_0_2735;
  wire       [7:0]    _zz_dataOut_payload_0_2736;
  wire                _zz_dataOut_payload_0_2737;
  wire       [7:0]    _zz_dataOut_payload_0_2738;
  wire       [7:0]    _zz_dataOut_payload_0_2739;
  wire                _zz_dataOut_payload_0_2740;
  wire       [7:0]    _zz_dataOut_payload_0_2741;
  wire       [7:0]    _zz_dataOut_payload_0_2742;
  wire                _zz_dataOut_payload_0_2743;
  wire       [7:0]    _zz_dataOut_payload_0_2744;
  wire       [7:0]    _zz_dataOut_payload_0_2745;
  wire                _zz_dataOut_payload_0_2746;
  wire                _zz_dataOut_payload_0_2747;
  reg        [7:0]    _zz_dataOut_payload_0_2748;
  reg        [7:0]    _zz_dataOut_payload_0_2749;
  reg        [7:0]    _zz_dataOut_payload_0_2750;
  reg        [7:0]    _zz_dataOut_payload_0_2751;
  wire                _zz_dataOut_payload_0_2752;
  wire       [7:0]    _zz_dataOut_payload_0_2753;
  wire       [7:0]    _zz_dataOut_payload_0_2754;
  wire                _zz_dataOut_payload_0_2755;
  wire       [7:0]    _zz_dataOut_payload_0_2756;
  wire       [7:0]    _zz_dataOut_payload_0_2757;
  wire                _zz_dataOut_payload_0_2758;
  wire                _zz_dataOut_payload_0_2759;
  reg        [7:0]    _zz_dataOut_payload_0_2760;
  reg        [7:0]    _zz_dataOut_payload_0_2761;
  reg        [7:0]    _zz_dataOut_payload_0_2762;
  reg        [7:0]    _zz_dataOut_payload_0_2763;
  reg        [7:0]    _zz_dataOut_payload_0_2764;
  reg        [7:0]    _zz_dataOut_payload_0_2765;
  reg        [7:0]    _zz_dataOut_payload_0_2766;
  reg        [7:0]    _zz_dataOut_payload_0_2767;
  reg        [7:0]    _zz_dataOut_payload_0_2768;
  reg        [7:0]    _zz_dataOut_payload_0_2769;
  reg        [7:0]    _zz_dataOut_payload_0_2770;
  reg        [7:0]    _zz_dataOut_payload_0_2771;
  wire                _zz_dataOut_payload_0_2772;
  wire       [7:0]    _zz_dataOut_payload_0_2773;
  wire       [7:0]    _zz_dataOut_payload_0_2774;
  wire                _zz_dataOut_payload_0_2775;
  wire       [7:0]    _zz_dataOut_payload_0_2776;
  wire       [7:0]    _zz_dataOut_payload_0_2777;
  wire                _zz_dataOut_payload_0_2778;
  wire       [7:0]    _zz_dataOut_payload_0_2779;
  wire       [7:0]    _zz_dataOut_payload_0_2780;
  wire                _zz_dataOut_payload_0_2781;
  wire       [7:0]    _zz_dataOut_payload_0_2782;
  wire       [7:0]    _zz_dataOut_payload_0_2783;
  wire                _zz_dataOut_payload_0_2784;
  wire       [7:0]    _zz_dataOut_payload_0_2785;
  wire       [7:0]    _zz_dataOut_payload_0_2786;
  wire                _zz_dataOut_payload_0_2787;
  wire       [7:0]    _zz_dataOut_payload_0_2788;
  wire       [7:0]    _zz_dataOut_payload_0_2789;
  wire                _zz_dataOut_payload_0_2790;
  wire                _zz_dataOut_payload_0_2791;
  reg        [7:0]    _zz_dataOut_payload_0_2792;
  reg        [7:0]    _zz_dataOut_payload_0_2793;
  reg        [7:0]    _zz_dataOut_payload_0_2794;
  reg        [7:0]    _zz_dataOut_payload_0_2795;
  wire                _zz_dataOut_payload_0_2796;
  wire       [7:0]    _zz_dataOut_payload_0_2797;
  wire       [7:0]    _zz_dataOut_payload_0_2798;
  wire                _zz_dataOut_payload_0_2799;
  wire       [7:0]    _zz_dataOut_payload_0_2800;
  wire       [7:0]    _zz_dataOut_payload_0_2801;
  wire                _zz_dataOut_payload_0_2802;
  wire                _zz_dataOut_payload_0_2803;
  reg        [7:0]    _zz_dataOut_payload_0_2804;
  reg        [7:0]    _zz_dataOut_payload_0_2805;
  reg        [7:0]    _zz_dataOut_payload_0_2806;
  reg        [7:0]    _zz_dataOut_payload_0_2807;
  reg        [7:0]    _zz_dataOut_payload_0_2808;
  reg        [7:0]    _zz_dataOut_payload_0_2809;
  reg        [7:0]    _zz_dataOut_payload_0_2810;
  reg        [7:0]    _zz_dataOut_payload_0_2811;
  reg        [7:0]    _zz_dataOut_payload_0_2812;
  reg        [7:0]    _zz_dataOut_payload_0_2813;
  reg        [7:0]    _zz_dataOut_payload_0_2814;
  reg        [7:0]    _zz_dataOut_payload_0_2815;
  reg        [7:0]    _zz_dataOut_payload_0_2816;
  reg        [7:0]    _zz_dataOut_payload_0_2817;
  reg        [7:0]    _zz_dataOut_payload_0_2818;
  reg        [7:0]    _zz_dataOut_payload_0_2819;
  reg        [7:0]    _zz_dataOut_payload_0_2820;
  reg        [7:0]    _zz_dataOut_payload_0_2821;
  reg        [7:0]    _zz_dataOut_payload_0_2822;
  reg        [7:0]    _zz_dataOut_payload_0_2823;
  reg        [7:0]    _zz_dataOut_payload_0_2824;
  reg        [7:0]    _zz_dataOut_payload_0_2825;
  reg        [7:0]    _zz_dataOut_payload_0_2826;
  reg        [7:0]    _zz_dataOut_payload_0_2827;
  reg        [7:0]    _zz_dataOut_payload_0_2828;
  reg        [7:0]    _zz_dataOut_payload_0_2829;
  reg        [7:0]    _zz_dataOut_payload_0_2830;
  reg        [7:0]    _zz_dataOut_payload_0_2831;
  reg        [7:0]    _zz_dataOut_payload_0_2832;
  reg        [7:0]    _zz_dataOut_payload_0_2833;
  reg        [7:0]    _zz_dataOut_payload_0_2834;
  reg        [7:0]    _zz_dataOut_payload_0_2835;
  reg        [7:0]    _zz_dataOut_payload_0_2836;
  reg        [7:0]    _zz_dataOut_payload_0_2837;
  reg        [7:0]    _zz_dataOut_payload_0_2838;
  reg        [7:0]    _zz_dataOut_payload_0_2839;
  reg        [7:0]    _zz_dataOut_payload_0_2840;
  reg        [7:0]    _zz_dataOut_payload_0_2841;
  reg        [7:0]    _zz_dataOut_payload_0_2842;
  reg        [7:0]    _zz_dataOut_payload_0_2843;
  reg        [7:0]    _zz_dataOut_payload_0_2844;
  reg        [7:0]    _zz_dataOut_payload_0_2845;
  reg        [7:0]    _zz_dataOut_payload_0_2846;
  reg        [7:0]    _zz_dataOut_payload_0_2847;
  reg        [7:0]    _zz_dataOut_payload_0_2848;
  reg        [7:0]    _zz_dataOut_payload_0_2849;
  reg        [7:0]    _zz_dataOut_payload_0_2850;
  reg        [7:0]    _zz_dataOut_payload_0_2851;
  reg        [7:0]    _zz_dataOut_payload_0_2852;
  reg        [7:0]    _zz_dataOut_payload_0_2853;
  reg        [7:0]    _zz_dataOut_payload_0_2854;
  reg        [7:0]    _zz_dataOut_payload_0_2855;
  reg        [7:0]    _zz_dataOut_payload_0_2856;
  reg        [7:0]    _zz_dataOut_payload_0_2857;
  reg        [7:0]    _zz_dataOut_payload_0_2858;
  reg        [7:0]    _zz_dataOut_payload_0_2859;
  reg        [7:0]    _zz_dataOut_payload_0_2860;
  reg        [7:0]    _zz_dataOut_payload_0_2861;
  reg        [7:0]    _zz_dataOut_payload_0_2862;
  reg        [7:0]    _zz_dataOut_payload_0_2863;
  reg        [7:0]    _zz_dataOut_payload_0_2864;
  reg        [7:0]    _zz_dataOut_payload_0_2865;
  reg        [7:0]    _zz_dataOut_payload_0_2866;
  reg        [7:0]    _zz_dataOut_payload_0_2867;
  reg        [7:0]    _zz_dataOut_payload_0_2868;
  reg        [7:0]    _zz_dataOut_payload_0_2869;
  reg        [7:0]    _zz_dataOut_payload_0_2870;
  reg        [7:0]    _zz_dataOut_payload_0_2871;
  reg        [7:0]    _zz_dataOut_payload_0_2872;
  reg        [7:0]    _zz_dataOut_payload_0_2873;
  reg        [7:0]    _zz_dataOut_payload_0_2874;
  reg        [7:0]    _zz_dataOut_payload_0_2875;
  reg        [7:0]    _zz_dataOut_payload_0_2876;
  reg        [7:0]    _zz_dataOut_payload_0_2877;
  reg        [7:0]    _zz_dataOut_payload_0_2878;
  reg        [7:0]    _zz_dataOut_payload_0_2879;
  reg        [7:0]    _zz_dataOut_payload_0_2880;
  reg        [7:0]    _zz_dataOut_payload_0_2881;
  reg        [7:0]    _zz_dataOut_payload_0_2882;
  reg        [7:0]    _zz_dataOut_payload_0_2883;
  reg        [7:0]    _zz_dataOut_payload_0_2884;
  reg        [7:0]    _zz_dataOut_payload_0_2885;
  reg        [7:0]    _zz_dataOut_payload_0_2886;
  reg        [7:0]    _zz_dataOut_payload_0_2887;
  reg        [7:0]    _zz_dataOut_payload_0_2888;
  reg        [7:0]    _zz_dataOut_payload_0_2889;
  reg        [7:0]    _zz_dataOut_payload_0_2890;
  reg        [7:0]    _zz_dataOut_payload_0_2891;
  reg        [7:0]    _zz_dataOut_payload_0_2892;
  reg        [7:0]    _zz_dataOut_payload_0_2893;
  reg        [7:0]    _zz_dataOut_payload_0_2894;
  reg        [7:0]    _zz_dataOut_payload_0_2895;
  reg        [7:0]    _zz_dataOut_payload_0_2896;
  reg        [7:0]    _zz_dataOut_payload_0_2897;
  reg        [7:0]    _zz_dataOut_payload_0_2898;
  reg        [7:0]    _zz_dataOut_payload_0_2899;
  reg        [7:0]    _zz_dataOut_payload_0_2900;
  reg        [7:0]    _zz_dataOut_payload_0_2901;
  reg        [7:0]    _zz_dataOut_payload_0_2902;
  reg        [7:0]    _zz_dataOut_payload_0_2903;
  reg        [7:0]    _zz_dataOut_payload_0_2904;
  reg        [7:0]    _zz_dataOut_payload_0_2905;
  reg        [7:0]    _zz_dataOut_payload_0_2906;
  reg        [7:0]    _zz_dataOut_payload_0_2907;
  reg        [7:0]    _zz_dataOut_payload_0_2908;
  reg        [7:0]    _zz_dataOut_payload_0_2909;
  reg        [7:0]    _zz_dataOut_payload_0_2910;
  reg        [7:0]    _zz_dataOut_payload_0_2911;
  reg        [7:0]    _zz_dataOut_payload_0_2912;
  reg        [7:0]    _zz_dataOut_payload_0_2913;
  reg        [7:0]    _zz_dataOut_payload_0_2914;
  reg        [7:0]    _zz_dataOut_payload_0_2915;
  reg        [7:0]    _zz_dataOut_payload_0_2916;
  reg        [7:0]    _zz_dataOut_payload_0_2917;
  reg        [7:0]    _zz_dataOut_payload_0_2918;
  reg        [7:0]    _zz_dataOut_payload_0_2919;
  reg        [7:0]    _zz_dataOut_payload_0_2920;
  reg        [7:0]    _zz_dataOut_payload_0_2921;
  reg        [7:0]    _zz_dataOut_payload_0_2922;
  reg        [7:0]    _zz_dataOut_payload_0_2923;
  reg        [7:0]    _zz_dataOut_payload_0_2924;
  reg        [7:0]    _zz_dataOut_payload_0_2925;
  reg        [7:0]    _zz_dataOut_payload_0_2926;
  reg        [7:0]    _zz_dataOut_payload_0_2927;
  reg        [7:0]    _zz_dataOut_payload_0_2928;
  reg        [7:0]    _zz_dataOut_payload_0_2929;
  reg        [7:0]    _zz_dataOut_payload_0_2930;
  reg        [7:0]    _zz_dataOut_payload_0_2931;
  reg        [7:0]    _zz_dataOut_payload_0_2932;
  reg        [7:0]    _zz_dataOut_payload_0_2933;
  reg        [7:0]    _zz_dataOut_payload_0_2934;
  reg        [7:0]    _zz_dataOut_payload_0_2935;
  reg        [7:0]    _zz_dataOut_payload_0_2936;
  reg        [7:0]    _zz_dataOut_payload_0_2937;
  reg        [7:0]    _zz_dataOut_payload_0_2938;
  reg        [7:0]    _zz_dataOut_payload_0_2939;
  reg        [7:0]    _zz_dataOut_payload_0_2940;
  reg        [7:0]    _zz_dataOut_payload_0_2941;
  reg        [7:0]    _zz_dataOut_payload_0_2942;
  reg        [7:0]    _zz_dataOut_payload_0_2943;
  reg        [7:0]    _zz_dataOut_payload_0_2944;
  reg        [7:0]    _zz_dataOut_payload_0_2945;
  reg        [7:0]    _zz_dataOut_payload_0_2946;
  reg        [7:0]    _zz_dataOut_payload_0_2947;
  reg        [7:0]    _zz_dataOut_payload_0_2948;
  reg        [7:0]    _zz_dataOut_payload_0_2949;
  reg        [7:0]    _zz_dataOut_payload_0_2950;
  reg        [7:0]    _zz_dataOut_payload_0_2951;
  reg        [7:0]    _zz_dataOut_payload_0_2952;
  reg        [7:0]    _zz_dataOut_payload_0_2953;
  reg        [7:0]    _zz_dataOut_payload_0_2954;
  reg        [7:0]    _zz_dataOut_payload_0_2955;
  reg        [7:0]    _zz_dataOut_payload_0_2956;
  reg        [7:0]    _zz_dataOut_payload_0_2957;
  reg        [7:0]    _zz_dataOut_payload_0_2958;
  reg        [7:0]    _zz_dataOut_payload_0_2959;
  reg        [7:0]    _zz_dataOut_payload_0_2960;
  reg        [7:0]    _zz_dataOut_payload_0_2961;
  reg        [7:0]    _zz_dataOut_payload_0_2962;
  reg        [7:0]    _zz_dataOut_payload_0_2963;
  reg        [7:0]    _zz_dataOut_payload_0_2964;
  reg        [7:0]    _zz_dataOut_payload_0_2965;
  reg        [7:0]    _zz_dataOut_payload_0_2966;
  reg        [7:0]    _zz_dataOut_payload_0_2967;
  reg        [7:0]    _zz_dataOut_payload_0_2968;
  reg        [7:0]    _zz_dataOut_payload_0_2969;
  reg        [7:0]    _zz_dataOut_payload_0_2970;
  reg        [7:0]    _zz_dataOut_payload_0_2971;
  reg        [7:0]    _zz_dataOut_payload_0_2972;
  reg        [7:0]    _zz_dataOut_payload_0_2973;
  reg        [7:0]    _zz_dataOut_payload_0_2974;
  reg        [7:0]    _zz_dataOut_payload_0_2975;
  reg        [7:0]    _zz_dataOut_payload_0_2976;
  reg        [7:0]    _zz_dataOut_payload_0_2977;
  reg        [7:0]    _zz_dataOut_payload_0_2978;
  reg        [7:0]    _zz_dataOut_payload_0_2979;
  reg        [7:0]    _zz_dataOut_payload_0_2980;
  reg        [7:0]    _zz_dataOut_payload_0_2981;
  reg        [7:0]    _zz_dataOut_payload_0_2982;
  reg        [7:0]    _zz_dataOut_payload_0_2983;
  reg        [7:0]    _zz_dataOut_payload_0_2984;
  reg        [7:0]    _zz_dataOut_payload_0_2985;
  reg        [7:0]    _zz_dataOut_payload_0_2986;
  reg        [7:0]    _zz_dataOut_payload_0_2987;
  reg        [7:0]    _zz_dataOut_payload_0_2988;
  reg        [7:0]    _zz_dataOut_payload_0_2989;
  reg        [7:0]    _zz_dataOut_payload_0_2990;
  reg        [7:0]    _zz_dataOut_payload_0_2991;
  reg        [7:0]    _zz_dataOut_payload_0_2992;
  reg        [7:0]    _zz_dataOut_payload_0_2993;
  reg        [7:0]    _zz_dataOut_payload_0_2994;
  reg        [7:0]    _zz_dataOut_payload_0_2995;
  reg        [7:0]    _zz_dataOut_payload_0_2996;
  reg        [7:0]    _zz_dataOut_payload_0_2997;
  reg        [7:0]    _zz_dataOut_payload_0_2998;
  reg        [7:0]    _zz_dataOut_payload_0_2999;
  reg        [7:0]    _zz_dataOut_payload_0_3000;
  reg        [7:0]    _zz_dataOut_payload_0_3001;
  reg        [7:0]    _zz_dataOut_payload_0_3002;
  reg        [7:0]    _zz_dataOut_payload_0_3003;
  reg        [7:0]    _zz_dataOut_payload_0_3004;
  reg        [7:0]    _zz_dataOut_payload_0_3005;
  reg        [7:0]    _zz_dataOut_payload_0_3006;
  reg        [7:0]    _zz_dataOut_payload_0_3007;
  reg        [7:0]    _zz_dataOut_payload_0_3008;
  reg        [7:0]    _zz_dataOut_payload_0_3009;
  reg        [7:0]    _zz_dataOut_payload_0_3010;
  reg        [7:0]    _zz_dataOut_payload_0_3011;
  reg        [7:0]    _zz_dataOut_payload_0_3012;
  reg        [7:0]    _zz_dataOut_payload_0_3013;
  reg        [7:0]    _zz_dataOut_payload_0_3014;
  reg        [7:0]    _zz_dataOut_payload_0_3015;
  reg        [7:0]    _zz_dataOut_payload_0_3016;
  reg        [7:0]    _zz_dataOut_payload_0_3017;
  reg        [7:0]    _zz_dataOut_payload_0_3018;
  reg        [7:0]    _zz_dataOut_payload_0_3019;
  reg        [7:0]    _zz_dataOut_payload_0_3020;
  reg        [7:0]    _zz_dataOut_payload_0_3021;
  reg        [7:0]    _zz_dataOut_payload_0_3022;
  reg        [7:0]    _zz_dataOut_payload_0_3023;
  reg        [7:0]    _zz_dataOut_payload_0_3024;
  reg        [7:0]    _zz_dataOut_payload_0_3025;
  reg        [7:0]    _zz_dataOut_payload_0_3026;
  reg        [7:0]    _zz_dataOut_payload_0_3027;
  reg        [7:0]    _zz_dataOut_payload_0_3028;
  reg        [7:0]    _zz_dataOut_payload_0_3029;
  reg        [7:0]    _zz_dataOut_payload_0_3030;
  reg        [7:0]    _zz_dataOut_payload_0_3031;
  reg        [7:0]    _zz_dataOut_payload_0_3032;
  reg        [7:0]    _zz_dataOut_payload_0_3033;
  reg        [7:0]    _zz_dataOut_payload_0_3034;
  reg        [7:0]    _zz_dataOut_payload_0_3035;
  reg        [7:0]    _zz_dataOut_payload_0_3036;
  reg        [7:0]    _zz_dataOut_payload_0_3037;
  reg        [7:0]    _zz_dataOut_payload_0_3038;
  reg        [7:0]    _zz_dataOut_payload_0_3039;
  reg        [7:0]    _zz_dataOut_payload_0_3040;
  reg        [7:0]    _zz_dataOut_payload_0_3041;
  reg        [7:0]    _zz_dataOut_payload_0_3042;
  reg        [7:0]    _zz_dataOut_payload_0_3043;
  reg        [7:0]    _zz_dataOut_payload_0_3044;
  reg        [7:0]    _zz_dataOut_payload_0_3045;
  reg        [7:0]    _zz_dataOut_payload_0_3046;
  reg        [7:0]    _zz_dataOut_payload_0_3047;
  reg        [7:0]    _zz_dataOut_payload_0_3048;
  reg        [7:0]    _zz_dataOut_payload_0_3049;
  reg        [7:0]    _zz_dataOut_payload_0_3050;
  reg        [7:0]    _zz_dataOut_payload_0_3051;
  reg        [7:0]    _zz_dataOut_payload_0_3052;
  reg        [7:0]    _zz_dataOut_payload_0_3053;
  reg        [7:0]    _zz_dataOut_payload_0_3054;
  reg        [7:0]    _zz_dataOut_payload_0_3055;
  reg        [7:0]    _zz_dataOut_payload_0_3056;
  reg        [7:0]    _zz_dataOut_payload_0_3057;
  reg        [7:0]    _zz_dataOut_payload_0_3058;
  reg        [7:0]    _zz_dataOut_payload_0_3059;
  reg        [7:0]    _zz_dataOut_payload_0_3060;
  reg        [7:0]    _zz_dataOut_payload_0_3061;
  reg        [7:0]    _zz_dataOut_payload_0_3062;
  reg        [7:0]    _zz_dataOut_payload_0_3063;
  reg        [7:0]    _zz_dataOut_payload_0_3064;
  reg        [7:0]    _zz_dataOut_payload_0_3065;
  reg        [7:0]    _zz_dataOut_payload_0_3066;
  reg        [7:0]    _zz_dataOut_payload_0_3067;
  reg        [7:0]    _zz_dataOut_payload_0_3068;
  reg        [7:0]    _zz_dataOut_payload_0_3069;
  reg        [7:0]    _zz_dataOut_payload_0_3070;
  reg        [7:0]    _zz_dataOut_payload_0_3071;
  wire                _zz_dataOut_payload_0_3072;
  wire       [7:0]    _zz_dataOut_payload_0_3073;
  wire       [7:0]    _zz_dataOut_payload_0_3074;
  wire                _zz_dataOut_payload_0_3075;
  wire       [7:0]    _zz_dataOut_payload_0_3076;
  wire       [7:0]    _zz_dataOut_payload_0_3077;
  wire                _zz_dataOut_payload_0_3078;
  wire       [7:0]    _zz_dataOut_payload_0_3079;
  wire       [7:0]    _zz_dataOut_payload_0_3080;
  wire                _zz_dataOut_payload_0_3081;
  wire       [7:0]    _zz_dataOut_payload_0_3082;
  wire       [7:0]    _zz_dataOut_payload_0_3083;
  wire                _zz_dataOut_payload_0_3084;
  wire       [7:0]    _zz_dataOut_payload_0_3085;
  wire       [7:0]    _zz_dataOut_payload_0_3086;
  wire                _zz_dataOut_payload_0_3087;
  wire       [7:0]    _zz_dataOut_payload_0_3088;
  wire       [7:0]    _zz_dataOut_payload_0_3089;
  wire                _zz_dataOut_payload_0_3090;
  wire       [7:0]    _zz_dataOut_payload_0_3091;
  wire       [7:0]    _zz_dataOut_payload_0_3092;
  wire                _zz_dataOut_payload_0_3093;
  wire       [7:0]    _zz_dataOut_payload_0_3094;
  wire       [7:0]    _zz_dataOut_payload_0_3095;
  wire                _zz_dataOut_payload_0_3096;
  wire       [7:0]    _zz_dataOut_payload_0_3097;
  wire       [7:0]    _zz_dataOut_payload_0_3098;
  wire                _zz_dataOut_payload_0_3099;
  wire       [7:0]    _zz_dataOut_payload_0_3100;
  wire       [7:0]    _zz_dataOut_payload_0_3101;
  wire                _zz_dataOut_payload_0_3102;
  wire       [7:0]    _zz_dataOut_payload_0_3103;
  wire       [7:0]    _zz_dataOut_payload_0_3104;
  wire                _zz_dataOut_payload_0_3105;
  wire       [7:0]    _zz_dataOut_payload_0_3106;
  wire       [7:0]    _zz_dataOut_payload_0_3107;
  wire                _zz_dataOut_payload_0_3108;
  wire       [7:0]    _zz_dataOut_payload_0_3109;
  wire       [7:0]    _zz_dataOut_payload_0_3110;
  wire                _zz_dataOut_payload_0_3111;
  wire       [7:0]    _zz_dataOut_payload_0_3112;
  wire       [7:0]    _zz_dataOut_payload_0_3113;
  wire                _zz_dataOut_payload_0_3114;
  wire                _zz_dataOut_payload_0_3115;
  reg        [7:0]    _zz_dataOut_payload_0_3116;
  reg        [7:0]    _zz_dataOut_payload_0_3117;
  reg        [7:0]    _zz_dataOut_payload_0_3118;
  reg        [7:0]    _zz_dataOut_payload_0_3119;
  wire                _zz_dataOut_payload_0_3120;
  wire       [7:0]    _zz_dataOut_payload_0_3121;
  wire       [7:0]    _zz_dataOut_payload_0_3122;
  wire                _zz_dataOut_payload_0_3123;
  wire       [7:0]    _zz_dataOut_payload_0_3124;
  wire       [7:0]    _zz_dataOut_payload_0_3125;
  wire                _zz_dataOut_payload_0_3126;
  wire                _zz_dataOut_payload_0_3127;
  reg        [7:0]    _zz_dataOut_payload_0_3128;
  reg        [7:0]    _zz_dataOut_payload_0_3129;
  reg        [7:0]    _zz_dataOut_payload_0_3130;
  reg        [7:0]    _zz_dataOut_payload_0_3131;
  reg        [7:0]    _zz_dataOut_payload_0_3132;
  reg        [7:0]    _zz_dataOut_payload_0_3133;
  reg        [7:0]    _zz_dataOut_payload_0_3134;
  reg        [7:0]    _zz_dataOut_payload_0_3135;
  reg        [7:0]    _zz_dataOut_payload_0_3136;
  reg        [7:0]    _zz_dataOut_payload_0_3137;
  reg        [7:0]    _zz_dataOut_payload_0_3138;
  reg        [7:0]    _zz_dataOut_payload_0_3139;
  wire                _zz_dataOut_payload_0_3140;
  wire       [7:0]    _zz_dataOut_payload_0_3141;
  wire       [7:0]    _zz_dataOut_payload_0_3142;
  wire                _zz_dataOut_payload_0_3143;
  wire       [7:0]    _zz_dataOut_payload_0_3144;
  wire       [7:0]    _zz_dataOut_payload_0_3145;
  wire                _zz_dataOut_payload_0_3146;
  wire       [7:0]    _zz_dataOut_payload_0_3147;
  wire       [7:0]    _zz_dataOut_payload_0_3148;
  wire                _zz_dataOut_payload_0_3149;
  wire       [7:0]    _zz_dataOut_payload_0_3150;
  wire       [7:0]    _zz_dataOut_payload_0_3151;
  wire                _zz_dataOut_payload_0_3152;
  wire       [7:0]    _zz_dataOut_payload_0_3153;
  wire       [7:0]    _zz_dataOut_payload_0_3154;
  wire                _zz_dataOut_payload_0_3155;
  wire       [7:0]    _zz_dataOut_payload_0_3156;
  wire       [7:0]    _zz_dataOut_payload_0_3157;
  wire                _zz_dataOut_payload_0_3158;
  wire                _zz_dataOut_payload_0_3159;
  reg        [7:0]    _zz_dataOut_payload_0_3160;
  reg        [7:0]    _zz_dataOut_payload_0_3161;
  reg        [7:0]    _zz_dataOut_payload_0_3162;
  reg        [7:0]    _zz_dataOut_payload_0_3163;
  wire                _zz_dataOut_payload_0_3164;
  wire       [7:0]    _zz_dataOut_payload_0_3165;
  wire       [7:0]    _zz_dataOut_payload_0_3166;
  wire                _zz_dataOut_payload_0_3167;
  wire       [7:0]    _zz_dataOut_payload_0_3168;
  wire       [7:0]    _zz_dataOut_payload_0_3169;
  wire                _zz_dataOut_payload_0_3170;
  wire                _zz_dataOut_payload_0_3171;
  reg        [7:0]    _zz_dataOut_payload_0_3172;
  reg        [7:0]    _zz_dataOut_payload_0_3173;
  reg        [7:0]    _zz_dataOut_payload_0_3174;
  reg        [7:0]    _zz_dataOut_payload_0_3175;
  reg        [7:0]    _zz_dataOut_payload_0_3176;
  reg        [7:0]    _zz_dataOut_payload_0_3177;
  reg        [7:0]    _zz_dataOut_payload_0_3178;
  reg        [7:0]    _zz_dataOut_payload_0_3179;
  reg        [7:0]    _zz_dataOut_payload_0_3180;
  reg        [7:0]    _zz_dataOut_payload_0_3181;
  reg        [7:0]    _zz_dataOut_payload_0_3182;
  reg        [7:0]    _zz_dataOut_payload_0_3183;
  reg        [7:0]    _zz_dataOut_payload_0_3184;
  reg        [7:0]    _zz_dataOut_payload_0_3185;
  reg        [7:0]    _zz_dataOut_payload_0_3186;
  reg        [7:0]    _zz_dataOut_payload_0_3187;
  reg        [7:0]    _zz_dataOut_payload_0_3188;
  reg        [7:0]    _zz_dataOut_payload_0_3189;
  reg        [7:0]    _zz_dataOut_payload_0_3190;
  reg        [7:0]    _zz_dataOut_payload_0_3191;
  reg        [7:0]    _zz_dataOut_payload_0_3192;
  reg        [7:0]    _zz_dataOut_payload_0_3193;
  reg        [7:0]    _zz_dataOut_payload_0_3194;
  reg        [7:0]    _zz_dataOut_payload_0_3195;
  reg        [7:0]    _zz_dataOut_payload_0_3196;
  reg        [7:0]    _zz_dataOut_payload_0_3197;
  reg        [7:0]    _zz_dataOut_payload_0_3198;
  reg        [7:0]    _zz_dataOut_payload_0_3199;
  wire                _zz_dataOut_payload_0_3200;
  wire       [7:0]    _zz_dataOut_payload_0_3201;
  wire       [7:0]    _zz_dataOut_payload_0_3202;
  wire                _zz_dataOut_payload_0_3203;
  wire       [7:0]    _zz_dataOut_payload_0_3204;
  wire       [7:0]    _zz_dataOut_payload_0_3205;
  wire                _zz_dataOut_payload_0_3206;
  wire       [7:0]    _zz_dataOut_payload_0_3207;
  wire       [7:0]    _zz_dataOut_payload_0_3208;
  wire                _zz_dataOut_payload_0_3209;
  wire       [7:0]    _zz_dataOut_payload_0_3210;
  wire       [7:0]    _zz_dataOut_payload_0_3211;
  wire                _zz_dataOut_payload_0_3212;
  wire       [7:0]    _zz_dataOut_payload_0_3213;
  wire       [7:0]    _zz_dataOut_payload_0_3214;
  wire                _zz_dataOut_payload_0_3215;
  wire       [7:0]    _zz_dataOut_payload_0_3216;
  wire       [7:0]    _zz_dataOut_payload_0_3217;
  wire                _zz_dataOut_payload_0_3218;
  wire       [7:0]    _zz_dataOut_payload_0_3219;
  wire       [7:0]    _zz_dataOut_payload_0_3220;
  wire                _zz_dataOut_payload_0_3221;
  wire       [7:0]    _zz_dataOut_payload_0_3222;
  wire       [7:0]    _zz_dataOut_payload_0_3223;
  wire                _zz_dataOut_payload_0_3224;
  wire       [7:0]    _zz_dataOut_payload_0_3225;
  wire       [7:0]    _zz_dataOut_payload_0_3226;
  wire                _zz_dataOut_payload_0_3227;
  wire       [7:0]    _zz_dataOut_payload_0_3228;
  wire       [7:0]    _zz_dataOut_payload_0_3229;
  wire                _zz_dataOut_payload_0_3230;
  wire       [7:0]    _zz_dataOut_payload_0_3231;
  wire       [7:0]    _zz_dataOut_payload_0_3232;
  wire                _zz_dataOut_payload_0_3233;
  wire       [7:0]    _zz_dataOut_payload_0_3234;
  wire       [7:0]    _zz_dataOut_payload_0_3235;
  wire                _zz_dataOut_payload_0_3236;
  wire       [7:0]    _zz_dataOut_payload_0_3237;
  wire       [7:0]    _zz_dataOut_payload_0_3238;
  wire                _zz_dataOut_payload_0_3239;
  wire       [7:0]    _zz_dataOut_payload_0_3240;
  wire       [7:0]    _zz_dataOut_payload_0_3241;
  wire                _zz_dataOut_payload_0_3242;
  wire                _zz_dataOut_payload_0_3243;
  reg        [7:0]    _zz_dataOut_payload_0_3244;
  reg        [7:0]    _zz_dataOut_payload_0_3245;
  reg        [7:0]    _zz_dataOut_payload_0_3246;
  reg        [7:0]    _zz_dataOut_payload_0_3247;
  wire                _zz_dataOut_payload_0_3248;
  wire       [7:0]    _zz_dataOut_payload_0_3249;
  wire       [7:0]    _zz_dataOut_payload_0_3250;
  wire                _zz_dataOut_payload_0_3251;
  wire       [7:0]    _zz_dataOut_payload_0_3252;
  wire       [7:0]    _zz_dataOut_payload_0_3253;
  wire                _zz_dataOut_payload_0_3254;
  wire                _zz_dataOut_payload_0_3255;
  reg        [7:0]    _zz_dataOut_payload_0_3256;
  reg        [7:0]    _zz_dataOut_payload_0_3257;
  reg        [7:0]    _zz_dataOut_payload_0_3258;
  reg        [7:0]    _zz_dataOut_payload_0_3259;
  reg        [7:0]    _zz_dataOut_payload_0_3260;
  reg        [7:0]    _zz_dataOut_payload_0_3261;
  reg        [7:0]    _zz_dataOut_payload_0_3262;
  reg        [7:0]    _zz_dataOut_payload_0_3263;
  reg        [7:0]    _zz_dataOut_payload_0_3264;
  reg        [7:0]    _zz_dataOut_payload_0_3265;
  reg        [7:0]    _zz_dataOut_payload_0_3266;
  reg        [7:0]    _zz_dataOut_payload_0_3267;
  wire                _zz_dataOut_payload_0_3268;
  wire       [7:0]    _zz_dataOut_payload_0_3269;
  wire       [7:0]    _zz_dataOut_payload_0_3270;
  wire                _zz_dataOut_payload_0_3271;
  wire       [7:0]    _zz_dataOut_payload_0_3272;
  wire       [7:0]    _zz_dataOut_payload_0_3273;
  wire                _zz_dataOut_payload_0_3274;
  wire       [7:0]    _zz_dataOut_payload_0_3275;
  wire       [7:0]    _zz_dataOut_payload_0_3276;
  wire                _zz_dataOut_payload_0_3277;
  wire       [7:0]    _zz_dataOut_payload_0_3278;
  wire       [7:0]    _zz_dataOut_payload_0_3279;
  wire                _zz_dataOut_payload_0_3280;
  wire       [7:0]    _zz_dataOut_payload_0_3281;
  wire       [7:0]    _zz_dataOut_payload_0_3282;
  wire                _zz_dataOut_payload_0_3283;
  wire       [7:0]    _zz_dataOut_payload_0_3284;
  wire       [7:0]    _zz_dataOut_payload_0_3285;
  wire                _zz_dataOut_payload_0_3286;
  wire                _zz_dataOut_payload_0_3287;
  reg        [7:0]    _zz_dataOut_payload_0_3288;
  reg        [7:0]    _zz_dataOut_payload_0_3289;
  reg        [7:0]    _zz_dataOut_payload_0_3290;
  reg        [7:0]    _zz_dataOut_payload_0_3291;
  wire                _zz_dataOut_payload_0_3292;
  wire       [7:0]    _zz_dataOut_payload_0_3293;
  wire       [7:0]    _zz_dataOut_payload_0_3294;
  wire                _zz_dataOut_payload_0_3295;
  wire       [7:0]    _zz_dataOut_payload_0_3296;
  wire       [7:0]    _zz_dataOut_payload_0_3297;
  wire                _zz_dataOut_payload_0_3298;
  wire                _zz_dataOut_payload_0_3299;
  reg        [7:0]    _zz_dataOut_payload_0_3300;
  reg        [7:0]    _zz_dataOut_payload_0_3301;
  reg        [7:0]    _zz_dataOut_payload_0_3302;
  reg        [7:0]    _zz_dataOut_payload_0_3303;
  reg        [7:0]    _zz_dataOut_payload_0_3304;
  reg        [7:0]    _zz_dataOut_payload_0_3305;
  reg        [7:0]    _zz_dataOut_payload_0_3306;
  reg        [7:0]    _zz_dataOut_payload_0_3307;
  reg        [7:0]    _zz_dataOut_payload_0_3308;
  reg        [7:0]    _zz_dataOut_payload_0_3309;
  reg        [7:0]    _zz_dataOut_payload_0_3310;
  reg        [7:0]    _zz_dataOut_payload_0_3311;
  reg        [7:0]    _zz_dataOut_payload_0_3312;
  reg        [7:0]    _zz_dataOut_payload_0_3313;
  reg        [7:0]    _zz_dataOut_payload_0_3314;
  reg        [7:0]    _zz_dataOut_payload_0_3315;
  reg        [7:0]    _zz_dataOut_payload_0_3316;
  reg        [7:0]    _zz_dataOut_payload_0_3317;
  reg        [7:0]    _zz_dataOut_payload_0_3318;
  reg        [7:0]    _zz_dataOut_payload_0_3319;
  reg        [7:0]    _zz_dataOut_payload_0_3320;
  reg        [7:0]    _zz_dataOut_payload_0_3321;
  reg        [7:0]    _zz_dataOut_payload_0_3322;
  reg        [7:0]    _zz_dataOut_payload_0_3323;
  reg        [7:0]    _zz_dataOut_payload_0_3324;
  reg        [7:0]    _zz_dataOut_payload_0_3325;
  reg        [7:0]    _zz_dataOut_payload_0_3326;
  reg        [7:0]    _zz_dataOut_payload_0_3327;
  wire                _zz_dataOut_payload_0_3328;
  wire       [7:0]    _zz_dataOut_payload_0_3329;
  wire       [7:0]    _zz_dataOut_payload_0_3330;
  wire                _zz_dataOut_payload_0_3331;
  wire       [7:0]    _zz_dataOut_payload_0_3332;
  wire       [7:0]    _zz_dataOut_payload_0_3333;
  wire                _zz_dataOut_payload_0_3334;
  wire       [7:0]    _zz_dataOut_payload_0_3335;
  wire       [7:0]    _zz_dataOut_payload_0_3336;
  wire                _zz_dataOut_payload_0_3337;
  wire       [7:0]    _zz_dataOut_payload_0_3338;
  wire       [7:0]    _zz_dataOut_payload_0_3339;
  wire                _zz_dataOut_payload_0_3340;
  wire       [7:0]    _zz_dataOut_payload_0_3341;
  wire       [7:0]    _zz_dataOut_payload_0_3342;
  wire                _zz_dataOut_payload_0_3343;
  wire       [7:0]    _zz_dataOut_payload_0_3344;
  wire       [7:0]    _zz_dataOut_payload_0_3345;
  wire                _zz_dataOut_payload_0_3346;
  wire       [7:0]    _zz_dataOut_payload_0_3347;
  wire       [7:0]    _zz_dataOut_payload_0_3348;
  wire                _zz_dataOut_payload_0_3349;
  wire       [7:0]    _zz_dataOut_payload_0_3350;
  wire       [7:0]    _zz_dataOut_payload_0_3351;
  wire                _zz_dataOut_payload_0_3352;
  wire       [7:0]    _zz_dataOut_payload_0_3353;
  wire       [7:0]    _zz_dataOut_payload_0_3354;
  wire                _zz_dataOut_payload_0_3355;
  wire       [7:0]    _zz_dataOut_payload_0_3356;
  wire       [7:0]    _zz_dataOut_payload_0_3357;
  wire                _zz_dataOut_payload_0_3358;
  wire       [7:0]    _zz_dataOut_payload_0_3359;
  wire       [7:0]    _zz_dataOut_payload_0_3360;
  wire                _zz_dataOut_payload_0_3361;
  wire       [7:0]    _zz_dataOut_payload_0_3362;
  wire       [7:0]    _zz_dataOut_payload_0_3363;
  wire                _zz_dataOut_payload_0_3364;
  wire       [7:0]    _zz_dataOut_payload_0_3365;
  wire       [7:0]    _zz_dataOut_payload_0_3366;
  wire                _zz_dataOut_payload_0_3367;
  wire       [7:0]    _zz_dataOut_payload_0_3368;
  wire       [7:0]    _zz_dataOut_payload_0_3369;
  wire                _zz_dataOut_payload_0_3370;
  wire                _zz_dataOut_payload_0_3371;
  reg        [7:0]    _zz_dataOut_payload_0_3372;
  reg        [7:0]    _zz_dataOut_payload_0_3373;
  reg        [7:0]    _zz_dataOut_payload_0_3374;
  reg        [7:0]    _zz_dataOut_payload_0_3375;
  wire                _zz_dataOut_payload_0_3376;
  wire       [7:0]    _zz_dataOut_payload_0_3377;
  wire       [7:0]    _zz_dataOut_payload_0_3378;
  wire                _zz_dataOut_payload_0_3379;
  wire       [7:0]    _zz_dataOut_payload_0_3380;
  wire       [7:0]    _zz_dataOut_payload_0_3381;
  wire                _zz_dataOut_payload_0_3382;
  wire                _zz_dataOut_payload_0_3383;
  reg        [7:0]    _zz_dataOut_payload_0_3384;
  reg        [7:0]    _zz_dataOut_payload_0_3385;
  reg        [7:0]    _zz_dataOut_payload_0_3386;
  reg        [7:0]    _zz_dataOut_payload_0_3387;
  reg        [7:0]    _zz_dataOut_payload_0_3388;
  reg        [7:0]    _zz_dataOut_payload_0_3389;
  reg        [7:0]    _zz_dataOut_payload_0_3390;
  reg        [7:0]    _zz_dataOut_payload_0_3391;
  reg        [7:0]    _zz_dataOut_payload_0_3392;
  reg        [7:0]    _zz_dataOut_payload_0_3393;
  reg        [7:0]    _zz_dataOut_payload_0_3394;
  reg        [7:0]    _zz_dataOut_payload_0_3395;
  wire                _zz_dataOut_payload_0_3396;
  wire       [7:0]    _zz_dataOut_payload_0_3397;
  wire       [7:0]    _zz_dataOut_payload_0_3398;
  wire                _zz_dataOut_payload_0_3399;
  wire       [7:0]    _zz_dataOut_payload_0_3400;
  wire       [7:0]    _zz_dataOut_payload_0_3401;
  wire                _zz_dataOut_payload_0_3402;
  wire       [7:0]    _zz_dataOut_payload_0_3403;
  wire       [7:0]    _zz_dataOut_payload_0_3404;
  wire                _zz_dataOut_payload_0_3405;
  wire       [7:0]    _zz_dataOut_payload_0_3406;
  wire       [7:0]    _zz_dataOut_payload_0_3407;
  wire                _zz_dataOut_payload_0_3408;
  wire       [7:0]    _zz_dataOut_payload_0_3409;
  wire       [7:0]    _zz_dataOut_payload_0_3410;
  wire                _zz_dataOut_payload_0_3411;
  wire       [7:0]    _zz_dataOut_payload_0_3412;
  wire       [7:0]    _zz_dataOut_payload_0_3413;
  wire                _zz_dataOut_payload_0_3414;
  wire                _zz_dataOut_payload_0_3415;
  reg        [7:0]    _zz_dataOut_payload_0_3416;
  reg        [7:0]    _zz_dataOut_payload_0_3417;
  reg        [7:0]    _zz_dataOut_payload_0_3418;
  reg        [7:0]    _zz_dataOut_payload_0_3419;
  wire                _zz_dataOut_payload_0_3420;
  wire       [7:0]    _zz_dataOut_payload_0_3421;
  wire       [7:0]    _zz_dataOut_payload_0_3422;
  wire                _zz_dataOut_payload_0_3423;
  wire       [7:0]    _zz_dataOut_payload_0_3424;
  wire       [7:0]    _zz_dataOut_payload_0_3425;
  wire                _zz_dataOut_payload_0_3426;
  wire                _zz_dataOut_payload_0_3427;
  reg        [7:0]    _zz_dataOut_payload_0_3428;
  reg        [7:0]    _zz_dataOut_payload_0_3429;
  reg        [7:0]    _zz_dataOut_payload_0_3430;
  reg        [7:0]    _zz_dataOut_payload_0_3431;
  reg        [7:0]    _zz_dataOut_payload_0_3432;
  reg        [7:0]    _zz_dataOut_payload_0_3433;
  reg        [7:0]    _zz_dataOut_payload_0_3434;
  reg        [7:0]    _zz_dataOut_payload_0_3435;
  reg        [7:0]    _zz_dataOut_payload_0_3436;
  reg        [7:0]    _zz_dataOut_payload_0_3437;
  reg        [7:0]    _zz_dataOut_payload_0_3438;
  reg        [7:0]    _zz_dataOut_payload_0_3439;
  reg        [7:0]    _zz_dataOut_payload_0_3440;
  reg        [7:0]    _zz_dataOut_payload_0_3441;
  reg        [7:0]    _zz_dataOut_payload_0_3442;
  reg        [7:0]    _zz_dataOut_payload_0_3443;
  reg        [7:0]    _zz_dataOut_payload_0_3444;
  reg        [7:0]    _zz_dataOut_payload_0_3445;
  reg        [7:0]    _zz_dataOut_payload_0_3446;
  reg        [7:0]    _zz_dataOut_payload_0_3447;
  reg        [7:0]    _zz_dataOut_payload_0_3448;
  reg        [7:0]    _zz_dataOut_payload_0_3449;
  reg        [7:0]    _zz_dataOut_payload_0_3450;
  reg        [7:0]    _zz_dataOut_payload_0_3451;
  reg        [7:0]    _zz_dataOut_payload_0_3452;
  reg        [7:0]    _zz_dataOut_payload_0_3453;
  reg        [7:0]    _zz_dataOut_payload_0_3454;
  reg        [7:0]    _zz_dataOut_payload_0_3455;
  wire                _zz_dataOut_payload_0_3456;
  wire       [7:0]    _zz_dataOut_payload_0_3457;
  wire       [7:0]    _zz_dataOut_payload_0_3458;
  wire                _zz_dataOut_payload_0_3459;
  wire       [7:0]    _zz_dataOut_payload_0_3460;
  wire       [7:0]    _zz_dataOut_payload_0_3461;
  wire                _zz_dataOut_payload_0_3462;
  wire       [7:0]    _zz_dataOut_payload_0_3463;
  wire       [7:0]    _zz_dataOut_payload_0_3464;
  wire                _zz_dataOut_payload_0_3465;
  wire       [7:0]    _zz_dataOut_payload_0_3466;
  wire       [7:0]    _zz_dataOut_payload_0_3467;
  wire                _zz_dataOut_payload_0_3468;
  wire       [7:0]    _zz_dataOut_payload_0_3469;
  wire       [7:0]    _zz_dataOut_payload_0_3470;
  wire                _zz_dataOut_payload_0_3471;
  wire       [7:0]    _zz_dataOut_payload_0_3472;
  wire       [7:0]    _zz_dataOut_payload_0_3473;
  wire                _zz_dataOut_payload_0_3474;
  wire       [7:0]    _zz_dataOut_payload_0_3475;
  wire       [7:0]    _zz_dataOut_payload_0_3476;
  wire                _zz_dataOut_payload_0_3477;
  wire       [7:0]    _zz_dataOut_payload_0_3478;
  wire       [7:0]    _zz_dataOut_payload_0_3479;
  wire                _zz_dataOut_payload_0_3480;
  wire       [7:0]    _zz_dataOut_payload_0_3481;
  wire       [7:0]    _zz_dataOut_payload_0_3482;
  wire                _zz_dataOut_payload_0_3483;
  wire       [7:0]    _zz_dataOut_payload_0_3484;
  wire       [7:0]    _zz_dataOut_payload_0_3485;
  wire                _zz_dataOut_payload_0_3486;
  wire       [7:0]    _zz_dataOut_payload_0_3487;
  wire       [7:0]    _zz_dataOut_payload_0_3488;
  wire                _zz_dataOut_payload_0_3489;
  wire       [7:0]    _zz_dataOut_payload_0_3490;
  wire       [7:0]    _zz_dataOut_payload_0_3491;
  wire                _zz_dataOut_payload_0_3492;
  wire       [7:0]    _zz_dataOut_payload_0_3493;
  wire       [7:0]    _zz_dataOut_payload_0_3494;
  wire                _zz_dataOut_payload_0_3495;
  wire       [7:0]    _zz_dataOut_payload_0_3496;
  wire       [7:0]    _zz_dataOut_payload_0_3497;
  wire                _zz_dataOut_payload_0_3498;
  wire                _zz_dataOut_payload_0_3499;
  reg        [7:0]    _zz_dataOut_payload_0_3500;
  reg        [7:0]    _zz_dataOut_payload_0_3501;
  reg        [7:0]    _zz_dataOut_payload_0_3502;
  reg        [7:0]    _zz_dataOut_payload_0_3503;
  wire                _zz_dataOut_payload_0_3504;
  wire       [7:0]    _zz_dataOut_payload_0_3505;
  wire       [7:0]    _zz_dataOut_payload_0_3506;
  wire                _zz_dataOut_payload_0_3507;
  wire       [7:0]    _zz_dataOut_payload_0_3508;
  wire       [7:0]    _zz_dataOut_payload_0_3509;
  wire                _zz_dataOut_payload_0_3510;
  wire                _zz_dataOut_payload_0_3511;
  reg        [7:0]    _zz_dataOut_payload_0_3512;
  reg        [7:0]    _zz_dataOut_payload_0_3513;
  reg        [7:0]    _zz_dataOut_payload_0_3514;
  reg        [7:0]    _zz_dataOut_payload_0_3515;
  reg        [7:0]    _zz_dataOut_payload_0_3516;
  reg        [7:0]    _zz_dataOut_payload_0_3517;
  reg        [7:0]    _zz_dataOut_payload_0_3518;
  reg        [7:0]    _zz_dataOut_payload_0_3519;
  reg        [7:0]    _zz_dataOut_payload_0_3520;
  reg        [7:0]    _zz_dataOut_payload_0_3521;
  reg        [7:0]    _zz_dataOut_payload_0_3522;
  reg        [7:0]    _zz_dataOut_payload_0_3523;
  wire                _zz_dataOut_payload_0_3524;
  wire       [7:0]    _zz_dataOut_payload_0_3525;
  wire       [7:0]    _zz_dataOut_payload_0_3526;
  wire                _zz_dataOut_payload_0_3527;
  wire       [7:0]    _zz_dataOut_payload_0_3528;
  wire       [7:0]    _zz_dataOut_payload_0_3529;
  wire                _zz_dataOut_payload_0_3530;
  wire       [7:0]    _zz_dataOut_payload_0_3531;
  wire       [7:0]    _zz_dataOut_payload_0_3532;
  wire                _zz_dataOut_payload_0_3533;
  wire       [7:0]    _zz_dataOut_payload_0_3534;
  wire       [7:0]    _zz_dataOut_payload_0_3535;
  wire                _zz_dataOut_payload_0_3536;
  wire       [7:0]    _zz_dataOut_payload_0_3537;
  wire       [7:0]    _zz_dataOut_payload_0_3538;
  wire                _zz_dataOut_payload_0_3539;
  wire       [7:0]    _zz_dataOut_payload_0_3540;
  wire       [7:0]    _zz_dataOut_payload_0_3541;
  wire                _zz_dataOut_payload_0_3542;
  wire                _zz_dataOut_payload_0_3543;
  reg        [7:0]    _zz_dataOut_payload_0_3544;
  reg        [7:0]    _zz_dataOut_payload_0_3545;
  reg        [7:0]    _zz_dataOut_payload_0_3546;
  reg        [7:0]    _zz_dataOut_payload_0_3547;
  wire                _zz_dataOut_payload_0_3548;
  wire       [7:0]    _zz_dataOut_payload_0_3549;
  wire       [7:0]    _zz_dataOut_payload_0_3550;
  wire                _zz_dataOut_payload_0_3551;
  wire       [7:0]    _zz_dataOut_payload_0_3552;
  wire       [7:0]    _zz_dataOut_payload_0_3553;
  wire                _zz_dataOut_payload_0_3554;
  wire                _zz_dataOut_payload_0_3555;
  reg        [7:0]    _zz_dataOut_payload_0_3556;
  reg        [7:0]    _zz_dataOut_payload_0_3557;
  reg        [7:0]    _zz_dataOut_payload_0_3558;
  reg        [7:0]    _zz_dataOut_payload_0_3559;
  reg        [7:0]    _zz_dataOut_payload_0_3560;
  reg        [7:0]    _zz_dataOut_payload_0_3561;
  reg        [7:0]    _zz_dataOut_payload_0_3562;
  reg        [7:0]    _zz_dataOut_payload_0_3563;
  reg        [7:0]    _zz_dataOut_payload_0_3564;
  reg        [7:0]    _zz_dataOut_payload_0_3565;
  reg        [7:0]    _zz_dataOut_payload_0_3566;
  reg        [7:0]    _zz_dataOut_payload_0_3567;
  reg        [7:0]    _zz_dataOut_payload_0_3568;
  reg        [7:0]    _zz_dataOut_payload_0_3569;
  reg        [7:0]    _zz_dataOut_payload_0_3570;
  reg        [7:0]    _zz_dataOut_payload_0_3571;
  reg        [7:0]    _zz_dataOut_payload_0_3572;
  reg        [7:0]    _zz_dataOut_payload_0_3573;
  reg        [7:0]    _zz_dataOut_payload_0_3574;
  reg        [7:0]    _zz_dataOut_payload_0_3575;
  reg        [7:0]    _zz_dataOut_payload_0_3576;
  reg        [7:0]    _zz_dataOut_payload_0_3577;
  reg        [7:0]    _zz_dataOut_payload_0_3578;
  reg        [7:0]    _zz_dataOut_payload_0_3579;
  reg        [7:0]    _zz_dataOut_payload_0_3580;
  reg        [7:0]    _zz_dataOut_payload_0_3581;
  reg        [7:0]    _zz_dataOut_payload_0_3582;
  reg        [7:0]    _zz_dataOut_payload_0_3583;
  wire                _zz_dataOut_payload_0_3584;
  wire       [7:0]    _zz_dataOut_payload_0_3585;
  wire       [7:0]    _zz_dataOut_payload_0_3586;
  wire                _zz_dataOut_payload_0_3587;
  wire       [7:0]    _zz_dataOut_payload_0_3588;
  wire       [7:0]    _zz_dataOut_payload_0_3589;
  wire                _zz_dataOut_payload_0_3590;
  wire       [7:0]    _zz_dataOut_payload_0_3591;
  wire       [7:0]    _zz_dataOut_payload_0_3592;
  wire                _zz_dataOut_payload_0_3593;
  wire       [7:0]    _zz_dataOut_payload_0_3594;
  wire       [7:0]    _zz_dataOut_payload_0_3595;
  wire                _zz_dataOut_payload_0_3596;
  wire       [7:0]    _zz_dataOut_payload_0_3597;
  wire       [7:0]    _zz_dataOut_payload_0_3598;
  wire                _zz_dataOut_payload_0_3599;
  wire       [7:0]    _zz_dataOut_payload_0_3600;
  wire       [7:0]    _zz_dataOut_payload_0_3601;
  wire                _zz_dataOut_payload_0_3602;
  wire       [7:0]    _zz_dataOut_payload_0_3603;
  wire       [7:0]    _zz_dataOut_payload_0_3604;
  wire                _zz_dataOut_payload_0_3605;
  wire       [7:0]    _zz_dataOut_payload_0_3606;
  wire       [7:0]    _zz_dataOut_payload_0_3607;
  wire                _zz_dataOut_payload_0_3608;
  wire       [7:0]    _zz_dataOut_payload_0_3609;
  wire       [7:0]    _zz_dataOut_payload_0_3610;
  wire                _zz_dataOut_payload_0_3611;
  wire       [7:0]    _zz_dataOut_payload_0_3612;
  wire       [7:0]    _zz_dataOut_payload_0_3613;
  wire                _zz_dataOut_payload_0_3614;
  wire       [7:0]    _zz_dataOut_payload_0_3615;
  wire       [7:0]    _zz_dataOut_payload_0_3616;
  wire                _zz_dataOut_payload_0_3617;
  wire       [7:0]    _zz_dataOut_payload_0_3618;
  wire       [7:0]    _zz_dataOut_payload_0_3619;
  wire                _zz_dataOut_payload_0_3620;
  wire       [7:0]    _zz_dataOut_payload_0_3621;
  wire       [7:0]    _zz_dataOut_payload_0_3622;
  wire                _zz_dataOut_payload_0_3623;
  wire       [7:0]    _zz_dataOut_payload_0_3624;
  wire       [7:0]    _zz_dataOut_payload_0_3625;
  wire                _zz_dataOut_payload_0_3626;
  wire                _zz_dataOut_payload_0_3627;
  reg        [7:0]    _zz_dataOut_payload_0_3628;
  reg        [7:0]    _zz_dataOut_payload_0_3629;
  reg        [7:0]    _zz_dataOut_payload_0_3630;
  reg        [7:0]    _zz_dataOut_payload_0_3631;
  wire                _zz_dataOut_payload_0_3632;
  wire       [7:0]    _zz_dataOut_payload_0_3633;
  wire       [7:0]    _zz_dataOut_payload_0_3634;
  wire                _zz_dataOut_payload_0_3635;
  wire       [7:0]    _zz_dataOut_payload_0_3636;
  wire       [7:0]    _zz_dataOut_payload_0_3637;
  wire                _zz_dataOut_payload_0_3638;
  wire                _zz_dataOut_payload_0_3639;
  reg        [7:0]    _zz_dataOut_payload_0_3640;
  reg        [7:0]    _zz_dataOut_payload_0_3641;
  reg        [7:0]    _zz_dataOut_payload_0_3642;
  reg        [7:0]    _zz_dataOut_payload_0_3643;
  reg        [7:0]    _zz_dataOut_payload_0_3644;
  reg        [7:0]    _zz_dataOut_payload_0_3645;
  reg        [7:0]    _zz_dataOut_payload_0_3646;
  reg        [7:0]    _zz_dataOut_payload_0_3647;
  reg        [7:0]    _zz_dataOut_payload_0_3648;
  reg        [7:0]    _zz_dataOut_payload_0_3649;
  reg        [7:0]    _zz_dataOut_payload_0_3650;
  reg        [7:0]    _zz_dataOut_payload_0_3651;
  wire                _zz_dataOut_payload_0_3652;
  wire       [7:0]    _zz_dataOut_payload_0_3653;
  wire       [7:0]    _zz_dataOut_payload_0_3654;
  wire                _zz_dataOut_payload_0_3655;
  wire       [7:0]    _zz_dataOut_payload_0_3656;
  wire       [7:0]    _zz_dataOut_payload_0_3657;
  wire                _zz_dataOut_payload_0_3658;
  wire       [7:0]    _zz_dataOut_payload_0_3659;
  wire       [7:0]    _zz_dataOut_payload_0_3660;
  wire                _zz_dataOut_payload_0_3661;
  wire       [7:0]    _zz_dataOut_payload_0_3662;
  wire       [7:0]    _zz_dataOut_payload_0_3663;
  wire                _zz_dataOut_payload_0_3664;
  wire       [7:0]    _zz_dataOut_payload_0_3665;
  wire       [7:0]    _zz_dataOut_payload_0_3666;
  wire                _zz_dataOut_payload_0_3667;
  wire       [7:0]    _zz_dataOut_payload_0_3668;
  wire       [7:0]    _zz_dataOut_payload_0_3669;
  wire                _zz_dataOut_payload_0_3670;
  wire                _zz_dataOut_payload_0_3671;
  reg        [7:0]    _zz_dataOut_payload_0_3672;
  reg        [7:0]    _zz_dataOut_payload_0_3673;
  reg        [7:0]    _zz_dataOut_payload_0_3674;
  reg        [7:0]    _zz_dataOut_payload_0_3675;
  wire                _zz_dataOut_payload_0_3676;
  wire       [7:0]    _zz_dataOut_payload_0_3677;
  wire       [7:0]    _zz_dataOut_payload_0_3678;
  wire                _zz_dataOut_payload_0_3679;
  wire       [7:0]    _zz_dataOut_payload_0_3680;
  wire       [7:0]    _zz_dataOut_payload_0_3681;
  wire                _zz_dataOut_payload_0_3682;
  wire                _zz_dataOut_payload_0_3683;
  reg        [7:0]    _zz_dataOut_payload_0_3684;
  reg        [7:0]    _zz_dataOut_payload_0_3685;
  reg        [7:0]    _zz_dataOut_payload_0_3686;
  reg        [7:0]    _zz_dataOut_payload_0_3687;
  reg        [7:0]    _zz_dataOut_payload_0_3688;
  reg        [7:0]    _zz_dataOut_payload_0_3689;
  reg        [7:0]    _zz_dataOut_payload_0_3690;
  reg        [7:0]    _zz_dataOut_payload_0_3691;
  reg        [7:0]    _zz_dataOut_payload_0_3692;
  reg        [7:0]    _zz_dataOut_payload_0_3693;
  reg        [7:0]    _zz_dataOut_payload_0_3694;
  reg        [7:0]    _zz_dataOut_payload_0_3695;
  reg        [7:0]    _zz_dataOut_payload_0_3696;
  reg        [7:0]    _zz_dataOut_payload_0_3697;
  reg        [7:0]    _zz_dataOut_payload_0_3698;
  reg        [7:0]    _zz_dataOut_payload_0_3699;
  reg        [7:0]    _zz_dataOut_payload_0_3700;
  reg        [7:0]    _zz_dataOut_payload_0_3701;
  reg        [7:0]    _zz_dataOut_payload_0_3702;
  reg        [7:0]    _zz_dataOut_payload_0_3703;
  reg        [7:0]    _zz_dataOut_payload_0_3704;
  reg        [7:0]    _zz_dataOut_payload_0_3705;
  reg        [7:0]    _zz_dataOut_payload_0_3706;
  reg        [7:0]    _zz_dataOut_payload_0_3707;
  reg        [7:0]    _zz_dataOut_payload_0_3708;
  reg        [7:0]    _zz_dataOut_payload_0_3709;
  reg        [7:0]    _zz_dataOut_payload_0_3710;
  reg        [7:0]    _zz_dataOut_payload_0_3711;
  wire                _zz_dataOut_payload_0_3712;
  wire       [7:0]    _zz_dataOut_payload_0_3713;
  wire       [7:0]    _zz_dataOut_payload_0_3714;
  wire                _zz_dataOut_payload_0_3715;
  wire       [7:0]    _zz_dataOut_payload_0_3716;
  wire       [7:0]    _zz_dataOut_payload_0_3717;
  wire                _zz_dataOut_payload_0_3718;
  wire       [7:0]    _zz_dataOut_payload_0_3719;
  wire       [7:0]    _zz_dataOut_payload_0_3720;
  wire                _zz_dataOut_payload_0_3721;
  wire       [7:0]    _zz_dataOut_payload_0_3722;
  wire       [7:0]    _zz_dataOut_payload_0_3723;
  wire                _zz_dataOut_payload_0_3724;
  wire       [7:0]    _zz_dataOut_payload_0_3725;
  wire       [7:0]    _zz_dataOut_payload_0_3726;
  wire                _zz_dataOut_payload_0_3727;
  wire       [7:0]    _zz_dataOut_payload_0_3728;
  wire       [7:0]    _zz_dataOut_payload_0_3729;
  wire                _zz_dataOut_payload_0_3730;
  wire       [7:0]    _zz_dataOut_payload_0_3731;
  wire       [7:0]    _zz_dataOut_payload_0_3732;
  wire                _zz_dataOut_payload_0_3733;
  wire       [7:0]    _zz_dataOut_payload_0_3734;
  wire       [7:0]    _zz_dataOut_payload_0_3735;
  wire                _zz_dataOut_payload_0_3736;
  wire       [7:0]    _zz_dataOut_payload_0_3737;
  wire       [7:0]    _zz_dataOut_payload_0_3738;
  wire                _zz_dataOut_payload_0_3739;
  wire       [7:0]    _zz_dataOut_payload_0_3740;
  wire       [7:0]    _zz_dataOut_payload_0_3741;
  wire                _zz_dataOut_payload_0_3742;
  wire       [7:0]    _zz_dataOut_payload_0_3743;
  wire       [7:0]    _zz_dataOut_payload_0_3744;
  wire                _zz_dataOut_payload_0_3745;
  wire       [7:0]    _zz_dataOut_payload_0_3746;
  wire       [7:0]    _zz_dataOut_payload_0_3747;
  wire                _zz_dataOut_payload_0_3748;
  wire       [7:0]    _zz_dataOut_payload_0_3749;
  wire       [7:0]    _zz_dataOut_payload_0_3750;
  wire                _zz_dataOut_payload_0_3751;
  wire       [7:0]    _zz_dataOut_payload_0_3752;
  wire       [7:0]    _zz_dataOut_payload_0_3753;
  wire                _zz_dataOut_payload_0_3754;
  wire                _zz_dataOut_payload_0_3755;
  reg        [7:0]    _zz_dataOut_payload_0_3756;
  reg        [7:0]    _zz_dataOut_payload_0_3757;
  reg        [7:0]    _zz_dataOut_payload_0_3758;
  reg        [7:0]    _zz_dataOut_payload_0_3759;
  wire                _zz_dataOut_payload_0_3760;
  wire       [7:0]    _zz_dataOut_payload_0_3761;
  wire       [7:0]    _zz_dataOut_payload_0_3762;
  wire                _zz_dataOut_payload_0_3763;
  wire       [7:0]    _zz_dataOut_payload_0_3764;
  wire       [7:0]    _zz_dataOut_payload_0_3765;
  wire                _zz_dataOut_payload_0_3766;
  wire                _zz_dataOut_payload_0_3767;
  reg        [7:0]    _zz_dataOut_payload_0_3768;
  reg        [7:0]    _zz_dataOut_payload_0_3769;
  reg        [7:0]    _zz_dataOut_payload_0_3770;
  reg        [7:0]    _zz_dataOut_payload_0_3771;
  reg        [7:0]    _zz_dataOut_payload_0_3772;
  reg        [7:0]    _zz_dataOut_payload_0_3773;
  reg        [7:0]    _zz_dataOut_payload_0_3774;
  reg        [7:0]    _zz_dataOut_payload_0_3775;
  reg        [7:0]    _zz_dataOut_payload_0_3776;
  reg        [7:0]    _zz_dataOut_payload_0_3777;
  reg        [7:0]    _zz_dataOut_payload_0_3778;
  reg        [7:0]    _zz_dataOut_payload_0_3779;
  wire                _zz_dataOut_payload_0_3780;
  wire       [7:0]    _zz_dataOut_payload_0_3781;
  wire       [7:0]    _zz_dataOut_payload_0_3782;
  wire                _zz_dataOut_payload_0_3783;
  wire       [7:0]    _zz_dataOut_payload_0_3784;
  wire       [7:0]    _zz_dataOut_payload_0_3785;
  wire                _zz_dataOut_payload_0_3786;
  wire       [7:0]    _zz_dataOut_payload_0_3787;
  wire       [7:0]    _zz_dataOut_payload_0_3788;
  wire                _zz_dataOut_payload_0_3789;
  wire       [7:0]    _zz_dataOut_payload_0_3790;
  wire       [7:0]    _zz_dataOut_payload_0_3791;
  wire                _zz_dataOut_payload_0_3792;
  wire       [7:0]    _zz_dataOut_payload_0_3793;
  wire       [7:0]    _zz_dataOut_payload_0_3794;
  wire                _zz_dataOut_payload_0_3795;
  wire       [7:0]    _zz_dataOut_payload_0_3796;
  wire       [7:0]    _zz_dataOut_payload_0_3797;
  wire                _zz_dataOut_payload_0_3798;
  wire                _zz_dataOut_payload_0_3799;
  reg        [7:0]    _zz_dataOut_payload_0_3800;
  reg        [7:0]    _zz_dataOut_payload_0_3801;
  reg        [7:0]    _zz_dataOut_payload_0_3802;
  reg        [7:0]    _zz_dataOut_payload_0_3803;
  wire                _zz_dataOut_payload_0_3804;
  wire       [7:0]    _zz_dataOut_payload_0_3805;
  wire       [7:0]    _zz_dataOut_payload_0_3806;
  wire                _zz_dataOut_payload_0_3807;
  wire       [7:0]    _zz_dataOut_payload_0_3808;
  wire       [7:0]    _zz_dataOut_payload_0_3809;
  wire                _zz_dataOut_payload_0_3810;
  wire                _zz_dataOut_payload_0_3811;
  reg        [7:0]    _zz_dataOut_payload_0_3812;
  reg        [7:0]    _zz_dataOut_payload_0_3813;
  reg        [7:0]    _zz_dataOut_payload_0_3814;
  reg        [7:0]    _zz_dataOut_payload_0_3815;
  reg        [7:0]    _zz_dataOut_payload_0_3816;
  reg        [7:0]    _zz_dataOut_payload_0_3817;
  reg        [7:0]    _zz_dataOut_payload_0_3818;
  reg        [7:0]    _zz_dataOut_payload_0_3819;
  reg        [7:0]    _zz_dataOut_payload_0_3820;
  reg        [7:0]    _zz_dataOut_payload_0_3821;
  reg        [7:0]    _zz_dataOut_payload_0_3822;
  reg        [7:0]    _zz_dataOut_payload_0_3823;
  reg        [7:0]    _zz_dataOut_payload_0_3824;
  reg        [7:0]    _zz_dataOut_payload_0_3825;
  reg        [7:0]    _zz_dataOut_payload_0_3826;
  reg        [7:0]    _zz_dataOut_payload_0_3827;
  reg        [7:0]    _zz_dataOut_payload_0_3828;
  reg        [7:0]    _zz_dataOut_payload_0_3829;
  reg        [7:0]    _zz_dataOut_payload_0_3830;
  reg        [7:0]    _zz_dataOut_payload_0_3831;
  reg        [7:0]    _zz_dataOut_payload_0_3832;
  reg        [7:0]    _zz_dataOut_payload_0_3833;
  reg        [7:0]    _zz_dataOut_payload_0_3834;
  reg        [7:0]    _zz_dataOut_payload_0_3835;
  reg        [7:0]    _zz_dataOut_payload_0_3836;
  reg        [7:0]    _zz_dataOut_payload_0_3837;
  reg        [7:0]    _zz_dataOut_payload_0_3838;
  reg        [7:0]    _zz_dataOut_payload_0_3839;
  wire                _zz_dataOut_payload_0_3840;
  wire       [7:0]    _zz_dataOut_payload_0_3841;
  wire       [7:0]    _zz_dataOut_payload_0_3842;
  wire                _zz_dataOut_payload_0_3843;
  wire       [7:0]    _zz_dataOut_payload_0_3844;
  wire       [7:0]    _zz_dataOut_payload_0_3845;
  wire                _zz_dataOut_payload_0_3846;
  wire       [7:0]    _zz_dataOut_payload_0_3847;
  wire       [7:0]    _zz_dataOut_payload_0_3848;
  wire                _zz_dataOut_payload_0_3849;
  wire       [7:0]    _zz_dataOut_payload_0_3850;
  wire       [7:0]    _zz_dataOut_payload_0_3851;
  wire                _zz_dataOut_payload_0_3852;
  wire       [7:0]    _zz_dataOut_payload_0_3853;
  wire       [7:0]    _zz_dataOut_payload_0_3854;
  wire                _zz_dataOut_payload_0_3855;
  wire       [7:0]    _zz_dataOut_payload_0_3856;
  wire       [7:0]    _zz_dataOut_payload_0_3857;
  wire                _zz_dataOut_payload_0_3858;
  wire       [7:0]    _zz_dataOut_payload_0_3859;
  wire       [7:0]    _zz_dataOut_payload_0_3860;
  wire                _zz_dataOut_payload_0_3861;
  wire       [7:0]    _zz_dataOut_payload_0_3862;
  wire       [7:0]    _zz_dataOut_payload_0_3863;
  wire                _zz_dataOut_payload_0_3864;
  wire       [7:0]    _zz_dataOut_payload_0_3865;
  wire       [7:0]    _zz_dataOut_payload_0_3866;
  wire                _zz_dataOut_payload_0_3867;
  wire       [7:0]    _zz_dataOut_payload_0_3868;
  wire       [7:0]    _zz_dataOut_payload_0_3869;
  wire                _zz_dataOut_payload_0_3870;
  wire       [7:0]    _zz_dataOut_payload_0_3871;
  wire       [7:0]    _zz_dataOut_payload_0_3872;
  wire                _zz_dataOut_payload_0_3873;
  wire       [7:0]    _zz_dataOut_payload_0_3874;
  wire       [7:0]    _zz_dataOut_payload_0_3875;
  wire                _zz_dataOut_payload_0_3876;
  wire       [7:0]    _zz_dataOut_payload_0_3877;
  wire       [7:0]    _zz_dataOut_payload_0_3878;
  wire                _zz_dataOut_payload_0_3879;
  wire       [7:0]    _zz_dataOut_payload_0_3880;
  wire       [7:0]    _zz_dataOut_payload_0_3881;
  wire                _zz_dataOut_payload_0_3882;
  wire                _zz_dataOut_payload_0_3883;
  reg        [7:0]    _zz_dataOut_payload_0_3884;
  reg        [7:0]    _zz_dataOut_payload_0_3885;
  reg        [7:0]    _zz_dataOut_payload_0_3886;
  reg        [7:0]    _zz_dataOut_payload_0_3887;
  wire                _zz_dataOut_payload_0_3888;
  wire       [7:0]    _zz_dataOut_payload_0_3889;
  wire       [7:0]    _zz_dataOut_payload_0_3890;
  wire                _zz_dataOut_payload_0_3891;
  wire       [7:0]    _zz_dataOut_payload_0_3892;
  wire       [7:0]    _zz_dataOut_payload_0_3893;
  wire                _zz_dataOut_payload_0_3894;
  wire                _zz_dataOut_payload_0_3895;
  reg        [7:0]    _zz_dataOut_payload_0_3896;
  reg        [7:0]    _zz_dataOut_payload_0_3897;
  reg        [7:0]    _zz_dataOut_payload_0_3898;
  reg        [7:0]    _zz_dataOut_payload_0_3899;
  reg        [7:0]    _zz_dataOut_payload_0_3900;
  reg        [7:0]    _zz_dataOut_payload_0_3901;
  reg        [7:0]    _zz_dataOut_payload_0_3902;
  reg        [7:0]    _zz_dataOut_payload_0_3903;
  reg        [7:0]    _zz_dataOut_payload_0_3904;
  reg        [7:0]    _zz_dataOut_payload_0_3905;
  reg        [7:0]    _zz_dataOut_payload_0_3906;
  reg        [7:0]    _zz_dataOut_payload_0_3907;
  wire                _zz_dataOut_payload_0_3908;
  wire       [7:0]    _zz_dataOut_payload_0_3909;
  wire       [7:0]    _zz_dataOut_payload_0_3910;
  wire                _zz_dataOut_payload_0_3911;
  wire       [7:0]    _zz_dataOut_payload_0_3912;
  wire       [7:0]    _zz_dataOut_payload_0_3913;
  wire                _zz_dataOut_payload_0_3914;
  wire       [7:0]    _zz_dataOut_payload_0_3915;
  wire       [7:0]    _zz_dataOut_payload_0_3916;
  wire                _zz_dataOut_payload_0_3917;
  wire       [7:0]    _zz_dataOut_payload_0_3918;
  wire       [7:0]    _zz_dataOut_payload_0_3919;
  wire                _zz_dataOut_payload_0_3920;
  wire       [7:0]    _zz_dataOut_payload_0_3921;
  wire       [7:0]    _zz_dataOut_payload_0_3922;
  wire                _zz_dataOut_payload_0_3923;
  wire       [7:0]    _zz_dataOut_payload_0_3924;
  wire       [7:0]    _zz_dataOut_payload_0_3925;
  wire                _zz_dataOut_payload_0_3926;
  wire                _zz_dataOut_payload_0_3927;
  reg        [7:0]    _zz_dataOut_payload_0_3928;
  reg        [7:0]    _zz_dataOut_payload_0_3929;
  reg        [7:0]    _zz_dataOut_payload_0_3930;
  reg        [7:0]    _zz_dataOut_payload_0_3931;
  wire                _zz_dataOut_payload_0_3932;
  wire       [7:0]    _zz_dataOut_payload_0_3933;
  wire       [7:0]    _zz_dataOut_payload_0_3934;
  wire                _zz_dataOut_payload_0_3935;
  wire       [7:0]    _zz_dataOut_payload_0_3936;
  wire       [7:0]    _zz_dataOut_payload_0_3937;
  wire                _zz_dataOut_payload_0_3938;
  wire                _zz_dataOut_payload_0_3939;
  reg        [7:0]    _zz_dataOut_payload_0_3940;
  reg        [7:0]    _zz_dataOut_payload_0_3941;
  reg        [7:0]    _zz_dataOut_payload_0_3942;
  reg        [7:0]    _zz_dataOut_payload_0_3943;
  reg        [7:0]    _zz_dataOut_payload_0_3944;
  reg        [7:0]    _zz_dataOut_payload_0_3945;
  reg        [7:0]    _zz_dataOut_payload_0_3946;
  reg        [7:0]    _zz_dataOut_payload_0_3947;
  reg        [7:0]    _zz_dataOut_payload_0_3948;
  reg        [7:0]    _zz_dataOut_payload_0_3949;
  reg        [7:0]    _zz_dataOut_payload_0_3950;
  reg        [7:0]    _zz_dataOut_payload_0_3951;
  reg        [7:0]    _zz_dataOut_payload_0_3952;
  reg        [7:0]    _zz_dataOut_payload_0_3953;
  reg        [7:0]    _zz_dataOut_payload_0_3954;
  reg        [7:0]    _zz_dataOut_payload_0_3955;
  reg        [7:0]    _zz_dataOut_payload_0_3956;
  reg        [7:0]    _zz_dataOut_payload_0_3957;
  reg        [7:0]    _zz_dataOut_payload_0_3958;
  reg        [7:0]    _zz_dataOut_payload_0_3959;
  reg        [7:0]    _zz_dataOut_payload_0_3960;
  reg        [7:0]    _zz_dataOut_payload_0_3961;
  reg        [7:0]    _zz_dataOut_payload_0_3962;
  reg        [7:0]    _zz_dataOut_payload_0_3963;
  reg        [7:0]    _zz_dataOut_payload_0_3964;
  reg        [7:0]    _zz_dataOut_payload_0_3965;
  reg        [7:0]    _zz_dataOut_payload_0_3966;
  reg        [7:0]    _zz_dataOut_payload_0_3967;
  wire                _zz_dataOut_payload_0_3968;
  wire       [7:0]    _zz_dataOut_payload_0_3969;
  wire       [7:0]    _zz_dataOut_payload_0_3970;
  wire                _zz_dataOut_payload_0_3971;
  wire       [7:0]    _zz_dataOut_payload_0_3972;
  wire       [7:0]    _zz_dataOut_payload_0_3973;
  wire                _zz_dataOut_payload_0_3974;
  wire       [7:0]    _zz_dataOut_payload_0_3975;
  wire       [7:0]    _zz_dataOut_payload_0_3976;
  wire                _zz_dataOut_payload_0_3977;
  wire       [7:0]    _zz_dataOut_payload_0_3978;
  wire       [7:0]    _zz_dataOut_payload_0_3979;
  wire                _zz_dataOut_payload_0_3980;
  wire       [7:0]    _zz_dataOut_payload_0_3981;
  wire       [7:0]    _zz_dataOut_payload_0_3982;
  wire                _zz_dataOut_payload_0_3983;
  wire       [7:0]    _zz_dataOut_payload_0_3984;
  wire       [7:0]    _zz_dataOut_payload_0_3985;
  wire                _zz_dataOut_payload_0_3986;
  wire       [7:0]    _zz_dataOut_payload_0_3987;
  wire       [7:0]    _zz_dataOut_payload_0_3988;
  wire                _zz_dataOut_payload_0_3989;
  wire       [7:0]    _zz_dataOut_payload_0_3990;
  wire       [7:0]    _zz_dataOut_payload_0_3991;
  wire                _zz_dataOut_payload_0_3992;
  wire       [7:0]    _zz_dataOut_payload_0_3993;
  wire       [7:0]    _zz_dataOut_payload_0_3994;
  wire                _zz_dataOut_payload_0_3995;
  wire       [7:0]    _zz_dataOut_payload_0_3996;
  wire       [7:0]    _zz_dataOut_payload_0_3997;
  wire                _zz_dataOut_payload_0_3998;
  wire       [7:0]    _zz_dataOut_payload_0_3999;
  wire       [7:0]    _zz_dataOut_payload_0_4000;
  wire                _zz_dataOut_payload_0_4001;
  wire       [7:0]    _zz_dataOut_payload_0_4002;
  wire       [7:0]    _zz_dataOut_payload_0_4003;
  wire                _zz_dataOut_payload_0_4004;
  wire       [7:0]    _zz_dataOut_payload_0_4005;
  wire       [7:0]    _zz_dataOut_payload_0_4006;
  wire                _zz_dataOut_payload_0_4007;
  wire       [7:0]    _zz_dataOut_payload_0_4008;
  wire       [7:0]    _zz_dataOut_payload_0_4009;
  wire                _zz_dataOut_payload_0_4010;
  wire                _zz_dataOut_payload_0_4011;
  reg        [7:0]    _zz_dataOut_payload_0_4012;
  reg        [7:0]    _zz_dataOut_payload_0_4013;
  reg        [7:0]    _zz_dataOut_payload_0_4014;
  reg        [7:0]    _zz_dataOut_payload_0_4015;
  wire                _zz_dataOut_payload_0_4016;
  wire       [7:0]    _zz_dataOut_payload_0_4017;
  wire       [7:0]    _zz_dataOut_payload_0_4018;
  wire                _zz_dataOut_payload_0_4019;
  wire       [7:0]    _zz_dataOut_payload_0_4020;
  wire       [7:0]    _zz_dataOut_payload_0_4021;
  wire                _zz_dataOut_payload_0_4022;
  wire                _zz_dataOut_payload_0_4023;
  reg        [7:0]    _zz_dataOut_payload_0_4024;
  reg        [7:0]    _zz_dataOut_payload_0_4025;
  reg        [7:0]    _zz_dataOut_payload_0_4026;
  reg        [7:0]    _zz_dataOut_payload_0_4027;
  reg        [7:0]    _zz_dataOut_payload_0_4028;
  reg        [7:0]    _zz_dataOut_payload_0_4029;
  reg        [7:0]    _zz_dataOut_payload_0_4030;
  reg        [7:0]    _zz_dataOut_payload_0_4031;
  reg        [7:0]    _zz_dataOut_payload_0_4032;
  reg        [7:0]    _zz_dataOut_payload_0_4033;
  reg        [7:0]    _zz_dataOut_payload_0_4034;
  reg        [7:0]    _zz_dataOut_payload_0_4035;
  wire                _zz_dataOut_payload_0_4036;
  wire       [7:0]    _zz_dataOut_payload_0_4037;
  wire       [7:0]    _zz_dataOut_payload_0_4038;
  wire                _zz_dataOut_payload_0_4039;
  wire       [7:0]    _zz_dataOut_payload_0_4040;
  wire       [7:0]    _zz_dataOut_payload_0_4041;
  wire                _zz_dataOut_payload_0_4042;
  wire       [7:0]    _zz_dataOut_payload_0_4043;
  wire       [7:0]    _zz_dataOut_payload_0_4044;
  wire                _zz_dataOut_payload_0_4045;
  wire       [7:0]    _zz_dataOut_payload_0_4046;
  wire       [7:0]    _zz_dataOut_payload_0_4047;
  wire                _zz_dataOut_payload_0_4048;
  wire       [7:0]    _zz_dataOut_payload_0_4049;
  wire       [7:0]    _zz_dataOut_payload_0_4050;
  wire                _zz_dataOut_payload_0_4051;
  wire       [7:0]    _zz_dataOut_payload_0_4052;
  wire       [7:0]    _zz_dataOut_payload_0_4053;
  wire                _zz_dataOut_payload_0_4054;
  wire                _zz_dataOut_payload_0_4055;
  reg        [7:0]    _zz_dataOut_payload_0_4056;
  reg        [7:0]    _zz_dataOut_payload_0_4057;
  reg        [7:0]    _zz_dataOut_payload_0_4058;
  reg        [7:0]    _zz_dataOut_payload_0_4059;
  wire                _zz_dataOut_payload_0_4060;
  wire       [7:0]    _zz_dataOut_payload_0_4061;
  wire       [7:0]    _zz_dataOut_payload_0_4062;
  wire                _zz_dataOut_payload_0_4063;
  wire       [7:0]    _zz_dataOut_payload_0_4064;
  wire       [7:0]    _zz_dataOut_payload_0_4065;
  wire                _zz_dataOut_payload_0_4066;
  wire                _zz_dataOut_payload_0_4067;
  reg        [7:0]    _zz_dataOut_payload_0_4068;
  reg        [7:0]    _zz_dataOut_payload_0_4069;
  reg        [7:0]    _zz_dataOut_payload_0_4070;
  reg        [7:0]    _zz_dataOut_payload_0_4071;
  reg        [7:0]    _zz_dataOut_payload_0_4072;
  reg        [7:0]    _zz_dataOut_payload_0_4073;
  reg        [7:0]    _zz_dataOut_payload_0_4074;
  reg        [7:0]    _zz_dataOut_payload_0_4075;
  reg        [7:0]    _zz_dataOut_payload_0_4076;
  reg        [7:0]    _zz_dataOut_payload_0_4077;
  reg        [7:0]    _zz_dataOut_payload_0_4078;
  reg        [7:0]    _zz_dataOut_payload_0_4079;
  reg        [7:0]    _zz_dataOut_payload_0_4080;
  reg        [7:0]    _zz_dataOut_payload_0_4081;
  reg        [7:0]    _zz_dataOut_payload_0_4082;
  reg        [7:0]    _zz_dataOut_payload_0_4083;
  reg        [7:0]    _zz_dataOut_payload_0_4084;
  reg        [7:0]    _zz_dataOut_payload_0_4085;
  reg        [7:0]    _zz_dataOut_payload_0_4086;
  reg        [7:0]    _zz_dataOut_payload_0_4087;
  reg        [7:0]    _zz_dataOut_payload_0_4088;
  reg        [7:0]    _zz_dataOut_payload_0_4089;
  reg        [7:0]    _zz_dataOut_payload_0_4090;
  reg        [7:0]    _zz_dataOut_payload_0_4091;
  reg        [7:0]    _zz_dataOut_payload_0_4092;
  reg        [7:0]    _zz_dataOut_payload_0_4093;
  reg        [7:0]    _zz_dataOut_payload_0_4094;
  reg        [7:0]    _zz_dataOut_payload_0_4095;
  wire                _zz_dataOut_payload_0_4096;
  wire       [7:0]    _zz_dataOut_payload_0_4097;
  wire       [7:0]    _zz_dataOut_payload_0_4098;
  wire                _zz_dataOut_payload_0_4099;
  wire       [7:0]    _zz_dataOut_payload_0_4100;
  wire       [7:0]    _zz_dataOut_payload_0_4101;
  wire                _zz_dataOut_payload_0_4102;
  wire       [7:0]    _zz_dataOut_payload_0_4103;
  wire       [7:0]    _zz_dataOut_payload_0_4104;
  wire                _zz_dataOut_payload_0_4105;
  wire       [7:0]    _zz_dataOut_payload_0_4106;
  wire       [7:0]    _zz_dataOut_payload_0_4107;
  wire                _zz_dataOut_payload_0_4108;
  wire       [7:0]    _zz_dataOut_payload_0_4109;
  wire       [7:0]    _zz_dataOut_payload_0_4110;
  wire                _zz_dataOut_payload_0_4111;
  wire       [7:0]    _zz_dataOut_payload_0_4112;
  wire       [7:0]    _zz_dataOut_payload_0_4113;
  wire                _zz_dataOut_payload_0_4114;
  wire       [7:0]    _zz_dataOut_payload_0_4115;
  wire       [7:0]    _zz_dataOut_payload_0_4116;
  wire                _zz_dataOut_payload_0_4117;
  wire       [7:0]    _zz_dataOut_payload_0_4118;
  wire       [7:0]    _zz_dataOut_payload_0_4119;
  wire                _zz_dataOut_payload_0_4120;
  wire       [7:0]    _zz_dataOut_payload_0_4121;
  wire       [7:0]    _zz_dataOut_payload_0_4122;
  wire                _zz_dataOut_payload_0_4123;
  wire       [7:0]    _zz_dataOut_payload_0_4124;
  wire       [7:0]    _zz_dataOut_payload_0_4125;
  wire                _zz_dataOut_payload_0_4126;
  wire       [7:0]    _zz_dataOut_payload_0_4127;
  wire       [7:0]    _zz_dataOut_payload_0_4128;
  wire                _zz_dataOut_payload_0_4129;
  wire       [7:0]    _zz_dataOut_payload_0_4130;
  wire       [7:0]    _zz_dataOut_payload_0_4131;
  wire                _zz_dataOut_payload_0_4132;
  wire       [7:0]    _zz_dataOut_payload_0_4133;
  wire       [7:0]    _zz_dataOut_payload_0_4134;
  wire                _zz_dataOut_payload_0_4135;
  wire       [7:0]    _zz_dataOut_payload_0_4136;
  wire       [7:0]    _zz_dataOut_payload_0_4137;
  wire                _zz_dataOut_payload_0_4138;
  wire                _zz_dataOut_payload_0_4139;
  reg        [7:0]    _zz_dataOut_payload_0_4140;
  reg        [7:0]    _zz_dataOut_payload_0_4141;
  reg        [7:0]    _zz_dataOut_payload_0_4142;
  reg        [7:0]    _zz_dataOut_payload_0_4143;
  wire                _zz_dataOut_payload_0_4144;
  wire       [7:0]    _zz_dataOut_payload_0_4145;
  wire       [7:0]    _zz_dataOut_payload_0_4146;
  wire                _zz_dataOut_payload_0_4147;
  wire       [7:0]    _zz_dataOut_payload_0_4148;
  wire       [7:0]    _zz_dataOut_payload_0_4149;
  wire                _zz_dataOut_payload_0_4150;
  wire                _zz_dataOut_payload_0_4151;
  reg        [7:0]    _zz_dataOut_payload_0_4152;
  reg        [7:0]    _zz_dataOut_payload_0_4153;
  reg        [7:0]    _zz_dataOut_payload_0_4154;
  reg        [7:0]    _zz_dataOut_payload_0_4155;
  reg        [7:0]    _zz_dataOut_payload_0_4156;
  reg        [7:0]    _zz_dataOut_payload_0_4157;
  reg        [7:0]    _zz_dataOut_payload_0_4158;
  reg        [7:0]    _zz_dataOut_payload_0_4159;
  reg        [7:0]    _zz_dataOut_payload_0_4160;
  reg        [7:0]    _zz_dataOut_payload_0_4161;
  reg        [7:0]    _zz_dataOut_payload_0_4162;
  reg        [7:0]    _zz_dataOut_payload_0_4163;
  wire                _zz_dataOut_payload_0_4164;
  wire       [7:0]    _zz_dataOut_payload_0_4165;
  wire       [7:0]    _zz_dataOut_payload_0_4166;
  wire                _zz_dataOut_payload_0_4167;
  wire       [7:0]    _zz_dataOut_payload_0_4168;
  wire       [7:0]    _zz_dataOut_payload_0_4169;
  wire                _zz_dataOut_payload_0_4170;
  wire       [7:0]    _zz_dataOut_payload_0_4171;
  wire       [7:0]    _zz_dataOut_payload_0_4172;
  wire                _zz_dataOut_payload_0_4173;
  wire       [7:0]    _zz_dataOut_payload_0_4174;
  wire       [7:0]    _zz_dataOut_payload_0_4175;
  wire                _zz_dataOut_payload_0_4176;
  wire       [7:0]    _zz_dataOut_payload_0_4177;
  wire       [7:0]    _zz_dataOut_payload_0_4178;
  wire                _zz_dataOut_payload_0_4179;
  wire       [7:0]    _zz_dataOut_payload_0_4180;
  wire       [7:0]    _zz_dataOut_payload_0_4181;
  wire                _zz_dataOut_payload_0_4182;
  wire                _zz_dataOut_payload_0_4183;
  reg        [7:0]    _zz_dataOut_payload_0_4184;
  reg        [7:0]    _zz_dataOut_payload_0_4185;
  reg        [7:0]    _zz_dataOut_payload_0_4186;
  reg        [7:0]    _zz_dataOut_payload_0_4187;
  wire                _zz_dataOut_payload_0_4188;
  wire       [7:0]    _zz_dataOut_payload_0_4189;
  wire       [7:0]    _zz_dataOut_payload_0_4190;
  wire                _zz_dataOut_payload_0_4191;
  wire       [7:0]    _zz_dataOut_payload_0_4192;
  wire       [7:0]    _zz_dataOut_payload_0_4193;
  wire                _zz_dataOut_payload_0_4194;
  wire                _zz_dataOut_payload_0_4195;
  reg        [7:0]    _zz_dataOut_payload_0_4196;
  reg        [7:0]    _zz_dataOut_payload_0_4197;
  reg        [7:0]    _zz_dataOut_payload_0_4198;
  reg        [7:0]    _zz_dataOut_payload_0_4199;
  reg        [7:0]    _zz_dataOut_payload_0_4200;
  reg        [7:0]    _zz_dataOut_payload_0_4201;
  reg        [7:0]    _zz_dataOut_payload_0_4202;
  reg        [7:0]    _zz_dataOut_payload_0_4203;
  reg        [7:0]    _zz_dataOut_payload_0_4204;
  reg        [7:0]    _zz_dataOut_payload_0_4205;
  reg        [7:0]    _zz_dataOut_payload_0_4206;
  reg        [7:0]    _zz_dataOut_payload_0_4207;
  reg        [7:0]    _zz_dataOut_payload_0_4208;
  reg        [7:0]    _zz_dataOut_payload_0_4209;
  reg        [7:0]    _zz_dataOut_payload_0_4210;
  reg        [7:0]    _zz_dataOut_payload_0_4211;
  reg        [7:0]    _zz_dataOut_payload_0_4212;
  reg        [7:0]    _zz_dataOut_payload_0_4213;
  reg        [7:0]    _zz_dataOut_payload_0_4214;
  reg        [7:0]    _zz_dataOut_payload_0_4215;
  reg        [7:0]    _zz_dataOut_payload_0_4216;
  reg        [7:0]    _zz_dataOut_payload_0_4217;
  reg        [7:0]    _zz_dataOut_payload_0_4218;
  reg        [7:0]    _zz_dataOut_payload_0_4219;
  reg        [7:0]    _zz_dataOut_payload_0_4220;
  reg        [7:0]    _zz_dataOut_payload_0_4221;
  reg        [7:0]    _zz_dataOut_payload_0_4222;
  reg        [7:0]    _zz_dataOut_payload_0_4223;
  wire                _zz_dataOut_payload_0_4224;
  wire       [7:0]    _zz_dataOut_payload_0_4225;
  wire       [7:0]    _zz_dataOut_payload_0_4226;
  wire                _zz_dataOut_payload_0_4227;
  wire       [7:0]    _zz_dataOut_payload_0_4228;
  wire       [7:0]    _zz_dataOut_payload_0_4229;
  wire                _zz_dataOut_payload_0_4230;
  wire       [7:0]    _zz_dataOut_payload_0_4231;
  wire       [7:0]    _zz_dataOut_payload_0_4232;
  wire                _zz_dataOut_payload_0_4233;
  wire       [7:0]    _zz_dataOut_payload_0_4234;
  wire       [7:0]    _zz_dataOut_payload_0_4235;
  wire                _zz_dataOut_payload_0_4236;
  wire       [7:0]    _zz_dataOut_payload_0_4237;
  wire       [7:0]    _zz_dataOut_payload_0_4238;
  wire                _zz_dataOut_payload_0_4239;
  wire       [7:0]    _zz_dataOut_payload_0_4240;
  wire       [7:0]    _zz_dataOut_payload_0_4241;
  wire                _zz_dataOut_payload_0_4242;
  wire       [7:0]    _zz_dataOut_payload_0_4243;
  wire       [7:0]    _zz_dataOut_payload_0_4244;
  wire                _zz_dataOut_payload_0_4245;
  wire       [7:0]    _zz_dataOut_payload_0_4246;
  wire       [7:0]    _zz_dataOut_payload_0_4247;
  wire                _zz_dataOut_payload_0_4248;
  wire       [7:0]    _zz_dataOut_payload_0_4249;
  wire       [7:0]    _zz_dataOut_payload_0_4250;
  wire                _zz_dataOut_payload_0_4251;
  wire       [7:0]    _zz_dataOut_payload_0_4252;
  wire       [7:0]    _zz_dataOut_payload_0_4253;
  wire                _zz_dataOut_payload_0_4254;
  wire       [7:0]    _zz_dataOut_payload_0_4255;
  wire       [7:0]    _zz_dataOut_payload_0_4256;
  wire                _zz_dataOut_payload_0_4257;
  wire       [7:0]    _zz_dataOut_payload_0_4258;
  wire       [7:0]    _zz_dataOut_payload_0_4259;
  wire                _zz_dataOut_payload_0_4260;
  wire       [7:0]    _zz_dataOut_payload_0_4261;
  wire       [7:0]    _zz_dataOut_payload_0_4262;
  wire                _zz_dataOut_payload_0_4263;
  wire       [7:0]    _zz_dataOut_payload_0_4264;
  wire       [7:0]    _zz_dataOut_payload_0_4265;
  wire                _zz_dataOut_payload_0_4266;
  wire                _zz_dataOut_payload_0_4267;
  reg        [7:0]    _zz_dataOut_payload_0_4268;
  reg        [7:0]    _zz_dataOut_payload_0_4269;
  reg        [7:0]    _zz_dataOut_payload_0_4270;
  reg        [7:0]    _zz_dataOut_payload_0_4271;
  wire                _zz_dataOut_payload_0_4272;
  wire       [7:0]    _zz_dataOut_payload_0_4273;
  wire       [7:0]    _zz_dataOut_payload_0_4274;
  wire                _zz_dataOut_payload_0_4275;
  wire       [7:0]    _zz_dataOut_payload_0_4276;
  wire       [7:0]    _zz_dataOut_payload_0_4277;
  wire                _zz_dataOut_payload_0_4278;
  wire                _zz_dataOut_payload_0_4279;
  reg        [7:0]    _zz_dataOut_payload_0_4280;
  reg        [7:0]    _zz_dataOut_payload_0_4281;
  reg        [7:0]    _zz_dataOut_payload_0_4282;
  reg        [7:0]    _zz_dataOut_payload_0_4283;
  reg        [7:0]    _zz_dataOut_payload_0_4284;
  reg        [7:0]    _zz_dataOut_payload_0_4285;
  reg        [7:0]    _zz_dataOut_payload_0_4286;
  reg        [7:0]    _zz_dataOut_payload_0_4287;
  reg        [7:0]    _zz_dataOut_payload_0_4288;
  reg        [7:0]    _zz_dataOut_payload_0_4289;
  reg        [7:0]    _zz_dataOut_payload_0_4290;
  reg        [7:0]    _zz_dataOut_payload_0_4291;
  wire                _zz_dataOut_payload_0_4292;
  wire       [7:0]    _zz_dataOut_payload_0_4293;
  wire       [7:0]    _zz_dataOut_payload_0_4294;
  wire                _zz_dataOut_payload_0_4295;
  wire       [7:0]    _zz_dataOut_payload_0_4296;
  wire       [7:0]    _zz_dataOut_payload_0_4297;
  wire                _zz_dataOut_payload_0_4298;
  wire       [7:0]    _zz_dataOut_payload_0_4299;
  wire       [7:0]    _zz_dataOut_payload_0_4300;
  wire                _zz_dataOut_payload_0_4301;
  wire       [7:0]    _zz_dataOut_payload_0_4302;
  wire       [7:0]    _zz_dataOut_payload_0_4303;
  wire                _zz_dataOut_payload_0_4304;
  wire       [7:0]    _zz_dataOut_payload_0_4305;
  wire       [7:0]    _zz_dataOut_payload_0_4306;
  wire                _zz_dataOut_payload_0_4307;
  wire       [7:0]    _zz_dataOut_payload_0_4308;
  wire       [7:0]    _zz_dataOut_payload_0_4309;
  wire                _zz_dataOut_payload_0_4310;
  wire                _zz_dataOut_payload_0_4311;
  reg        [7:0]    _zz_dataOut_payload_0_4312;
  reg        [7:0]    _zz_dataOut_payload_0_4313;
  reg        [7:0]    _zz_dataOut_payload_0_4314;
  reg        [7:0]    _zz_dataOut_payload_0_4315;
  wire                _zz_dataOut_payload_0_4316;
  wire       [7:0]    _zz_dataOut_payload_0_4317;
  wire       [7:0]    _zz_dataOut_payload_0_4318;
  wire                _zz_dataOut_payload_0_4319;
  wire       [7:0]    _zz_dataOut_payload_0_4320;
  wire       [7:0]    _zz_dataOut_payload_0_4321;
  wire                _zz_dataOut_payload_0_4322;
  wire                _zz_dataOut_payload_0_4323;
  reg        [7:0]    _zz_dataOut_payload_0_4324;
  reg        [7:0]    _zz_dataOut_payload_0_4325;
  reg        [7:0]    _zz_dataOut_payload_0_4326;
  reg        [7:0]    _zz_dataOut_payload_0_4327;
  reg        [7:0]    _zz_dataOut_payload_0_4328;
  reg        [7:0]    _zz_dataOut_payload_0_4329;
  reg        [7:0]    _zz_dataOut_payload_0_4330;
  reg        [7:0]    _zz_dataOut_payload_0_4331;
  reg        [7:0]    _zz_dataOut_payload_0_4332;
  reg        [7:0]    _zz_dataOut_payload_0_4333;
  reg        [7:0]    _zz_dataOut_payload_0_4334;
  reg        [7:0]    _zz_dataOut_payload_0_4335;
  reg        [7:0]    _zz_dataOut_payload_0_4336;
  reg        [7:0]    _zz_dataOut_payload_0_4337;
  reg        [7:0]    _zz_dataOut_payload_0_4338;
  reg        [7:0]    _zz_dataOut_payload_0_4339;
  reg        [7:0]    _zz_dataOut_payload_0_4340;
  reg        [7:0]    _zz_dataOut_payload_0_4341;
  reg        [7:0]    _zz_dataOut_payload_0_4342;
  reg        [7:0]    _zz_dataOut_payload_0_4343;
  reg        [7:0]    _zz_dataOut_payload_0_4344;
  reg        [7:0]    _zz_dataOut_payload_0_4345;
  reg        [7:0]    _zz_dataOut_payload_0_4346;
  reg        [7:0]    _zz_dataOut_payload_0_4347;
  reg        [7:0]    _zz_dataOut_payload_0_4348;
  reg        [7:0]    _zz_dataOut_payload_0_4349;
  reg        [7:0]    _zz_dataOut_payload_0_4350;
  reg        [7:0]    _zz_dataOut_payload_0_4351;
  wire                _zz_dataOut_payload_0_4352;
  wire       [7:0]    _zz_dataOut_payload_0_4353;
  wire       [7:0]    _zz_dataOut_payload_0_4354;
  wire                _zz_dataOut_payload_0_4355;
  wire       [7:0]    _zz_dataOut_payload_0_4356;
  wire       [7:0]    _zz_dataOut_payload_0_4357;
  wire                _zz_dataOut_payload_0_4358;
  wire       [7:0]    _zz_dataOut_payload_0_4359;
  wire       [7:0]    _zz_dataOut_payload_0_4360;
  wire                _zz_dataOut_payload_0_4361;
  wire       [7:0]    _zz_dataOut_payload_0_4362;
  wire       [7:0]    _zz_dataOut_payload_0_4363;
  wire                _zz_dataOut_payload_0_4364;
  wire       [7:0]    _zz_dataOut_payload_0_4365;
  wire       [7:0]    _zz_dataOut_payload_0_4366;
  wire                _zz_dataOut_payload_0_4367;
  wire       [7:0]    _zz_dataOut_payload_0_4368;
  wire       [7:0]    _zz_dataOut_payload_0_4369;
  wire                _zz_dataOut_payload_0_4370;
  wire       [7:0]    _zz_dataOut_payload_0_4371;
  wire       [7:0]    _zz_dataOut_payload_0_4372;
  wire                _zz_dataOut_payload_0_4373;
  wire       [7:0]    _zz_dataOut_payload_0_4374;
  wire       [7:0]    _zz_dataOut_payload_0_4375;
  wire                _zz_dataOut_payload_0_4376;
  wire       [7:0]    _zz_dataOut_payload_0_4377;
  wire       [7:0]    _zz_dataOut_payload_0_4378;
  wire                _zz_dataOut_payload_0_4379;
  wire       [7:0]    _zz_dataOut_payload_0_4380;
  wire       [7:0]    _zz_dataOut_payload_0_4381;
  wire                _zz_dataOut_payload_0_4382;
  wire       [7:0]    _zz_dataOut_payload_0_4383;
  wire       [7:0]    _zz_dataOut_payload_0_4384;
  wire                _zz_dataOut_payload_0_4385;
  wire       [7:0]    _zz_dataOut_payload_0_4386;
  wire       [7:0]    _zz_dataOut_payload_0_4387;
  wire                _zz_dataOut_payload_0_4388;
  wire       [7:0]    _zz_dataOut_payload_0_4389;
  wire       [7:0]    _zz_dataOut_payload_0_4390;
  wire                _zz_dataOut_payload_0_4391;
  wire       [7:0]    _zz_dataOut_payload_0_4392;
  wire       [7:0]    _zz_dataOut_payload_0_4393;
  wire                _zz_dataOut_payload_0_4394;
  wire                _zz_dataOut_payload_0_4395;
  reg        [7:0]    _zz_dataOut_payload_0_4396;
  reg        [7:0]    _zz_dataOut_payload_0_4397;
  reg        [7:0]    _zz_dataOut_payload_0_4398;
  reg        [7:0]    _zz_dataOut_payload_0_4399;
  wire                _zz_dataOut_payload_0_4400;
  wire       [7:0]    _zz_dataOut_payload_0_4401;
  wire       [7:0]    _zz_dataOut_payload_0_4402;
  wire                _zz_dataOut_payload_0_4403;
  wire       [7:0]    _zz_dataOut_payload_0_4404;
  wire       [7:0]    _zz_dataOut_payload_0_4405;
  wire                _zz_dataOut_payload_0_4406;
  wire                _zz_dataOut_payload_0_4407;
  reg        [7:0]    _zz_dataOut_payload_0_4408;
  reg        [7:0]    _zz_dataOut_payload_0_4409;
  reg        [7:0]    _zz_dataOut_payload_0_4410;
  reg        [7:0]    _zz_dataOut_payload_0_4411;
  reg        [7:0]    _zz_dataOut_payload_0_4412;
  reg        [7:0]    _zz_dataOut_payload_0_4413;
  reg        [7:0]    _zz_dataOut_payload_0_4414;
  reg        [7:0]    _zz_dataOut_payload_0_4415;
  reg        [7:0]    _zz_dataOut_payload_0_4416;
  reg        [7:0]    _zz_dataOut_payload_0_4417;
  reg        [7:0]    _zz_dataOut_payload_0_4418;
  reg        [7:0]    _zz_dataOut_payload_0_4419;
  wire                _zz_dataOut_payload_0_4420;
  wire       [7:0]    _zz_dataOut_payload_0_4421;
  wire       [7:0]    _zz_dataOut_payload_0_4422;
  wire                _zz_dataOut_payload_0_4423;
  wire       [7:0]    _zz_dataOut_payload_0_4424;
  wire       [7:0]    _zz_dataOut_payload_0_4425;
  wire                _zz_dataOut_payload_0_4426;
  wire       [7:0]    _zz_dataOut_payload_0_4427;
  wire       [7:0]    _zz_dataOut_payload_0_4428;
  wire                _zz_dataOut_payload_0_4429;
  wire       [7:0]    _zz_dataOut_payload_0_4430;
  wire       [7:0]    _zz_dataOut_payload_0_4431;
  wire                _zz_dataOut_payload_0_4432;
  wire       [7:0]    _zz_dataOut_payload_0_4433;
  wire       [7:0]    _zz_dataOut_payload_0_4434;
  wire                _zz_dataOut_payload_0_4435;
  wire       [7:0]    _zz_dataOut_payload_0_4436;
  wire       [7:0]    _zz_dataOut_payload_0_4437;
  wire                _zz_dataOut_payload_0_4438;
  wire                _zz_dataOut_payload_0_4439;
  reg        [7:0]    _zz_dataOut_payload_0_4440;
  reg        [7:0]    _zz_dataOut_payload_0_4441;
  reg        [7:0]    _zz_dataOut_payload_0_4442;
  reg        [7:0]    _zz_dataOut_payload_0_4443;
  wire                _zz_dataOut_payload_0_4444;
  wire       [7:0]    _zz_dataOut_payload_0_4445;
  wire       [7:0]    _zz_dataOut_payload_0_4446;
  wire                _zz_dataOut_payload_0_4447;
  wire       [7:0]    _zz_dataOut_payload_0_4448;
  wire       [7:0]    _zz_dataOut_payload_0_4449;
  wire                _zz_dataOut_payload_0_4450;
  wire                _zz_dataOut_payload_0_4451;
  reg        [7:0]    _zz_dataOut_payload_0_4452;
  reg        [7:0]    _zz_dataOut_payload_0_4453;
  reg        [7:0]    _zz_dataOut_payload_0_4454;
  reg        [7:0]    _zz_dataOut_payload_0_4455;
  reg        [7:0]    _zz_dataOut_payload_0_4456;
  reg        [7:0]    _zz_dataOut_payload_0_4457;
  reg        [7:0]    _zz_dataOut_payload_0_4458;
  reg        [7:0]    _zz_dataOut_payload_0_4459;
  reg        [7:0]    _zz_dataOut_payload_0_4460;
  reg        [7:0]    _zz_dataOut_payload_0_4461;
  reg        [7:0]    _zz_dataOut_payload_0_4462;
  reg        [7:0]    _zz_dataOut_payload_0_4463;
  reg        [7:0]    _zz_dataOut_payload_0_4464;
  reg        [7:0]    _zz_dataOut_payload_0_4465;
  reg        [7:0]    _zz_dataOut_payload_0_4466;
  reg        [7:0]    _zz_dataOut_payload_0_4467;
  reg        [7:0]    _zz_dataOut_payload_0_4468;
  reg        [7:0]    _zz_dataOut_payload_0_4469;
  reg        [7:0]    _zz_dataOut_payload_0_4470;
  reg        [7:0]    _zz_dataOut_payload_0_4471;
  reg        [7:0]    _zz_dataOut_payload_0_4472;
  reg        [7:0]    _zz_dataOut_payload_0_4473;
  reg        [7:0]    _zz_dataOut_payload_0_4474;
  reg        [7:0]    _zz_dataOut_payload_0_4475;
  reg        [7:0]    _zz_dataOut_payload_0_4476;
  reg        [7:0]    _zz_dataOut_payload_0_4477;
  reg        [7:0]    _zz_dataOut_payload_0_4478;
  reg        [7:0]    _zz_dataOut_payload_0_4479;
  wire                _zz_dataOut_payload_0_4480;
  wire       [7:0]    _zz_dataOut_payload_0_4481;
  wire       [7:0]    _zz_dataOut_payload_0_4482;
  wire                _zz_dataOut_payload_0_4483;
  wire       [7:0]    _zz_dataOut_payload_0_4484;
  wire       [7:0]    _zz_dataOut_payload_0_4485;
  wire                _zz_dataOut_payload_0_4486;
  wire       [7:0]    _zz_dataOut_payload_0_4487;
  wire       [7:0]    _zz_dataOut_payload_0_4488;
  wire                _zz_dataOut_payload_0_4489;
  wire       [7:0]    _zz_dataOut_payload_0_4490;
  wire       [7:0]    _zz_dataOut_payload_0_4491;
  wire                _zz_dataOut_payload_0_4492;
  wire       [7:0]    _zz_dataOut_payload_0_4493;
  wire       [7:0]    _zz_dataOut_payload_0_4494;
  wire                _zz_dataOut_payload_0_4495;
  wire       [7:0]    _zz_dataOut_payload_0_4496;
  wire       [7:0]    _zz_dataOut_payload_0_4497;
  wire                _zz_dataOut_payload_0_4498;
  wire       [7:0]    _zz_dataOut_payload_0_4499;
  wire       [7:0]    _zz_dataOut_payload_0_4500;
  wire                _zz_dataOut_payload_0_4501;
  wire       [7:0]    _zz_dataOut_payload_0_4502;
  wire       [7:0]    _zz_dataOut_payload_0_4503;
  wire                _zz_dataOut_payload_0_4504;
  wire       [7:0]    _zz_dataOut_payload_0_4505;
  wire       [7:0]    _zz_dataOut_payload_0_4506;
  wire                _zz_dataOut_payload_0_4507;
  wire       [7:0]    _zz_dataOut_payload_0_4508;
  wire       [7:0]    _zz_dataOut_payload_0_4509;
  wire                _zz_dataOut_payload_0_4510;
  wire       [7:0]    _zz_dataOut_payload_0_4511;
  wire       [7:0]    _zz_dataOut_payload_0_4512;
  wire                _zz_dataOut_payload_0_4513;
  wire       [7:0]    _zz_dataOut_payload_0_4514;
  wire       [7:0]    _zz_dataOut_payload_0_4515;
  wire                _zz_dataOut_payload_0_4516;
  wire       [7:0]    _zz_dataOut_payload_0_4517;
  wire       [7:0]    _zz_dataOut_payload_0_4518;
  wire                _zz_dataOut_payload_0_4519;
  wire       [7:0]    _zz_dataOut_payload_0_4520;
  wire       [7:0]    _zz_dataOut_payload_0_4521;
  wire                _zz_dataOut_payload_0_4522;
  wire                _zz_dataOut_payload_0_4523;
  reg        [7:0]    _zz_dataOut_payload_0_4524;
  reg        [7:0]    _zz_dataOut_payload_0_4525;
  reg        [7:0]    _zz_dataOut_payload_0_4526;
  reg        [7:0]    _zz_dataOut_payload_0_4527;
  wire                _zz_dataOut_payload_0_4528;
  wire       [7:0]    _zz_dataOut_payload_0_4529;
  wire       [7:0]    _zz_dataOut_payload_0_4530;
  wire                _zz_dataOut_payload_0_4531;
  wire       [7:0]    _zz_dataOut_payload_0_4532;
  wire       [7:0]    _zz_dataOut_payload_0_4533;
  wire                _zz_dataOut_payload_0_4534;
  wire                _zz_dataOut_payload_0_4535;
  reg        [7:0]    _zz_dataOut_payload_0_4536;
  reg        [7:0]    _zz_dataOut_payload_0_4537;
  reg        [7:0]    _zz_dataOut_payload_0_4538;
  reg        [7:0]    _zz_dataOut_payload_0_4539;
  reg        [7:0]    _zz_dataOut_payload_0_4540;
  reg        [7:0]    _zz_dataOut_payload_0_4541;
  reg        [7:0]    _zz_dataOut_payload_0_4542;
  reg        [7:0]    _zz_dataOut_payload_0_4543;
  reg        [7:0]    _zz_dataOut_payload_0_4544;
  reg        [7:0]    _zz_dataOut_payload_0_4545;
  reg        [7:0]    _zz_dataOut_payload_0_4546;
  reg        [7:0]    _zz_dataOut_payload_0_4547;
  wire                _zz_dataOut_payload_0_4548;
  wire       [7:0]    _zz_dataOut_payload_0_4549;
  wire       [7:0]    _zz_dataOut_payload_0_4550;
  wire                _zz_dataOut_payload_0_4551;
  wire       [7:0]    _zz_dataOut_payload_0_4552;
  wire       [7:0]    _zz_dataOut_payload_0_4553;
  wire                _zz_dataOut_payload_0_4554;
  wire       [7:0]    _zz_dataOut_payload_0_4555;
  wire       [7:0]    _zz_dataOut_payload_0_4556;
  wire                _zz_dataOut_payload_0_4557;
  wire       [7:0]    _zz_dataOut_payload_0_4558;
  wire       [7:0]    _zz_dataOut_payload_0_4559;
  wire                _zz_dataOut_payload_0_4560;
  wire       [7:0]    _zz_dataOut_payload_0_4561;
  wire       [7:0]    _zz_dataOut_payload_0_4562;
  wire                _zz_dataOut_payload_0_4563;
  wire       [7:0]    _zz_dataOut_payload_0_4564;
  wire       [7:0]    _zz_dataOut_payload_0_4565;
  wire                _zz_dataOut_payload_0_4566;
  wire                _zz_dataOut_payload_0_4567;
  reg        [7:0]    _zz_dataOut_payload_0_4568;
  reg        [7:0]    _zz_dataOut_payload_0_4569;
  reg        [7:0]    _zz_dataOut_payload_0_4570;
  reg        [7:0]    _zz_dataOut_payload_0_4571;
  wire                _zz_dataOut_payload_0_4572;
  wire       [7:0]    _zz_dataOut_payload_0_4573;
  wire       [7:0]    _zz_dataOut_payload_0_4574;
  wire                _zz_dataOut_payload_0_4575;
  wire       [7:0]    _zz_dataOut_payload_0_4576;
  wire       [7:0]    _zz_dataOut_payload_0_4577;
  wire                _zz_dataOut_payload_0_4578;
  wire                _zz_dataOut_payload_0_4579;
  reg        [7:0]    _zz_dataOut_payload_0_4580;
  reg        [7:0]    _zz_dataOut_payload_0_4581;
  reg        [7:0]    _zz_dataOut_payload_0_4582;
  reg        [7:0]    _zz_dataOut_payload_0_4583;
  reg        [7:0]    _zz_dataOut_payload_0_4584;
  reg        [7:0]    _zz_dataOut_payload_0_4585;
  reg        [7:0]    _zz_dataOut_payload_0_4586;
  reg        [7:0]    _zz_dataOut_payload_0_4587;
  reg        [7:0]    _zz_dataOut_payload_0_4588;
  reg        [7:0]    _zz_dataOut_payload_0_4589;
  reg        [7:0]    _zz_dataOut_payload_0_4590;
  reg        [7:0]    _zz_dataOut_payload_0_4591;
  reg        [7:0]    _zz_dataOut_payload_0_4592;
  reg        [7:0]    _zz_dataOut_payload_0_4593;
  reg        [7:0]    _zz_dataOut_payload_0_4594;
  reg        [7:0]    _zz_dataOut_payload_0_4595;
  reg        [7:0]    _zz_dataOut_payload_0_4596;
  reg        [7:0]    _zz_dataOut_payload_0_4597;
  reg        [7:0]    _zz_dataOut_payload_0_4598;
  reg        [7:0]    _zz_dataOut_payload_0_4599;
  reg        [7:0]    _zz_dataOut_payload_0_4600;
  reg        [7:0]    _zz_dataOut_payload_0_4601;
  reg        [7:0]    _zz_dataOut_payload_0_4602;
  reg        [7:0]    _zz_dataOut_payload_0_4603;
  reg        [7:0]    _zz_dataOut_payload_0_4604;
  reg        [7:0]    _zz_dataOut_payload_0_4605;
  reg        [7:0]    _zz_dataOut_payload_0_4606;
  reg        [7:0]    _zz_dataOut_payload_0_4607;
  wire                _zz_dataOut_payload_0_4608;
  wire       [7:0]    _zz_dataOut_payload_0_4609;
  wire       [7:0]    _zz_dataOut_payload_0_4610;
  wire                _zz_dataOut_payload_0_4611;
  wire       [7:0]    _zz_dataOut_payload_0_4612;
  wire       [7:0]    _zz_dataOut_payload_0_4613;
  wire                _zz_dataOut_payload_0_4614;
  wire       [7:0]    _zz_dataOut_payload_0_4615;
  wire       [7:0]    _zz_dataOut_payload_0_4616;
  wire                _zz_dataOut_payload_0_4617;
  wire       [7:0]    _zz_dataOut_payload_0_4618;
  wire       [7:0]    _zz_dataOut_payload_0_4619;
  wire                _zz_dataOut_payload_0_4620;
  wire       [7:0]    _zz_dataOut_payload_0_4621;
  wire       [7:0]    _zz_dataOut_payload_0_4622;
  wire                _zz_dataOut_payload_0_4623;
  wire       [7:0]    _zz_dataOut_payload_0_4624;
  wire       [7:0]    _zz_dataOut_payload_0_4625;
  wire                _zz_dataOut_payload_0_4626;
  wire       [7:0]    _zz_dataOut_payload_0_4627;
  wire       [7:0]    _zz_dataOut_payload_0_4628;
  wire                _zz_dataOut_payload_0_4629;
  wire       [7:0]    _zz_dataOut_payload_0_4630;
  wire       [7:0]    _zz_dataOut_payload_0_4631;
  wire                _zz_dataOut_payload_0_4632;
  wire       [7:0]    _zz_dataOut_payload_0_4633;
  wire       [7:0]    _zz_dataOut_payload_0_4634;
  wire                _zz_dataOut_payload_0_4635;
  wire       [7:0]    _zz_dataOut_payload_0_4636;
  wire       [7:0]    _zz_dataOut_payload_0_4637;
  wire                _zz_dataOut_payload_0_4638;
  wire       [7:0]    _zz_dataOut_payload_0_4639;
  wire       [7:0]    _zz_dataOut_payload_0_4640;
  wire                _zz_dataOut_payload_0_4641;
  wire       [7:0]    _zz_dataOut_payload_0_4642;
  wire       [7:0]    _zz_dataOut_payload_0_4643;
  wire                _zz_dataOut_payload_0_4644;
  wire       [7:0]    _zz_dataOut_payload_0_4645;
  wire       [7:0]    _zz_dataOut_payload_0_4646;
  wire                _zz_dataOut_payload_0_4647;
  wire       [7:0]    _zz_dataOut_payload_0_4648;
  wire       [7:0]    _zz_dataOut_payload_0_4649;
  wire                _zz_dataOut_payload_0_4650;
  wire                _zz_dataOut_payload_0_4651;
  reg        [7:0]    _zz_dataOut_payload_0_4652;
  reg        [7:0]    _zz_dataOut_payload_0_4653;
  reg        [7:0]    _zz_dataOut_payload_0_4654;
  reg        [7:0]    _zz_dataOut_payload_0_4655;
  wire                _zz_dataOut_payload_0_4656;
  wire       [7:0]    _zz_dataOut_payload_0_4657;
  wire       [7:0]    _zz_dataOut_payload_0_4658;
  wire                _zz_dataOut_payload_0_4659;
  wire       [7:0]    _zz_dataOut_payload_0_4660;
  wire       [7:0]    _zz_dataOut_payload_0_4661;
  wire                _zz_dataOut_payload_0_4662;
  wire                _zz_dataOut_payload_0_4663;
  reg        [7:0]    _zz_dataOut_payload_0_4664;
  reg        [7:0]    _zz_dataOut_payload_0_4665;
  reg        [7:0]    _zz_dataOut_payload_0_4666;
  reg        [7:0]    _zz_dataOut_payload_0_4667;
  reg        [7:0]    _zz_dataOut_payload_0_4668;
  reg        [7:0]    _zz_dataOut_payload_0_4669;
  reg        [7:0]    _zz_dataOut_payload_0_4670;
  reg        [7:0]    _zz_dataOut_payload_0_4671;
  reg        [7:0]    _zz_dataOut_payload_0_4672;
  reg        [7:0]    _zz_dataOut_payload_0_4673;
  reg        [7:0]    _zz_dataOut_payload_0_4674;
  reg        [7:0]    _zz_dataOut_payload_0_4675;
  wire                _zz_dataOut_payload_0_4676;
  wire       [7:0]    _zz_dataOut_payload_0_4677;
  wire       [7:0]    _zz_dataOut_payload_0_4678;
  wire                _zz_dataOut_payload_0_4679;
  wire       [7:0]    _zz_dataOut_payload_0_4680;
  wire       [7:0]    _zz_dataOut_payload_0_4681;
  wire                _zz_dataOut_payload_0_4682;
  wire       [7:0]    _zz_dataOut_payload_0_4683;
  wire       [7:0]    _zz_dataOut_payload_0_4684;
  wire                _zz_dataOut_payload_0_4685;
  wire       [7:0]    _zz_dataOut_payload_0_4686;
  wire       [7:0]    _zz_dataOut_payload_0_4687;
  wire                _zz_dataOut_payload_0_4688;
  wire       [7:0]    _zz_dataOut_payload_0_4689;
  wire       [7:0]    _zz_dataOut_payload_0_4690;
  wire                _zz_dataOut_payload_0_4691;
  wire       [7:0]    _zz_dataOut_payload_0_4692;
  wire       [7:0]    _zz_dataOut_payload_0_4693;
  wire                _zz_dataOut_payload_0_4694;
  wire                _zz_dataOut_payload_0_4695;
  reg        [7:0]    _zz_dataOut_payload_0_4696;
  reg        [7:0]    _zz_dataOut_payload_0_4697;
  reg        [7:0]    _zz_dataOut_payload_0_4698;
  reg        [7:0]    _zz_dataOut_payload_0_4699;
  wire                _zz_dataOut_payload_0_4700;
  wire       [7:0]    _zz_dataOut_payload_0_4701;
  wire       [7:0]    _zz_dataOut_payload_0_4702;
  wire                _zz_dataOut_payload_0_4703;
  wire       [7:0]    _zz_dataOut_payload_0_4704;
  wire       [7:0]    _zz_dataOut_payload_0_4705;
  wire                _zz_dataOut_payload_0_4706;
  wire                _zz_dataOut_payload_0_4707;
  reg        [7:0]    _zz_dataOut_payload_0_4708;
  reg        [7:0]    _zz_dataOut_payload_0_4709;
  reg        [7:0]    _zz_dataOut_payload_0_4710;
  reg        [7:0]    _zz_dataOut_payload_0_4711;
  reg        [7:0]    _zz_dataOut_payload_0_4712;
  reg        [7:0]    _zz_dataOut_payload_0_4713;
  reg        [7:0]    _zz_dataOut_payload_0_4714;
  reg        [7:0]    _zz_dataOut_payload_0_4715;
  reg        [7:0]    _zz_dataOut_payload_0_4716;
  reg        [7:0]    _zz_dataOut_payload_0_4717;
  reg        [7:0]    _zz_dataOut_payload_0_4718;
  reg        [7:0]    _zz_dataOut_payload_0_4719;
  reg        [7:0]    _zz_dataOut_payload_0_4720;
  reg        [7:0]    _zz_dataOut_payload_0_4721;
  reg        [7:0]    _zz_dataOut_payload_0_4722;
  reg        [7:0]    _zz_dataOut_payload_0_4723;
  reg        [7:0]    _zz_dataOut_payload_0_4724;
  reg        [7:0]    _zz_dataOut_payload_0_4725;
  reg        [7:0]    _zz_dataOut_payload_0_4726;
  reg        [7:0]    _zz_dataOut_payload_0_4727;
  reg        [7:0]    _zz_dataOut_payload_0_4728;
  reg        [7:0]    _zz_dataOut_payload_0_4729;
  reg        [7:0]    _zz_dataOut_payload_0_4730;
  reg        [7:0]    _zz_dataOut_payload_0_4731;
  reg        [7:0]    _zz_dataOut_payload_0_4732;
  reg        [7:0]    _zz_dataOut_payload_0_4733;
  reg        [7:0]    _zz_dataOut_payload_0_4734;
  reg        [7:0]    _zz_dataOut_payload_0_4735;
  wire                _zz_dataOut_payload_0_4736;
  wire       [7:0]    _zz_dataOut_payload_0_4737;
  wire       [7:0]    _zz_dataOut_payload_0_4738;
  wire                _zz_dataOut_payload_0_4739;
  wire       [7:0]    _zz_dataOut_payload_0_4740;
  wire       [7:0]    _zz_dataOut_payload_0_4741;
  wire                _zz_dataOut_payload_0_4742;
  wire       [7:0]    _zz_dataOut_payload_0_4743;
  wire       [7:0]    _zz_dataOut_payload_0_4744;
  wire                _zz_dataOut_payload_0_4745;
  wire       [7:0]    _zz_dataOut_payload_0_4746;
  wire       [7:0]    _zz_dataOut_payload_0_4747;
  wire                _zz_dataOut_payload_0_4748;
  wire       [7:0]    _zz_dataOut_payload_0_4749;
  wire       [7:0]    _zz_dataOut_payload_0_4750;
  wire                _zz_dataOut_payload_0_4751;
  wire       [7:0]    _zz_dataOut_payload_0_4752;
  wire       [7:0]    _zz_dataOut_payload_0_4753;
  wire                _zz_dataOut_payload_0_4754;
  wire       [7:0]    _zz_dataOut_payload_0_4755;
  wire       [7:0]    _zz_dataOut_payload_0_4756;
  wire                _zz_dataOut_payload_0_4757;
  wire       [7:0]    _zz_dataOut_payload_0_4758;
  wire       [7:0]    _zz_dataOut_payload_0_4759;
  wire                _zz_dataOut_payload_0_4760;
  wire       [7:0]    _zz_dataOut_payload_0_4761;
  wire       [7:0]    _zz_dataOut_payload_0_4762;
  wire                _zz_dataOut_payload_0_4763;
  wire       [7:0]    _zz_dataOut_payload_0_4764;
  wire       [7:0]    _zz_dataOut_payload_0_4765;
  wire                _zz_dataOut_payload_0_4766;
  wire       [7:0]    _zz_dataOut_payload_0_4767;
  wire       [7:0]    _zz_dataOut_payload_0_4768;
  wire                _zz_dataOut_payload_0_4769;
  wire       [7:0]    _zz_dataOut_payload_0_4770;
  wire       [7:0]    _zz_dataOut_payload_0_4771;
  wire                _zz_dataOut_payload_0_4772;
  wire       [7:0]    _zz_dataOut_payload_0_4773;
  wire       [7:0]    _zz_dataOut_payload_0_4774;
  wire                _zz_dataOut_payload_0_4775;
  wire       [7:0]    _zz_dataOut_payload_0_4776;
  wire       [7:0]    _zz_dataOut_payload_0_4777;
  wire                _zz_dataOut_payload_0_4778;
  wire                _zz_dataOut_payload_0_4779;
  reg        [7:0]    _zz_dataOut_payload_0_4780;
  reg        [7:0]    _zz_dataOut_payload_0_4781;
  reg        [7:0]    _zz_dataOut_payload_0_4782;
  reg        [7:0]    _zz_dataOut_payload_0_4783;
  wire                _zz_dataOut_payload_0_4784;
  wire       [7:0]    _zz_dataOut_payload_0_4785;
  wire       [7:0]    _zz_dataOut_payload_0_4786;
  wire                _zz_dataOut_payload_0_4787;
  wire       [7:0]    _zz_dataOut_payload_0_4788;
  wire       [7:0]    _zz_dataOut_payload_0_4789;
  wire                _zz_dataOut_payload_0_4790;
  wire                _zz_dataOut_payload_0_4791;
  reg        [7:0]    _zz_dataOut_payload_0_4792;
  reg        [7:0]    _zz_dataOut_payload_0_4793;
  reg        [7:0]    _zz_dataOut_payload_0_4794;
  reg        [7:0]    _zz_dataOut_payload_0_4795;
  reg        [7:0]    _zz_dataOut_payload_0_4796;
  reg        [7:0]    _zz_dataOut_payload_0_4797;
  reg        [7:0]    _zz_dataOut_payload_0_4798;
  reg        [7:0]    _zz_dataOut_payload_0_4799;
  reg        [7:0]    _zz_dataOut_payload_0_4800;
  reg        [7:0]    _zz_dataOut_payload_0_4801;
  reg        [7:0]    _zz_dataOut_payload_0_4802;
  reg        [7:0]    _zz_dataOut_payload_0_4803;
  wire                _zz_dataOut_payload_0_4804;
  wire       [7:0]    _zz_dataOut_payload_0_4805;
  wire       [7:0]    _zz_dataOut_payload_0_4806;
  wire                _zz_dataOut_payload_0_4807;
  wire       [7:0]    _zz_dataOut_payload_0_4808;
  wire       [7:0]    _zz_dataOut_payload_0_4809;
  wire                _zz_dataOut_payload_0_4810;
  wire       [7:0]    _zz_dataOut_payload_0_4811;
  wire       [7:0]    _zz_dataOut_payload_0_4812;
  wire                _zz_dataOut_payload_0_4813;
  wire       [7:0]    _zz_dataOut_payload_0_4814;
  wire       [7:0]    _zz_dataOut_payload_0_4815;
  wire                _zz_dataOut_payload_0_4816;
  wire       [7:0]    _zz_dataOut_payload_0_4817;
  wire       [7:0]    _zz_dataOut_payload_0_4818;
  wire                _zz_dataOut_payload_0_4819;
  wire       [7:0]    _zz_dataOut_payload_0_4820;
  wire       [7:0]    _zz_dataOut_payload_0_4821;
  wire                _zz_dataOut_payload_0_4822;
  wire                _zz_dataOut_payload_0_4823;
  reg        [7:0]    _zz_dataOut_payload_0_4824;
  reg        [7:0]    _zz_dataOut_payload_0_4825;
  reg        [7:0]    _zz_dataOut_payload_0_4826;
  reg        [7:0]    _zz_dataOut_payload_0_4827;
  wire                _zz_dataOut_payload_0_4828;
  wire       [7:0]    _zz_dataOut_payload_0_4829;
  wire       [7:0]    _zz_dataOut_payload_0_4830;
  wire                _zz_dataOut_payload_0_4831;
  wire       [7:0]    _zz_dataOut_payload_0_4832;
  wire       [7:0]    _zz_dataOut_payload_0_4833;
  wire                _zz_dataOut_payload_0_4834;
  wire                _zz_dataOut_payload_0_4835;
  reg        [7:0]    _zz_dataOut_payload_0_4836;
  reg        [7:0]    _zz_dataOut_payload_0_4837;
  reg        [7:0]    _zz_dataOut_payload_0_4838;
  reg        [7:0]    _zz_dataOut_payload_0_4839;
  reg        [7:0]    _zz_dataOut_payload_0_4840;
  reg        [7:0]    _zz_dataOut_payload_0_4841;
  reg        [7:0]    _zz_dataOut_payload_0_4842;
  reg        [7:0]    _zz_dataOut_payload_0_4843;
  reg        [7:0]    _zz_dataOut_payload_0_4844;
  reg        [7:0]    _zz_dataOut_payload_0_4845;
  reg        [7:0]    _zz_dataOut_payload_0_4846;
  reg        [7:0]    _zz_dataOut_payload_0_4847;
  reg        [7:0]    _zz_dataOut_payload_0_4848;
  reg        [7:0]    _zz_dataOut_payload_0_4849;
  reg        [7:0]    _zz_dataOut_payload_0_4850;
  reg        [7:0]    _zz_dataOut_payload_0_4851;
  reg        [7:0]    _zz_dataOut_payload_0_4852;
  reg        [7:0]    _zz_dataOut_payload_0_4853;
  reg        [7:0]    _zz_dataOut_payload_0_4854;
  reg        [7:0]    _zz_dataOut_payload_0_4855;
  reg        [7:0]    _zz_dataOut_payload_0_4856;
  reg        [7:0]    _zz_dataOut_payload_0_4857;
  reg        [7:0]    _zz_dataOut_payload_0_4858;
  reg        [7:0]    _zz_dataOut_payload_0_4859;
  reg        [7:0]    _zz_dataOut_payload_0_4860;
  reg        [7:0]    _zz_dataOut_payload_0_4861;
  reg        [7:0]    _zz_dataOut_payload_0_4862;
  reg        [7:0]    _zz_dataOut_payload_0_4863;
  wire                _zz_dataOut_payload_0_4864;
  wire       [7:0]    _zz_dataOut_payload_0_4865;
  wire       [7:0]    _zz_dataOut_payload_0_4866;
  wire                _zz_dataOut_payload_0_4867;
  wire       [7:0]    _zz_dataOut_payload_0_4868;
  wire       [7:0]    _zz_dataOut_payload_0_4869;
  wire                _zz_dataOut_payload_0_4870;
  wire       [7:0]    _zz_dataOut_payload_0_4871;
  wire       [7:0]    _zz_dataOut_payload_0_4872;
  wire                _zz_dataOut_payload_0_4873;
  wire       [7:0]    _zz_dataOut_payload_0_4874;
  wire       [7:0]    _zz_dataOut_payload_0_4875;
  wire                _zz_dataOut_payload_0_4876;
  wire       [7:0]    _zz_dataOut_payload_0_4877;
  wire       [7:0]    _zz_dataOut_payload_0_4878;
  wire                _zz_dataOut_payload_0_4879;
  wire       [7:0]    _zz_dataOut_payload_0_4880;
  wire       [7:0]    _zz_dataOut_payload_0_4881;
  wire                _zz_dataOut_payload_0_4882;
  wire       [7:0]    _zz_dataOut_payload_0_4883;
  wire       [7:0]    _zz_dataOut_payload_0_4884;
  wire                _zz_dataOut_payload_0_4885;
  wire       [7:0]    _zz_dataOut_payload_0_4886;
  wire       [7:0]    _zz_dataOut_payload_0_4887;
  wire                _zz_dataOut_payload_0_4888;
  wire       [7:0]    _zz_dataOut_payload_0_4889;
  wire       [7:0]    _zz_dataOut_payload_0_4890;
  wire                _zz_dataOut_payload_0_4891;
  wire       [7:0]    _zz_dataOut_payload_0_4892;
  wire       [7:0]    _zz_dataOut_payload_0_4893;
  wire                _zz_dataOut_payload_0_4894;
  wire       [7:0]    _zz_dataOut_payload_0_4895;
  wire       [7:0]    _zz_dataOut_payload_0_4896;
  wire                _zz_dataOut_payload_0_4897;
  wire       [7:0]    _zz_dataOut_payload_0_4898;
  wire       [7:0]    _zz_dataOut_payload_0_4899;
  wire                _zz_dataOut_payload_0_4900;
  wire       [7:0]    _zz_dataOut_payload_0_4901;
  wire       [7:0]    _zz_dataOut_payload_0_4902;
  wire                _zz_dataOut_payload_0_4903;
  wire       [7:0]    _zz_dataOut_payload_0_4904;
  wire       [7:0]    _zz_dataOut_payload_0_4905;
  wire                _zz_dataOut_payload_0_4906;
  wire                _zz_dataOut_payload_0_4907;
  reg        [7:0]    _zz_dataOut_payload_0_4908;
  reg        [7:0]    _zz_dataOut_payload_0_4909;
  reg        [7:0]    _zz_dataOut_payload_0_4910;
  reg        [7:0]    _zz_dataOut_payload_0_4911;
  wire                _zz_dataOut_payload_0_4912;
  wire       [7:0]    _zz_dataOut_payload_0_4913;
  wire       [7:0]    _zz_dataOut_payload_0_4914;
  wire                _zz_dataOut_payload_0_4915;
  wire       [7:0]    _zz_dataOut_payload_0_4916;
  wire       [7:0]    _zz_dataOut_payload_0_4917;
  wire                _zz_dataOut_payload_0_4918;
  wire                _zz_dataOut_payload_0_4919;
  reg        [7:0]    _zz_dataOut_payload_0_4920;
  reg        [7:0]    _zz_dataOut_payload_0_4921;
  reg        [7:0]    _zz_dataOut_payload_0_4922;
  reg        [7:0]    _zz_dataOut_payload_0_4923;
  reg        [7:0]    _zz_dataOut_payload_0_4924;
  reg        [7:0]    _zz_dataOut_payload_0_4925;
  reg        [7:0]    _zz_dataOut_payload_0_4926;
  reg        [7:0]    _zz_dataOut_payload_0_4927;
  reg        [7:0]    _zz_dataOut_payload_0_4928;
  reg        [7:0]    _zz_dataOut_payload_0_4929;
  reg        [7:0]    _zz_dataOut_payload_0_4930;
  reg        [7:0]    _zz_dataOut_payload_0_4931;
  wire                _zz_dataOut_payload_0_4932;
  wire       [7:0]    _zz_dataOut_payload_0_4933;
  wire       [7:0]    _zz_dataOut_payload_0_4934;
  wire                _zz_dataOut_payload_0_4935;
  wire       [7:0]    _zz_dataOut_payload_0_4936;
  wire       [7:0]    _zz_dataOut_payload_0_4937;
  wire                _zz_dataOut_payload_0_4938;
  wire       [7:0]    _zz_dataOut_payload_0_4939;
  wire       [7:0]    _zz_dataOut_payload_0_4940;
  wire                _zz_dataOut_payload_0_4941;
  wire       [7:0]    _zz_dataOut_payload_0_4942;
  wire       [7:0]    _zz_dataOut_payload_0_4943;
  wire                _zz_dataOut_payload_0_4944;
  wire       [7:0]    _zz_dataOut_payload_0_4945;
  wire       [7:0]    _zz_dataOut_payload_0_4946;
  wire                _zz_dataOut_payload_0_4947;
  wire       [7:0]    _zz_dataOut_payload_0_4948;
  wire       [7:0]    _zz_dataOut_payload_0_4949;
  wire                _zz_dataOut_payload_0_4950;
  wire                _zz_dataOut_payload_0_4951;
  reg        [7:0]    _zz_dataOut_payload_0_4952;
  reg        [7:0]    _zz_dataOut_payload_0_4953;
  reg        [7:0]    _zz_dataOut_payload_0_4954;
  reg        [7:0]    _zz_dataOut_payload_0_4955;
  wire                _zz_dataOut_payload_0_4956;
  wire       [7:0]    _zz_dataOut_payload_0_4957;
  wire       [7:0]    _zz_dataOut_payload_0_4958;
  wire                _zz_dataOut_payload_0_4959;
  wire       [7:0]    _zz_dataOut_payload_0_4960;
  wire       [7:0]    _zz_dataOut_payload_0_4961;
  wire                _zz_dataOut_payload_0_4962;
  wire                _zz_dataOut_payload_0_4963;
  reg        [7:0]    _zz_dataOut_payload_0_4964;
  reg        [7:0]    _zz_dataOut_payload_0_4965;
  reg        [7:0]    _zz_dataOut_payload_0_4966;
  reg        [7:0]    _zz_dataOut_payload_0_4967;
  reg        [7:0]    _zz_dataOut_payload_0_4968;
  reg        [7:0]    _zz_dataOut_payload_0_4969;
  reg        [7:0]    _zz_dataOut_payload_0_4970;
  reg        [7:0]    _zz_dataOut_payload_0_4971;
  reg        [7:0]    _zz_dataOut_payload_0_4972;
  reg        [7:0]    _zz_dataOut_payload_0_4973;
  reg        [7:0]    _zz_dataOut_payload_0_4974;
  reg        [7:0]    _zz_dataOut_payload_0_4975;
  reg        [7:0]    _zz_dataOut_payload_0_4976;
  reg        [7:0]    _zz_dataOut_payload_0_4977;
  reg        [7:0]    _zz_dataOut_payload_0_4978;
  reg        [7:0]    _zz_dataOut_payload_0_4979;
  reg        [7:0]    _zz_dataOut_payload_0_4980;
  reg        [7:0]    _zz_dataOut_payload_0_4981;
  reg        [7:0]    _zz_dataOut_payload_0_4982;
  reg        [7:0]    _zz_dataOut_payload_0_4983;
  reg        [7:0]    _zz_dataOut_payload_0_4984;
  reg        [7:0]    _zz_dataOut_payload_0_4985;
  reg        [7:0]    _zz_dataOut_payload_0_4986;
  reg        [7:0]    _zz_dataOut_payload_0_4987;
  reg        [7:0]    _zz_dataOut_payload_0_4988;
  reg        [7:0]    _zz_dataOut_payload_0_4989;
  reg        [7:0]    _zz_dataOut_payload_0_4990;
  reg        [7:0]    _zz_dataOut_payload_0_4991;
  wire                _zz_dataOut_payload_0_4992;
  wire       [7:0]    _zz_dataOut_payload_0_4993;
  wire       [7:0]    _zz_dataOut_payload_0_4994;
  wire                _zz_dataOut_payload_0_4995;
  wire       [7:0]    _zz_dataOut_payload_0_4996;
  wire       [7:0]    _zz_dataOut_payload_0_4997;
  wire                _zz_dataOut_payload_0_4998;
  wire       [7:0]    _zz_dataOut_payload_0_4999;
  wire       [7:0]    _zz_dataOut_payload_0_5000;
  wire                _zz_dataOut_payload_0_5001;
  wire       [7:0]    _zz_dataOut_payload_0_5002;
  wire       [7:0]    _zz_dataOut_payload_0_5003;
  wire                _zz_dataOut_payload_0_5004;
  wire       [7:0]    _zz_dataOut_payload_0_5005;
  wire       [7:0]    _zz_dataOut_payload_0_5006;
  wire                _zz_dataOut_payload_0_5007;
  wire       [7:0]    _zz_dataOut_payload_0_5008;
  wire       [7:0]    _zz_dataOut_payload_0_5009;
  wire                _zz_dataOut_payload_0_5010;
  wire       [7:0]    _zz_dataOut_payload_0_5011;
  wire       [7:0]    _zz_dataOut_payload_0_5012;
  wire                _zz_dataOut_payload_0_5013;
  wire       [7:0]    _zz_dataOut_payload_0_5014;
  wire       [7:0]    _zz_dataOut_payload_0_5015;
  wire                _zz_dataOut_payload_0_5016;
  wire       [7:0]    _zz_dataOut_payload_0_5017;
  wire       [7:0]    _zz_dataOut_payload_0_5018;
  wire                _zz_dataOut_payload_0_5019;
  wire       [7:0]    _zz_dataOut_payload_0_5020;
  wire       [7:0]    _zz_dataOut_payload_0_5021;
  wire                _zz_dataOut_payload_0_5022;
  wire       [7:0]    _zz_dataOut_payload_0_5023;
  wire       [7:0]    _zz_dataOut_payload_0_5024;
  wire                _zz_dataOut_payload_0_5025;
  wire       [7:0]    _zz_dataOut_payload_0_5026;
  wire       [7:0]    _zz_dataOut_payload_0_5027;
  wire                _zz_dataOut_payload_0_5028;
  wire       [7:0]    _zz_dataOut_payload_0_5029;
  wire       [7:0]    _zz_dataOut_payload_0_5030;
  wire                _zz_dataOut_payload_0_5031;
  wire       [7:0]    _zz_dataOut_payload_0_5032;
  wire       [7:0]    _zz_dataOut_payload_0_5033;
  wire                _zz_dataOut_payload_0_5034;
  wire                _zz_dataOut_payload_0_5035;
  reg        [7:0]    _zz_dataOut_payload_0_5036;
  reg        [7:0]    _zz_dataOut_payload_0_5037;
  reg        [7:0]    _zz_dataOut_payload_0_5038;
  reg        [7:0]    _zz_dataOut_payload_0_5039;
  wire                _zz_dataOut_payload_0_5040;
  wire       [7:0]    _zz_dataOut_payload_0_5041;
  wire       [7:0]    _zz_dataOut_payload_0_5042;
  wire                _zz_dataOut_payload_0_5043;
  wire       [7:0]    _zz_dataOut_payload_0_5044;
  wire       [7:0]    _zz_dataOut_payload_0_5045;
  wire                _zz_dataOut_payload_0_5046;
  wire                _zz_dataOut_payload_0_5047;
  reg        [7:0]    _zz_dataOut_payload_0_5048;
  reg        [7:0]    _zz_dataOut_payload_0_5049;
  reg        [7:0]    _zz_dataOut_payload_0_5050;
  reg        [7:0]    _zz_dataOut_payload_0_5051;
  reg        [7:0]    _zz_dataOut_payload_0_5052;
  reg        [7:0]    _zz_dataOut_payload_0_5053;
  reg        [7:0]    _zz_dataOut_payload_0_5054;
  reg        [7:0]    _zz_dataOut_payload_0_5055;
  reg        [7:0]    _zz_dataOut_payload_0_5056;
  reg        [7:0]    _zz_dataOut_payload_0_5057;
  reg        [7:0]    _zz_dataOut_payload_0_5058;
  reg        [7:0]    _zz_dataOut_payload_0_5059;
  wire                _zz_dataOut_payload_0_5060;
  wire       [7:0]    _zz_dataOut_payload_0_5061;
  wire       [7:0]    _zz_dataOut_payload_0_5062;
  wire                _zz_dataOut_payload_0_5063;
  wire       [7:0]    _zz_dataOut_payload_0_5064;
  wire       [7:0]    _zz_dataOut_payload_0_5065;
  wire                _zz_dataOut_payload_0_5066;
  wire       [7:0]    _zz_dataOut_payload_0_5067;
  wire       [7:0]    _zz_dataOut_payload_0_5068;
  wire                _zz_dataOut_payload_0_5069;
  wire       [7:0]    _zz_dataOut_payload_0_5070;
  wire       [7:0]    _zz_dataOut_payload_0_5071;
  wire                _zz_dataOut_payload_0_5072;
  wire       [7:0]    _zz_dataOut_payload_0_5073;
  wire       [7:0]    _zz_dataOut_payload_0_5074;
  wire                _zz_dataOut_payload_0_5075;
  wire       [7:0]    _zz_dataOut_payload_0_5076;
  wire       [7:0]    _zz_dataOut_payload_0_5077;
  wire                _zz_dataOut_payload_0_5078;
  wire                _zz_dataOut_payload_0_5079;
  reg        [7:0]    _zz_dataOut_payload_0_5080;
  reg        [7:0]    _zz_dataOut_payload_0_5081;
  reg        [7:0]    _zz_dataOut_payload_0_5082;
  reg        [7:0]    _zz_dataOut_payload_0_5083;
  wire                _zz_dataOut_payload_0_5084;
  wire       [7:0]    _zz_dataOut_payload_0_5085;
  wire       [7:0]    _zz_dataOut_payload_0_5086;
  wire                _zz_dataOut_payload_0_5087;
  wire       [7:0]    _zz_dataOut_payload_0_5088;
  wire       [7:0]    _zz_dataOut_payload_0_5089;
  wire                _zz_dataOut_payload_0_5090;
  wire                _zz_dataOut_payload_0_5091;
  reg        [7:0]    _zz_dataOut_payload_0_5092;
  reg        [7:0]    _zz_dataOut_payload_0_5093;
  reg        [7:0]    _zz_dataOut_payload_0_5094;
  reg        [7:0]    _zz_dataOut_payload_0_5095;
  reg        [7:0]    _zz_dataOut_payload_0_5096;
  reg        [7:0]    _zz_dataOut_payload_0_5097;
  reg        [7:0]    _zz_dataOut_payload_0_5098;
  reg        [7:0]    _zz_dataOut_payload_0_5099;
  reg        [7:0]    _zz_dataOut_payload_0_5100;
  reg        [7:0]    _zz_dataOut_payload_0_5101;
  reg        [7:0]    _zz_dataOut_payload_0_5102;
  reg        [7:0]    _zz_dataOut_payload_0_5103;
  reg        [7:0]    _zz_dataOut_payload_0_5104;
  reg        [7:0]    _zz_dataOut_payload_0_5105;
  reg        [7:0]    _zz_dataOut_payload_0_5106;
  reg        [7:0]    _zz_dataOut_payload_0_5107;
  reg        [7:0]    _zz_dataOut_payload_0_5108;
  reg        [7:0]    _zz_dataOut_payload_0_5109;
  reg        [7:0]    _zz_dataOut_payload_0_5110;
  reg        [7:0]    _zz_dataOut_payload_0_5111;
  reg        [7:0]    _zz_dataOut_payload_0_5112;
  reg        [7:0]    _zz_dataOut_payload_0_5113;
  reg        [7:0]    _zz_dataOut_payload_0_5114;
  reg        [7:0]    _zz_dataOut_payload_0_5115;
  reg        [7:0]    _zz_dataOut_payload_0_5116;
  reg        [7:0]    _zz_dataOut_payload_0_5117;
  reg        [7:0]    _zz_dataOut_payload_0_5118;
  reg        [7:0]    _zz_dataOut_payload_0_5119;
  reg        [7:0]    _zz_dataOut_payload_0_5120;
  reg        [7:0]    _zz_dataOut_payload_0_5121;
  reg        [7:0]    _zz_dataOut_payload_0_5122;
  reg        [7:0]    _zz_dataOut_payload_0_5123;
  reg        [7:0]    _zz_dataOut_payload_0_5124;
  reg        [7:0]    _zz_dataOut_payload_0_5125;
  reg        [7:0]    _zz_dataOut_payload_0_5126;
  reg        [7:0]    _zz_dataOut_payload_0_5127;
  reg        [7:0]    _zz_dataOut_payload_0_5128;
  reg        [7:0]    _zz_dataOut_payload_0_5129;
  reg        [7:0]    _zz_dataOut_payload_0_5130;
  reg        [7:0]    _zz_dataOut_payload_0_5131;
  reg        [7:0]    _zz_dataOut_payload_0_5132;
  reg        [7:0]    _zz_dataOut_payload_0_5133;
  reg        [7:0]    _zz_dataOut_payload_0_5134;
  reg        [7:0]    _zz_dataOut_payload_0_5135;
  reg        [7:0]    _zz_dataOut_payload_0_5136;
  reg        [7:0]    _zz_dataOut_payload_0_5137;
  reg        [7:0]    _zz_dataOut_payload_0_5138;
  reg        [7:0]    _zz_dataOut_payload_0_5139;
  reg        [7:0]    _zz_dataOut_payload_0_5140;
  reg        [7:0]    _zz_dataOut_payload_0_5141;
  reg        [7:0]    _zz_dataOut_payload_0_5142;
  reg        [7:0]    _zz_dataOut_payload_0_5143;
  reg        [7:0]    _zz_dataOut_payload_0_5144;
  reg        [7:0]    _zz_dataOut_payload_0_5145;
  reg        [7:0]    _zz_dataOut_payload_0_5146;
  reg        [7:0]    _zz_dataOut_payload_0_5147;
  reg        [7:0]    _zz_dataOut_payload_0_5148;
  reg        [7:0]    _zz_dataOut_payload_0_5149;
  reg        [7:0]    _zz_dataOut_payload_0_5150;
  reg        [7:0]    _zz_dataOut_payload_0_5151;
  reg        [7:0]    _zz_dataOut_payload_0_5152;
  reg        [7:0]    _zz_dataOut_payload_0_5153;
  reg        [7:0]    _zz_dataOut_payload_0_5154;
  reg        [7:0]    _zz_dataOut_payload_0_5155;
  reg        [7:0]    _zz_dataOut_payload_0_5156;
  reg        [7:0]    _zz_dataOut_payload_0_5157;
  reg        [7:0]    _zz_dataOut_payload_0_5158;
  reg        [7:0]    _zz_dataOut_payload_0_5159;
  reg        [7:0]    _zz_dataOut_payload_0_5160;
  reg        [7:0]    _zz_dataOut_payload_0_5161;
  reg        [7:0]    _zz_dataOut_payload_0_5162;
  reg        [7:0]    _zz_dataOut_payload_0_5163;
  reg        [7:0]    _zz_dataOut_payload_0_5164;
  reg        [7:0]    _zz_dataOut_payload_0_5165;
  reg        [7:0]    _zz_dataOut_payload_0_5166;
  reg        [7:0]    _zz_dataOut_payload_0_5167;
  reg        [7:0]    _zz_dataOut_payload_0_5168;
  reg        [7:0]    _zz_dataOut_payload_0_5169;
  reg        [7:0]    _zz_dataOut_payload_0_5170;
  reg        [7:0]    _zz_dataOut_payload_0_5171;
  reg        [7:0]    _zz_dataOut_payload_0_5172;
  reg        [7:0]    _zz_dataOut_payload_0_5173;
  reg        [7:0]    _zz_dataOut_payload_0_5174;
  reg        [7:0]    _zz_dataOut_payload_0_5175;
  reg        [7:0]    _zz_dataOut_payload_0_5176;
  reg        [7:0]    _zz_dataOut_payload_0_5177;
  reg        [7:0]    _zz_dataOut_payload_0_5178;
  reg        [7:0]    _zz_dataOut_payload_0_5179;
  reg        [7:0]    _zz_dataOut_payload_0_5180;
  reg        [7:0]    _zz_dataOut_payload_0_5181;
  reg        [7:0]    _zz_dataOut_payload_0_5182;
  reg        [7:0]    _zz_dataOut_payload_0_5183;
  reg        [7:0]    _zz_dataOut_payload_0_5184;
  reg        [7:0]    _zz_dataOut_payload_0_5185;
  reg        [7:0]    _zz_dataOut_payload_0_5186;
  reg        [7:0]    _zz_dataOut_payload_0_5187;
  reg        [7:0]    _zz_dataOut_payload_0_5188;
  reg        [7:0]    _zz_dataOut_payload_0_5189;
  reg        [7:0]    _zz_dataOut_payload_0_5190;
  reg        [7:0]    _zz_dataOut_payload_0_5191;
  reg        [7:0]    _zz_dataOut_payload_0_5192;
  reg        [7:0]    _zz_dataOut_payload_0_5193;
  reg        [7:0]    _zz_dataOut_payload_0_5194;
  reg        [7:0]    _zz_dataOut_payload_0_5195;
  reg        [7:0]    _zz_dataOut_payload_0_5196;
  reg        [7:0]    _zz_dataOut_payload_0_5197;
  reg        [7:0]    _zz_dataOut_payload_0_5198;
  reg        [7:0]    _zz_dataOut_payload_0_5199;
  reg        [7:0]    _zz_dataOut_payload_0_5200;
  reg        [7:0]    _zz_dataOut_payload_0_5201;
  reg        [7:0]    _zz_dataOut_payload_0_5202;
  reg        [7:0]    _zz_dataOut_payload_0_5203;
  reg        [7:0]    _zz_dataOut_payload_0_5204;
  reg        [7:0]    _zz_dataOut_payload_0_5205;
  reg        [7:0]    _zz_dataOut_payload_0_5206;
  reg        [7:0]    _zz_dataOut_payload_0_5207;
  reg        [7:0]    _zz_dataOut_payload_0_5208;
  reg        [7:0]    _zz_dataOut_payload_0_5209;
  reg        [7:0]    _zz_dataOut_payload_0_5210;
  reg        [7:0]    _zz_dataOut_payload_0_5211;
  reg        [7:0]    _zz_dataOut_payload_0_5212;
  reg        [7:0]    _zz_dataOut_payload_0_5213;
  reg        [7:0]    _zz_dataOut_payload_0_5214;
  reg        [7:0]    _zz_dataOut_payload_0_5215;
  reg        [7:0]    _zz_dataOut_payload_0_5216;
  reg        [7:0]    _zz_dataOut_payload_0_5217;
  reg        [7:0]    _zz_dataOut_payload_0_5218;
  reg        [7:0]    _zz_dataOut_payload_0_5219;
  reg        [7:0]    _zz_dataOut_payload_0_5220;
  reg        [7:0]    _zz_dataOut_payload_0_5221;
  reg        [7:0]    _zz_dataOut_payload_0_5222;
  reg        [7:0]    _zz_dataOut_payload_0_5223;
  reg        [7:0]    _zz_dataOut_payload_0_5224;
  reg        [7:0]    _zz_dataOut_payload_0_5225;
  reg        [7:0]    _zz_dataOut_payload_0_5226;
  reg        [7:0]    _zz_dataOut_payload_0_5227;
  reg        [7:0]    _zz_dataOut_payload_0_5228;
  reg        [7:0]    _zz_dataOut_payload_0_5229;
  reg        [7:0]    _zz_dataOut_payload_0_5230;
  reg        [7:0]    _zz_dataOut_payload_0_5231;
  reg        [7:0]    _zz_dataOut_payload_0_5232;
  reg        [7:0]    _zz_dataOut_payload_0_5233;
  reg        [7:0]    _zz_dataOut_payload_0_5234;
  reg        [7:0]    _zz_dataOut_payload_0_5235;
  reg        [7:0]    _zz_dataOut_payload_0_5236;
  reg        [7:0]    _zz_dataOut_payload_0_5237;
  reg        [7:0]    _zz_dataOut_payload_0_5238;
  reg        [7:0]    _zz_dataOut_payload_0_5239;
  reg        [7:0]    _zz_dataOut_payload_0_5240;
  reg        [7:0]    _zz_dataOut_payload_0_5241;
  reg        [7:0]    _zz_dataOut_payload_0_5242;
  reg        [7:0]    _zz_dataOut_payload_0_5243;
  reg        [7:0]    _zz_dataOut_payload_0_5244;
  reg        [7:0]    _zz_dataOut_payload_0_5245;
  reg        [7:0]    _zz_dataOut_payload_0_5246;
  reg        [7:0]    _zz_dataOut_payload_0_5247;
  reg        [7:0]    _zz_dataOut_payload_0_5248;
  reg        [7:0]    _zz_dataOut_payload_0_5249;
  reg        [7:0]    _zz_dataOut_payload_0_5250;
  reg        [7:0]    _zz_dataOut_payload_0_5251;
  reg        [7:0]    _zz_dataOut_payload_0_5252;
  reg        [7:0]    _zz_dataOut_payload_0_5253;
  reg        [7:0]    _zz_dataOut_payload_0_5254;
  reg        [7:0]    _zz_dataOut_payload_0_5255;
  reg        [7:0]    _zz_dataOut_payload_0_5256;
  reg        [7:0]    _zz_dataOut_payload_0_5257;
  reg        [7:0]    _zz_dataOut_payload_0_5258;
  reg        [7:0]    _zz_dataOut_payload_0_5259;
  reg        [7:0]    _zz_dataOut_payload_0_5260;
  reg        [7:0]    _zz_dataOut_payload_0_5261;
  reg        [7:0]    _zz_dataOut_payload_0_5262;
  reg        [7:0]    _zz_dataOut_payload_0_5263;
  reg        [7:0]    _zz_dataOut_payload_0_5264;
  reg        [7:0]    _zz_dataOut_payload_0_5265;
  reg        [7:0]    _zz_dataOut_payload_0_5266;
  reg        [7:0]    _zz_dataOut_payload_0_5267;
  reg        [7:0]    _zz_dataOut_payload_0_5268;
  reg        [7:0]    _zz_dataOut_payload_0_5269;
  reg        [7:0]    _zz_dataOut_payload_0_5270;
  reg        [7:0]    _zz_dataOut_payload_0_5271;
  reg        [7:0]    _zz_dataOut_payload_0_5272;
  reg        [7:0]    _zz_dataOut_payload_0_5273;
  reg        [7:0]    _zz_dataOut_payload_0_5274;
  reg        [7:0]    _zz_dataOut_payload_0_5275;
  reg        [7:0]    _zz_dataOut_payload_0_5276;
  reg        [7:0]    _zz_dataOut_payload_0_5277;
  reg        [7:0]    _zz_dataOut_payload_0_5278;
  reg        [7:0]    _zz_dataOut_payload_0_5279;
  reg        [7:0]    _zz_dataOut_payload_0_5280;
  reg        [7:0]    _zz_dataOut_payload_0_5281;
  reg        [7:0]    _zz_dataOut_payload_0_5282;
  reg        [7:0]    _zz_dataOut_payload_0_5283;
  reg        [7:0]    _zz_dataOut_payload_0_5284;
  reg        [7:0]    _zz_dataOut_payload_0_5285;
  reg        [7:0]    _zz_dataOut_payload_0_5286;
  reg        [7:0]    _zz_dataOut_payload_0_5287;
  reg        [7:0]    _zz_dataOut_payload_0_5288;
  reg        [7:0]    _zz_dataOut_payload_0_5289;
  reg        [7:0]    _zz_dataOut_payload_0_5290;
  reg        [7:0]    _zz_dataOut_payload_0_5291;
  reg        [7:0]    _zz_dataOut_payload_0_5292;
  reg        [7:0]    _zz_dataOut_payload_0_5293;
  reg        [7:0]    _zz_dataOut_payload_0_5294;
  reg        [7:0]    _zz_dataOut_payload_0_5295;
  reg        [7:0]    _zz_dataOut_payload_0_5296;
  reg        [7:0]    _zz_dataOut_payload_0_5297;
  reg        [7:0]    _zz_dataOut_payload_0_5298;
  reg        [7:0]    _zz_dataOut_payload_0_5299;
  reg        [7:0]    _zz_dataOut_payload_0_5300;
  reg        [7:0]    _zz_dataOut_payload_0_5301;
  reg        [7:0]    _zz_dataOut_payload_0_5302;
  reg        [7:0]    _zz_dataOut_payload_0_5303;
  reg        [7:0]    _zz_dataOut_payload_0_5304;
  reg        [7:0]    _zz_dataOut_payload_0_5305;
  reg        [7:0]    _zz_dataOut_payload_0_5306;
  reg        [7:0]    _zz_dataOut_payload_0_5307;
  reg        [7:0]    _zz_dataOut_payload_0_5308;
  reg        [7:0]    _zz_dataOut_payload_0_5309;
  reg        [7:0]    _zz_dataOut_payload_0_5310;
  reg        [7:0]    _zz_dataOut_payload_0_5311;
  reg        [7:0]    _zz_dataOut_payload_0_5312;
  reg        [7:0]    _zz_dataOut_payload_0_5313;
  reg        [7:0]    _zz_dataOut_payload_0_5314;
  reg        [7:0]    _zz_dataOut_payload_0_5315;
  reg        [7:0]    _zz_dataOut_payload_0_5316;
  reg        [7:0]    _zz_dataOut_payload_0_5317;
  reg        [7:0]    _zz_dataOut_payload_0_5318;
  reg        [7:0]    _zz_dataOut_payload_0_5319;
  reg        [7:0]    _zz_dataOut_payload_0_5320;
  reg        [7:0]    _zz_dataOut_payload_0_5321;
  reg        [7:0]    _zz_dataOut_payload_0_5322;
  reg        [7:0]    _zz_dataOut_payload_0_5323;
  reg        [7:0]    _zz_dataOut_payload_0_5324;
  reg        [7:0]    _zz_dataOut_payload_0_5325;
  reg        [7:0]    _zz_dataOut_payload_0_5326;
  reg        [7:0]    _zz_dataOut_payload_0_5327;
  reg        [7:0]    _zz_dataOut_payload_0_5328;
  reg        [7:0]    _zz_dataOut_payload_0_5329;
  reg        [7:0]    _zz_dataOut_payload_0_5330;
  reg        [7:0]    _zz_dataOut_payload_0_5331;
  reg        [7:0]    _zz_dataOut_payload_0_5332;
  reg        [7:0]    _zz_dataOut_payload_0_5333;
  reg        [7:0]    _zz_dataOut_payload_0_5334;
  reg        [7:0]    _zz_dataOut_payload_0_5335;
  reg        [7:0]    _zz_dataOut_payload_0_5336;
  reg        [7:0]    _zz_dataOut_payload_0_5337;
  reg        [7:0]    _zz_dataOut_payload_0_5338;
  reg        [7:0]    _zz_dataOut_payload_0_5339;
  reg        [7:0]    _zz_dataOut_payload_0_5340;
  reg        [7:0]    _zz_dataOut_payload_0_5341;
  reg        [7:0]    _zz_dataOut_payload_0_5342;
  reg        [7:0]    _zz_dataOut_payload_0_5343;
  reg        [7:0]    _zz_dataOut_payload_0_5344;
  reg        [7:0]    _zz_dataOut_payload_0_5345;
  reg        [7:0]    _zz_dataOut_payload_0_5346;
  reg        [7:0]    _zz_dataOut_payload_0_5347;
  reg        [7:0]    _zz_dataOut_payload_0_5348;
  reg        [7:0]    _zz_dataOut_payload_0_5349;
  reg        [7:0]    _zz_dataOut_payload_0_5350;
  reg        [7:0]    _zz_dataOut_payload_0_5351;
  reg        [7:0]    _zz_dataOut_payload_0_5352;
  reg        [7:0]    _zz_dataOut_payload_0_5353;
  reg        [7:0]    _zz_dataOut_payload_0_5354;
  reg        [7:0]    _zz_dataOut_payload_0_5355;
  reg        [7:0]    _zz_dataOut_payload_0_5356;
  reg        [7:0]    _zz_dataOut_payload_0_5357;
  reg        [7:0]    _zz_dataOut_payload_0_5358;
  reg        [7:0]    _zz_dataOut_payload_0_5359;
  reg        [7:0]    _zz_dataOut_payload_0_5360;
  reg        [7:0]    _zz_dataOut_payload_0_5361;
  reg        [7:0]    _zz_dataOut_payload_0_5362;
  reg        [7:0]    _zz_dataOut_payload_0_5363;
  reg        [7:0]    _zz_dataOut_payload_0_5364;
  reg        [7:0]    _zz_dataOut_payload_0_5365;
  reg        [7:0]    _zz_dataOut_payload_0_5366;
  reg        [7:0]    _zz_dataOut_payload_0_5367;
  reg        [7:0]    _zz_dataOut_payload_0_5368;
  reg        [7:0]    _zz_dataOut_payload_0_5369;
  reg        [7:0]    _zz_dataOut_payload_0_5370;
  reg        [7:0]    _zz_dataOut_payload_0_5371;
  reg        [7:0]    _zz_dataOut_payload_0_5372;
  reg        [7:0]    _zz_dataOut_payload_0_5373;
  reg        [7:0]    _zz_dataOut_payload_0_5374;
  reg        [7:0]    _zz_dataOut_payload_0_5375;
  wire                _zz_dataOut_payload_0_5376;
  wire       [7:0]    _zz_dataOut_payload_0_5377;
  wire       [7:0]    _zz_dataOut_payload_0_5378;
  wire                _zz_dataOut_payload_0_5379;
  wire       [7:0]    _zz_dataOut_payload_0_5380;
  wire       [7:0]    _zz_dataOut_payload_0_5381;
  wire                _zz_dataOut_payload_0_5382;
  wire       [7:0]    _zz_dataOut_payload_0_5383;
  wire       [7:0]    _zz_dataOut_payload_0_5384;
  wire                _zz_dataOut_payload_0_5385;
  wire       [7:0]    _zz_dataOut_payload_0_5386;
  wire       [7:0]    _zz_dataOut_payload_0_5387;
  wire                _zz_dataOut_payload_0_5388;
  wire       [7:0]    _zz_dataOut_payload_0_5389;
  wire       [7:0]    _zz_dataOut_payload_0_5390;
  wire                _zz_dataOut_payload_0_5391;
  wire       [7:0]    _zz_dataOut_payload_0_5392;
  wire       [7:0]    _zz_dataOut_payload_0_5393;
  wire                _zz_dataOut_payload_0_5394;
  wire       [7:0]    _zz_dataOut_payload_0_5395;
  wire       [7:0]    _zz_dataOut_payload_0_5396;
  wire                _zz_dataOut_payload_0_5397;
  wire       [7:0]    _zz_dataOut_payload_0_5398;
  wire       [7:0]    _zz_dataOut_payload_0_5399;
  wire                _zz_dataOut_payload_0_5400;
  wire       [7:0]    _zz_dataOut_payload_0_5401;
  wire       [7:0]    _zz_dataOut_payload_0_5402;
  wire                _zz_dataOut_payload_0_5403;
  wire       [7:0]    _zz_dataOut_payload_0_5404;
  wire       [7:0]    _zz_dataOut_payload_0_5405;
  wire                _zz_dataOut_payload_0_5406;
  wire       [7:0]    _zz_dataOut_payload_0_5407;
  wire       [7:0]    _zz_dataOut_payload_0_5408;
  wire                _zz_dataOut_payload_0_5409;
  wire       [7:0]    _zz_dataOut_payload_0_5410;
  wire       [7:0]    _zz_dataOut_payload_0_5411;
  wire                _zz_dataOut_payload_0_5412;
  wire       [7:0]    _zz_dataOut_payload_0_5413;
  wire       [7:0]    _zz_dataOut_payload_0_5414;
  wire                _zz_dataOut_payload_0_5415;
  wire       [7:0]    _zz_dataOut_payload_0_5416;
  wire       [7:0]    _zz_dataOut_payload_0_5417;
  wire                _zz_dataOut_payload_0_5418;
  wire       [7:0]    _zz_dataOut_payload_0_5419;
  wire       [7:0]    _zz_dataOut_payload_0_5420;
  wire                _zz_dataOut_payload_0_5421;
  wire       [7:0]    _zz_dataOut_payload_0_5422;
  wire       [7:0]    _zz_dataOut_payload_0_5423;
  wire                _zz_dataOut_payload_0_5424;
  wire       [7:0]    _zz_dataOut_payload_0_5425;
  wire       [7:0]    _zz_dataOut_payload_0_5426;
  wire                _zz_dataOut_payload_0_5427;
  wire       [7:0]    _zz_dataOut_payload_0_5428;
  wire       [7:0]    _zz_dataOut_payload_0_5429;
  wire                _zz_dataOut_payload_0_5430;
  wire       [7:0]    _zz_dataOut_payload_0_5431;
  wire       [7:0]    _zz_dataOut_payload_0_5432;
  wire                _zz_dataOut_payload_0_5433;
  wire       [7:0]    _zz_dataOut_payload_0_5434;
  wire       [7:0]    _zz_dataOut_payload_0_5435;
  wire                _zz_dataOut_payload_0_5436;
  wire       [7:0]    _zz_dataOut_payload_0_5437;
  wire       [7:0]    _zz_dataOut_payload_0_5438;
  wire                _zz_dataOut_payload_0_5439;
  wire       [7:0]    _zz_dataOut_payload_0_5440;
  wire       [7:0]    _zz_dataOut_payload_0_5441;
  wire                _zz_dataOut_payload_0_5442;
  wire       [7:0]    _zz_dataOut_payload_0_5443;
  wire       [7:0]    _zz_dataOut_payload_0_5444;
  wire                _zz_dataOut_payload_0_5445;
  wire       [7:0]    _zz_dataOut_payload_0_5446;
  wire       [7:0]    _zz_dataOut_payload_0_5447;
  wire                _zz_dataOut_payload_0_5448;
  wire       [7:0]    _zz_dataOut_payload_0_5449;
  wire       [7:0]    _zz_dataOut_payload_0_5450;
  wire                _zz_dataOut_payload_0_5451;
  wire       [7:0]    _zz_dataOut_payload_0_5452;
  wire       [7:0]    _zz_dataOut_payload_0_5453;
  wire                _zz_dataOut_payload_0_5454;
  wire       [7:0]    _zz_dataOut_payload_0_5455;
  wire       [7:0]    _zz_dataOut_payload_0_5456;
  wire                _zz_dataOut_payload_0_5457;
  wire       [7:0]    _zz_dataOut_payload_0_5458;
  wire       [7:0]    _zz_dataOut_payload_0_5459;
  wire                _zz_dataOut_payload_0_5460;
  wire       [7:0]    _zz_dataOut_payload_0_5461;
  wire       [7:0]    _zz_dataOut_payload_0_5462;
  wire                _zz_dataOut_payload_0_5463;
  wire       [7:0]    _zz_dataOut_payload_0_5464;
  wire       [7:0]    _zz_dataOut_payload_0_5465;
  wire                _zz_dataOut_payload_0_5466;
  wire                _zz_dataOut_payload_0_5467;
  reg        [7:0]    _zz_dataOut_payload_0_5468;
  reg        [7:0]    _zz_dataOut_payload_0_5469;
  reg        [7:0]    _zz_dataOut_payload_0_5470;
  reg        [7:0]    _zz_dataOut_payload_0_5471;
  wire                _zz_dataOut_payload_0_5472;
  wire       [7:0]    _zz_dataOut_payload_0_5473;
  wire       [7:0]    _zz_dataOut_payload_0_5474;
  wire                _zz_dataOut_payload_0_5475;
  wire       [7:0]    _zz_dataOut_payload_0_5476;
  wire       [7:0]    _zz_dataOut_payload_0_5477;
  wire                _zz_dataOut_payload_0_5478;
  wire                _zz_dataOut_payload_0_5479;
  reg        [7:0]    _zz_dataOut_payload_0_5480;
  reg        [7:0]    _zz_dataOut_payload_0_5481;
  reg        [7:0]    _zz_dataOut_payload_0_5482;
  reg        [7:0]    _zz_dataOut_payload_0_5483;
  reg        [7:0]    _zz_dataOut_payload_0_5484;
  reg        [7:0]    _zz_dataOut_payload_0_5485;
  reg        [7:0]    _zz_dataOut_payload_0_5486;
  reg        [7:0]    _zz_dataOut_payload_0_5487;
  reg        [7:0]    _zz_dataOut_payload_0_5488;
  reg        [7:0]    _zz_dataOut_payload_0_5489;
  reg        [7:0]    _zz_dataOut_payload_0_5490;
  reg        [7:0]    _zz_dataOut_payload_0_5491;
  wire                _zz_dataOut_payload_0_5492;
  wire       [7:0]    _zz_dataOut_payload_0_5493;
  wire       [7:0]    _zz_dataOut_payload_0_5494;
  wire                _zz_dataOut_payload_0_5495;
  wire       [7:0]    _zz_dataOut_payload_0_5496;
  wire       [7:0]    _zz_dataOut_payload_0_5497;
  wire                _zz_dataOut_payload_0_5498;
  wire       [7:0]    _zz_dataOut_payload_0_5499;
  wire       [7:0]    _zz_dataOut_payload_0_5500;
  wire                _zz_dataOut_payload_0_5501;
  wire       [7:0]    _zz_dataOut_payload_0_5502;
  wire       [7:0]    _zz_dataOut_payload_0_5503;
  wire                _zz_dataOut_payload_0_5504;
  wire       [7:0]    _zz_dataOut_payload_0_5505;
  wire       [7:0]    _zz_dataOut_payload_0_5506;
  wire                _zz_dataOut_payload_0_5507;
  wire       [7:0]    _zz_dataOut_payload_0_5508;
  wire       [7:0]    _zz_dataOut_payload_0_5509;
  wire                _zz_dataOut_payload_0_5510;
  wire                _zz_dataOut_payload_0_5511;
  reg        [7:0]    _zz_dataOut_payload_0_5512;
  reg        [7:0]    _zz_dataOut_payload_0_5513;
  reg        [7:0]    _zz_dataOut_payload_0_5514;
  reg        [7:0]    _zz_dataOut_payload_0_5515;
  wire                _zz_dataOut_payload_0_5516;
  wire       [7:0]    _zz_dataOut_payload_0_5517;
  wire       [7:0]    _zz_dataOut_payload_0_5518;
  wire                _zz_dataOut_payload_0_5519;
  wire       [7:0]    _zz_dataOut_payload_0_5520;
  wire       [7:0]    _zz_dataOut_payload_0_5521;
  wire                _zz_dataOut_payload_0_5522;
  wire                _zz_dataOut_payload_0_5523;
  reg        [7:0]    _zz_dataOut_payload_0_5524;
  reg        [7:0]    _zz_dataOut_payload_0_5525;
  reg        [7:0]    _zz_dataOut_payload_0_5526;
  reg        [7:0]    _zz_dataOut_payload_0_5527;
  reg        [7:0]    _zz_dataOut_payload_0_5528;
  reg        [7:0]    _zz_dataOut_payload_0_5529;
  reg        [7:0]    _zz_dataOut_payload_0_5530;
  reg        [7:0]    _zz_dataOut_payload_0_5531;
  reg        [7:0]    _zz_dataOut_payload_0_5532;
  reg        [7:0]    _zz_dataOut_payload_0_5533;
  reg        [7:0]    _zz_dataOut_payload_0_5534;
  reg        [7:0]    _zz_dataOut_payload_0_5535;
  reg        [7:0]    _zz_dataOut_payload_0_5536;
  reg        [7:0]    _zz_dataOut_payload_0_5537;
  reg        [7:0]    _zz_dataOut_payload_0_5538;
  reg        [7:0]    _zz_dataOut_payload_0_5539;
  reg        [7:0]    _zz_dataOut_payload_0_5540;
  reg        [7:0]    _zz_dataOut_payload_0_5541;
  reg        [7:0]    _zz_dataOut_payload_0_5542;
  reg        [7:0]    _zz_dataOut_payload_0_5543;
  reg        [7:0]    _zz_dataOut_payload_0_5544;
  reg        [7:0]    _zz_dataOut_payload_0_5545;
  reg        [7:0]    _zz_dataOut_payload_0_5546;
  reg        [7:0]    _zz_dataOut_payload_0_5547;
  reg        [7:0]    _zz_dataOut_payload_0_5548;
  reg        [7:0]    _zz_dataOut_payload_0_5549;
  reg        [7:0]    _zz_dataOut_payload_0_5550;
  reg        [7:0]    _zz_dataOut_payload_0_5551;
  wire                _zz_dataOut_payload_0_5552;
  wire       [7:0]    _zz_dataOut_payload_0_5553;
  wire       [7:0]    _zz_dataOut_payload_0_5554;
  wire                _zz_dataOut_payload_0_5555;
  wire       [7:0]    _zz_dataOut_payload_0_5556;
  wire       [7:0]    _zz_dataOut_payload_0_5557;
  wire                _zz_dataOut_payload_0_5558;
  wire       [7:0]    _zz_dataOut_payload_0_5559;
  wire       [7:0]    _zz_dataOut_payload_0_5560;
  wire                _zz_dataOut_payload_0_5561;
  wire       [7:0]    _zz_dataOut_payload_0_5562;
  wire       [7:0]    _zz_dataOut_payload_0_5563;
  wire                _zz_dataOut_payload_0_5564;
  wire       [7:0]    _zz_dataOut_payload_0_5565;
  wire       [7:0]    _zz_dataOut_payload_0_5566;
  wire                _zz_dataOut_payload_0_5567;
  wire       [7:0]    _zz_dataOut_payload_0_5568;
  wire       [7:0]    _zz_dataOut_payload_0_5569;
  wire                _zz_dataOut_payload_0_5570;
  wire       [7:0]    _zz_dataOut_payload_0_5571;
  wire       [7:0]    _zz_dataOut_payload_0_5572;
  wire                _zz_dataOut_payload_0_5573;
  wire       [7:0]    _zz_dataOut_payload_0_5574;
  wire       [7:0]    _zz_dataOut_payload_0_5575;
  wire                _zz_dataOut_payload_0_5576;
  wire       [7:0]    _zz_dataOut_payload_0_5577;
  wire       [7:0]    _zz_dataOut_payload_0_5578;
  wire                _zz_dataOut_payload_0_5579;
  wire       [7:0]    _zz_dataOut_payload_0_5580;
  wire       [7:0]    _zz_dataOut_payload_0_5581;
  wire                _zz_dataOut_payload_0_5582;
  wire       [7:0]    _zz_dataOut_payload_0_5583;
  wire       [7:0]    _zz_dataOut_payload_0_5584;
  wire                _zz_dataOut_payload_0_5585;
  wire       [7:0]    _zz_dataOut_payload_0_5586;
  wire       [7:0]    _zz_dataOut_payload_0_5587;
  wire                _zz_dataOut_payload_0_5588;
  wire       [7:0]    _zz_dataOut_payload_0_5589;
  wire       [7:0]    _zz_dataOut_payload_0_5590;
  wire                _zz_dataOut_payload_0_5591;
  wire       [7:0]    _zz_dataOut_payload_0_5592;
  wire       [7:0]    _zz_dataOut_payload_0_5593;
  wire                _zz_dataOut_payload_0_5594;
  wire                _zz_dataOut_payload_0_5595;
  reg        [7:0]    _zz_dataOut_payload_0_5596;
  reg        [7:0]    _zz_dataOut_payload_0_5597;
  reg        [7:0]    _zz_dataOut_payload_0_5598;
  reg        [7:0]    _zz_dataOut_payload_0_5599;
  wire                _zz_dataOut_payload_0_5600;
  wire       [7:0]    _zz_dataOut_payload_0_5601;
  wire       [7:0]    _zz_dataOut_payload_0_5602;
  wire                _zz_dataOut_payload_0_5603;
  wire       [7:0]    _zz_dataOut_payload_0_5604;
  wire       [7:0]    _zz_dataOut_payload_0_5605;
  wire                _zz_dataOut_payload_0_5606;
  wire                _zz_dataOut_payload_0_5607;
  reg        [7:0]    _zz_dataOut_payload_0_5608;
  reg        [7:0]    _zz_dataOut_payload_0_5609;
  reg        [7:0]    _zz_dataOut_payload_0_5610;
  reg        [7:0]    _zz_dataOut_payload_0_5611;
  reg        [7:0]    _zz_dataOut_payload_0_5612;
  reg        [7:0]    _zz_dataOut_payload_0_5613;
  reg        [7:0]    _zz_dataOut_payload_0_5614;
  reg        [7:0]    _zz_dataOut_payload_0_5615;
  reg        [7:0]    _zz_dataOut_payload_0_5616;
  reg        [7:0]    _zz_dataOut_payload_0_5617;
  reg        [7:0]    _zz_dataOut_payload_0_5618;
  reg        [7:0]    _zz_dataOut_payload_0_5619;
  wire                _zz_dataOut_payload_0_5620;
  wire       [7:0]    _zz_dataOut_payload_0_5621;
  wire       [7:0]    _zz_dataOut_payload_0_5622;
  wire                _zz_dataOut_payload_0_5623;
  wire       [7:0]    _zz_dataOut_payload_0_5624;
  wire       [7:0]    _zz_dataOut_payload_0_5625;
  wire                _zz_dataOut_payload_0_5626;
  wire       [7:0]    _zz_dataOut_payload_0_5627;
  wire       [7:0]    _zz_dataOut_payload_0_5628;
  wire                _zz_dataOut_payload_0_5629;
  wire       [7:0]    _zz_dataOut_payload_0_5630;
  wire       [7:0]    _zz_dataOut_payload_0_5631;
  wire                _zz_dataOut_payload_0_5632;
  wire       [7:0]    _zz_dataOut_payload_0_5633;
  wire       [7:0]    _zz_dataOut_payload_0_5634;
  wire                _zz_dataOut_payload_0_5635;
  wire       [7:0]    _zz_dataOut_payload_0_5636;
  wire       [7:0]    _zz_dataOut_payload_0_5637;
  wire                _zz_dataOut_payload_0_5638;
  wire                _zz_dataOut_payload_0_5639;
  reg        [7:0]    _zz_dataOut_payload_0_5640;
  reg        [7:0]    _zz_dataOut_payload_0_5641;
  reg        [7:0]    _zz_dataOut_payload_0_5642;
  reg        [7:0]    _zz_dataOut_payload_0_5643;
  wire                _zz_dataOut_payload_0_5644;
  wire       [7:0]    _zz_dataOut_payload_0_5645;
  wire       [7:0]    _zz_dataOut_payload_0_5646;
  wire                _zz_dataOut_payload_0_5647;
  wire       [7:0]    _zz_dataOut_payload_0_5648;
  wire       [7:0]    _zz_dataOut_payload_0_5649;
  wire                _zz_dataOut_payload_0_5650;
  wire                _zz_dataOut_payload_0_5651;
  reg        [7:0]    _zz_dataOut_payload_0_5652;
  reg        [7:0]    _zz_dataOut_payload_0_5653;
  reg        [7:0]    _zz_dataOut_payload_0_5654;
  reg        [7:0]    _zz_dataOut_payload_0_5655;
  reg        [7:0]    _zz_dataOut_payload_0_5656;
  reg        [7:0]    _zz_dataOut_payload_0_5657;
  reg        [7:0]    _zz_dataOut_payload_0_5658;
  reg        [7:0]    _zz_dataOut_payload_0_5659;
  reg        [7:0]    _zz_dataOut_payload_0_5660;
  reg        [7:0]    _zz_dataOut_payload_0_5661;
  reg        [7:0]    _zz_dataOut_payload_0_5662;
  reg        [7:0]    _zz_dataOut_payload_0_5663;
  reg        [7:0]    _zz_dataOut_payload_0_5664;
  reg        [7:0]    _zz_dataOut_payload_0_5665;
  reg        [7:0]    _zz_dataOut_payload_0_5666;
  reg        [7:0]    _zz_dataOut_payload_0_5667;
  reg        [7:0]    _zz_dataOut_payload_0_5668;
  reg        [7:0]    _zz_dataOut_payload_0_5669;
  reg        [7:0]    _zz_dataOut_payload_0_5670;
  reg        [7:0]    _zz_dataOut_payload_0_5671;
  reg        [7:0]    _zz_dataOut_payload_0_5672;
  reg        [7:0]    _zz_dataOut_payload_0_5673;
  reg        [7:0]    _zz_dataOut_payload_0_5674;
  reg        [7:0]    _zz_dataOut_payload_0_5675;
  reg        [7:0]    _zz_dataOut_payload_0_5676;
  reg        [7:0]    _zz_dataOut_payload_0_5677;
  reg        [7:0]    _zz_dataOut_payload_0_5678;
  reg        [7:0]    _zz_dataOut_payload_0_5679;
  reg        [7:0]    _zz_dataOut_payload_0_5680;
  reg        [7:0]    _zz_dataOut_payload_0_5681;
  reg        [7:0]    _zz_dataOut_payload_0_5682;
  reg        [7:0]    _zz_dataOut_payload_0_5683;
  reg        [7:0]    _zz_dataOut_payload_0_5684;
  reg        [7:0]    _zz_dataOut_payload_0_5685;
  reg        [7:0]    _zz_dataOut_payload_0_5686;
  reg        [7:0]    _zz_dataOut_payload_0_5687;
  reg        [7:0]    _zz_dataOut_payload_0_5688;
  reg        [7:0]    _zz_dataOut_payload_0_5689;
  reg        [7:0]    _zz_dataOut_payload_0_5690;
  reg        [7:0]    _zz_dataOut_payload_0_5691;
  reg        [7:0]    _zz_dataOut_payload_0_5692;
  reg        [7:0]    _zz_dataOut_payload_0_5693;
  reg        [7:0]    _zz_dataOut_payload_0_5694;
  reg        [7:0]    _zz_dataOut_payload_0_5695;
  reg        [7:0]    _zz_dataOut_payload_0_5696;
  reg        [7:0]    _zz_dataOut_payload_0_5697;
  reg        [7:0]    _zz_dataOut_payload_0_5698;
  reg        [7:0]    _zz_dataOut_payload_0_5699;
  reg        [7:0]    _zz_dataOut_payload_0_5700;
  reg        [7:0]    _zz_dataOut_payload_0_5701;
  reg        [7:0]    _zz_dataOut_payload_0_5702;
  reg        [7:0]    _zz_dataOut_payload_0_5703;
  reg        [7:0]    _zz_dataOut_payload_0_5704;
  reg        [7:0]    _zz_dataOut_payload_0_5705;
  reg        [7:0]    _zz_dataOut_payload_0_5706;
  reg        [7:0]    _zz_dataOut_payload_0_5707;
  reg        [7:0]    _zz_dataOut_payload_0_5708;
  reg        [7:0]    _zz_dataOut_payload_0_5709;
  reg        [7:0]    _zz_dataOut_payload_0_5710;
  reg        [7:0]    _zz_dataOut_payload_0_5711;
  wire                _zz_dataOut_payload_0_5712;
  wire       [7:0]    _zz_dataOut_payload_0_5713;
  wire       [7:0]    _zz_dataOut_payload_0_5714;
  wire                _zz_dataOut_payload_0_5715;
  wire       [7:0]    _zz_dataOut_payload_0_5716;
  wire       [7:0]    _zz_dataOut_payload_0_5717;
  wire                _zz_dataOut_payload_0_5718;
  wire       [7:0]    _zz_dataOut_payload_0_5719;
  wire       [7:0]    _zz_dataOut_payload_0_5720;
  wire                _zz_dataOut_payload_0_5721;
  wire       [7:0]    _zz_dataOut_payload_0_5722;
  wire       [7:0]    _zz_dataOut_payload_0_5723;
  wire                _zz_dataOut_payload_0_5724;
  wire       [7:0]    _zz_dataOut_payload_0_5725;
  wire       [7:0]    _zz_dataOut_payload_0_5726;
  wire                _zz_dataOut_payload_0_5727;
  wire       [7:0]    _zz_dataOut_payload_0_5728;
  wire       [7:0]    _zz_dataOut_payload_0_5729;
  wire                _zz_dataOut_payload_0_5730;
  wire       [7:0]    _zz_dataOut_payload_0_5731;
  wire       [7:0]    _zz_dataOut_payload_0_5732;
  wire                _zz_dataOut_payload_0_5733;
  wire       [7:0]    _zz_dataOut_payload_0_5734;
  wire       [7:0]    _zz_dataOut_payload_0_5735;
  wire                _zz_dataOut_payload_0_5736;
  wire       [7:0]    _zz_dataOut_payload_0_5737;
  wire       [7:0]    _zz_dataOut_payload_0_5738;
  wire                _zz_dataOut_payload_0_5739;
  wire       [7:0]    _zz_dataOut_payload_0_5740;
  wire       [7:0]    _zz_dataOut_payload_0_5741;
  wire                _zz_dataOut_payload_0_5742;
  wire       [7:0]    _zz_dataOut_payload_0_5743;
  wire       [7:0]    _zz_dataOut_payload_0_5744;
  wire                _zz_dataOut_payload_0_5745;
  wire       [7:0]    _zz_dataOut_payload_0_5746;
  wire       [7:0]    _zz_dataOut_payload_0_5747;
  wire                _zz_dataOut_payload_0_5748;
  wire       [7:0]    _zz_dataOut_payload_0_5749;
  wire       [7:0]    _zz_dataOut_payload_0_5750;
  wire                _zz_dataOut_payload_0_5751;
  wire       [7:0]    _zz_dataOut_payload_0_5752;
  wire       [7:0]    _zz_dataOut_payload_0_5753;
  wire                _zz_dataOut_payload_0_5754;
  wire       [7:0]    _zz_dataOut_payload_0_5755;
  wire       [7:0]    _zz_dataOut_payload_0_5756;
  wire                _zz_dataOut_payload_0_5757;
  wire       [7:0]    _zz_dataOut_payload_0_5758;
  wire       [7:0]    _zz_dataOut_payload_0_5759;
  wire                _zz_dataOut_payload_0_5760;
  wire       [7:0]    _zz_dataOut_payload_0_5761;
  wire       [7:0]    _zz_dataOut_payload_0_5762;
  wire                _zz_dataOut_payload_0_5763;
  wire       [7:0]    _zz_dataOut_payload_0_5764;
  wire       [7:0]    _zz_dataOut_payload_0_5765;
  wire                _zz_dataOut_payload_0_5766;
  wire       [7:0]    _zz_dataOut_payload_0_5767;
  wire       [7:0]    _zz_dataOut_payload_0_5768;
  wire                _zz_dataOut_payload_0_5769;
  wire       [7:0]    _zz_dataOut_payload_0_5770;
  wire       [7:0]    _zz_dataOut_payload_0_5771;
  wire                _zz_dataOut_payload_0_5772;
  wire       [7:0]    _zz_dataOut_payload_0_5773;
  wire       [7:0]    _zz_dataOut_payload_0_5774;
  wire                _zz_dataOut_payload_0_5775;
  wire       [7:0]    _zz_dataOut_payload_0_5776;
  wire       [7:0]    _zz_dataOut_payload_0_5777;
  wire                _zz_dataOut_payload_0_5778;
  wire       [7:0]    _zz_dataOut_payload_0_5779;
  wire       [7:0]    _zz_dataOut_payload_0_5780;
  wire                _zz_dataOut_payload_0_5781;
  wire       [7:0]    _zz_dataOut_payload_0_5782;
  wire       [7:0]    _zz_dataOut_payload_0_5783;
  wire                _zz_dataOut_payload_0_5784;
  wire       [7:0]    _zz_dataOut_payload_0_5785;
  wire       [7:0]    _zz_dataOut_payload_0_5786;
  wire                _zz_dataOut_payload_0_5787;
  wire       [7:0]    _zz_dataOut_payload_0_5788;
  wire       [7:0]    _zz_dataOut_payload_0_5789;
  wire                _zz_dataOut_payload_0_5790;
  wire       [7:0]    _zz_dataOut_payload_0_5791;
  wire       [7:0]    _zz_dataOut_payload_0_5792;
  wire                _zz_dataOut_payload_0_5793;
  wire       [7:0]    _zz_dataOut_payload_0_5794;
  wire       [7:0]    _zz_dataOut_payload_0_5795;
  wire                _zz_dataOut_payload_0_5796;
  wire       [7:0]    _zz_dataOut_payload_0_5797;
  wire       [7:0]    _zz_dataOut_payload_0_5798;
  wire                _zz_dataOut_payload_0_5799;
  wire       [7:0]    _zz_dataOut_payload_0_5800;
  wire       [7:0]    _zz_dataOut_payload_0_5801;
  wire                _zz_dataOut_payload_0_5802;
  wire                _zz_dataOut_payload_0_5803;
  reg        [7:0]    _zz_dataOut_payload_0_5804;
  reg        [7:0]    _zz_dataOut_payload_0_5805;
  reg        [7:0]    _zz_dataOut_payload_0_5806;
  reg        [7:0]    _zz_dataOut_payload_0_5807;
  wire                _zz_dataOut_payload_0_5808;
  wire       [7:0]    _zz_dataOut_payload_0_5809;
  wire       [7:0]    _zz_dataOut_payload_0_5810;
  wire                _zz_dataOut_payload_0_5811;
  wire       [7:0]    _zz_dataOut_payload_0_5812;
  wire       [7:0]    _zz_dataOut_payload_0_5813;
  wire                _zz_dataOut_payload_0_5814;
  wire                _zz_dataOut_payload_0_5815;
  reg        [7:0]    _zz_dataOut_payload_0_5816;
  reg        [7:0]    _zz_dataOut_payload_0_5817;
  reg        [7:0]    _zz_dataOut_payload_0_5818;
  reg        [7:0]    _zz_dataOut_payload_0_5819;
  reg        [7:0]    _zz_dataOut_payload_0_5820;
  reg        [7:0]    _zz_dataOut_payload_0_5821;
  reg        [7:0]    _zz_dataOut_payload_0_5822;
  reg        [7:0]    _zz_dataOut_payload_0_5823;
  reg        [7:0]    _zz_dataOut_payload_0_5824;
  reg        [7:0]    _zz_dataOut_payload_0_5825;
  reg        [7:0]    _zz_dataOut_payload_0_5826;
  reg        [7:0]    _zz_dataOut_payload_0_5827;
  wire                _zz_dataOut_payload_0_5828;
  wire       [7:0]    _zz_dataOut_payload_0_5829;
  wire       [7:0]    _zz_dataOut_payload_0_5830;
  wire                _zz_dataOut_payload_0_5831;
  wire       [7:0]    _zz_dataOut_payload_0_5832;
  wire       [7:0]    _zz_dataOut_payload_0_5833;
  wire                _zz_dataOut_payload_0_5834;
  wire       [7:0]    _zz_dataOut_payload_0_5835;
  wire       [7:0]    _zz_dataOut_payload_0_5836;
  wire                _zz_dataOut_payload_0_5837;
  wire       [7:0]    _zz_dataOut_payload_0_5838;
  wire       [7:0]    _zz_dataOut_payload_0_5839;
  wire                _zz_dataOut_payload_0_5840;
  wire       [7:0]    _zz_dataOut_payload_0_5841;
  wire       [7:0]    _zz_dataOut_payload_0_5842;
  wire                _zz_dataOut_payload_0_5843;
  wire       [7:0]    _zz_dataOut_payload_0_5844;
  wire       [7:0]    _zz_dataOut_payload_0_5845;
  wire                _zz_dataOut_payload_0_5846;
  wire                _zz_dataOut_payload_0_5847;
  reg        [7:0]    _zz_dataOut_payload_0_5848;
  reg        [7:0]    _zz_dataOut_payload_0_5849;
  reg        [7:0]    _zz_dataOut_payload_0_5850;
  reg        [7:0]    _zz_dataOut_payload_0_5851;
  wire                _zz_dataOut_payload_0_5852;
  wire       [7:0]    _zz_dataOut_payload_0_5853;
  wire       [7:0]    _zz_dataOut_payload_0_5854;
  wire                _zz_dataOut_payload_0_5855;
  wire       [7:0]    _zz_dataOut_payload_0_5856;
  wire       [7:0]    _zz_dataOut_payload_0_5857;
  wire                _zz_dataOut_payload_0_5858;
  wire                _zz_dataOut_payload_0_5859;
  reg        [7:0]    _zz_dataOut_payload_0_5860;
  reg        [7:0]    _zz_dataOut_payload_0_5861;
  reg        [7:0]    _zz_dataOut_payload_0_5862;
  reg        [7:0]    _zz_dataOut_payload_0_5863;
  reg        [7:0]    _zz_dataOut_payload_0_5864;
  reg        [7:0]    _zz_dataOut_payload_0_5865;
  reg        [7:0]    _zz_dataOut_payload_0_5866;
  reg        [7:0]    _zz_dataOut_payload_0_5867;
  reg        [7:0]    _zz_dataOut_payload_0_5868;
  reg        [7:0]    _zz_dataOut_payload_0_5869;
  reg        [7:0]    _zz_dataOut_payload_0_5870;
  reg        [7:0]    _zz_dataOut_payload_0_5871;
  reg        [7:0]    _zz_dataOut_payload_0_5872;
  reg        [7:0]    _zz_dataOut_payload_0_5873;
  reg        [7:0]    _zz_dataOut_payload_0_5874;
  reg        [7:0]    _zz_dataOut_payload_0_5875;
  reg        [7:0]    _zz_dataOut_payload_0_5876;
  reg        [7:0]    _zz_dataOut_payload_0_5877;
  reg        [7:0]    _zz_dataOut_payload_0_5878;
  reg        [7:0]    _zz_dataOut_payload_0_5879;
  reg        [7:0]    _zz_dataOut_payload_0_5880;
  reg        [7:0]    _zz_dataOut_payload_0_5881;
  reg        [7:0]    _zz_dataOut_payload_0_5882;
  reg        [7:0]    _zz_dataOut_payload_0_5883;
  reg        [7:0]    _zz_dataOut_payload_0_5884;
  reg        [7:0]    _zz_dataOut_payload_0_5885;
  reg        [7:0]    _zz_dataOut_payload_0_5886;
  reg        [7:0]    _zz_dataOut_payload_0_5887;
  wire                _zz_dataOut_payload_0_5888;
  wire       [7:0]    _zz_dataOut_payload_0_5889;
  wire       [7:0]    _zz_dataOut_payload_0_5890;
  wire                _zz_dataOut_payload_0_5891;
  wire       [7:0]    _zz_dataOut_payload_0_5892;
  wire       [7:0]    _zz_dataOut_payload_0_5893;
  wire                _zz_dataOut_payload_0_5894;
  wire       [7:0]    _zz_dataOut_payload_0_5895;
  wire       [7:0]    _zz_dataOut_payload_0_5896;
  wire                _zz_dataOut_payload_0_5897;
  wire       [7:0]    _zz_dataOut_payload_0_5898;
  wire       [7:0]    _zz_dataOut_payload_0_5899;
  wire                _zz_dataOut_payload_0_5900;
  wire       [7:0]    _zz_dataOut_payload_0_5901;
  wire       [7:0]    _zz_dataOut_payload_0_5902;
  wire                _zz_dataOut_payload_0_5903;
  wire       [7:0]    _zz_dataOut_payload_0_5904;
  wire       [7:0]    _zz_dataOut_payload_0_5905;
  wire                _zz_dataOut_payload_0_5906;
  wire       [7:0]    _zz_dataOut_payload_0_5907;
  wire       [7:0]    _zz_dataOut_payload_0_5908;
  wire                _zz_dataOut_payload_0_5909;
  wire       [7:0]    _zz_dataOut_payload_0_5910;
  wire       [7:0]    _zz_dataOut_payload_0_5911;
  wire                _zz_dataOut_payload_0_5912;
  wire       [7:0]    _zz_dataOut_payload_0_5913;
  wire       [7:0]    _zz_dataOut_payload_0_5914;
  wire                _zz_dataOut_payload_0_5915;
  wire       [7:0]    _zz_dataOut_payload_0_5916;
  wire       [7:0]    _zz_dataOut_payload_0_5917;
  wire                _zz_dataOut_payload_0_5918;
  wire       [7:0]    _zz_dataOut_payload_0_5919;
  wire       [7:0]    _zz_dataOut_payload_0_5920;
  wire                _zz_dataOut_payload_0_5921;
  wire       [7:0]    _zz_dataOut_payload_0_5922;
  wire       [7:0]    _zz_dataOut_payload_0_5923;
  wire                _zz_dataOut_payload_0_5924;
  wire       [7:0]    _zz_dataOut_payload_0_5925;
  wire       [7:0]    _zz_dataOut_payload_0_5926;
  wire                _zz_dataOut_payload_0_5927;
  wire       [7:0]    _zz_dataOut_payload_0_5928;
  wire       [7:0]    _zz_dataOut_payload_0_5929;
  wire                _zz_dataOut_payload_0_5930;
  wire                _zz_dataOut_payload_0_5931;
  reg        [7:0]    _zz_dataOut_payload_0_5932;
  reg        [7:0]    _zz_dataOut_payload_0_5933;
  reg        [7:0]    _zz_dataOut_payload_0_5934;
  reg        [7:0]    _zz_dataOut_payload_0_5935;
  wire                _zz_dataOut_payload_0_5936;
  wire       [7:0]    _zz_dataOut_payload_0_5937;
  wire       [7:0]    _zz_dataOut_payload_0_5938;
  wire                _zz_dataOut_payload_0_5939;
  wire       [7:0]    _zz_dataOut_payload_0_5940;
  wire       [7:0]    _zz_dataOut_payload_0_5941;
  wire                _zz_dataOut_payload_0_5942;
  wire                _zz_dataOut_payload_0_5943;
  reg        [7:0]    _zz_dataOut_payload_0_5944;
  reg        [7:0]    _zz_dataOut_payload_0_5945;
  reg        [7:0]    _zz_dataOut_payload_0_5946;
  reg        [7:0]    _zz_dataOut_payload_0_5947;
  reg        [7:0]    _zz_dataOut_payload_0_5948;
  reg        [7:0]    _zz_dataOut_payload_0_5949;
  reg        [7:0]    _zz_dataOut_payload_0_5950;
  reg        [7:0]    _zz_dataOut_payload_0_5951;
  reg        [7:0]    _zz_dataOut_payload_0_5952;
  reg        [7:0]    _zz_dataOut_payload_0_5953;
  reg        [7:0]    _zz_dataOut_payload_0_5954;
  reg        [7:0]    _zz_dataOut_payload_0_5955;
  wire                _zz_dataOut_payload_0_5956;
  wire       [7:0]    _zz_dataOut_payload_0_5957;
  wire       [7:0]    _zz_dataOut_payload_0_5958;
  wire                _zz_dataOut_payload_0_5959;
  wire       [7:0]    _zz_dataOut_payload_0_5960;
  wire       [7:0]    _zz_dataOut_payload_0_5961;
  wire                _zz_dataOut_payload_0_5962;
  wire       [7:0]    _zz_dataOut_payload_0_5963;
  wire       [7:0]    _zz_dataOut_payload_0_5964;
  wire                _zz_dataOut_payload_0_5965;
  wire       [7:0]    _zz_dataOut_payload_0_5966;
  wire       [7:0]    _zz_dataOut_payload_0_5967;
  wire                _zz_dataOut_payload_0_5968;
  wire       [7:0]    _zz_dataOut_payload_0_5969;
  wire       [7:0]    _zz_dataOut_payload_0_5970;
  wire                _zz_dataOut_payload_0_5971;
  wire       [7:0]    _zz_dataOut_payload_0_5972;
  wire       [7:0]    _zz_dataOut_payload_0_5973;
  wire                _zz_dataOut_payload_0_5974;
  wire                _zz_dataOut_payload_0_5975;
  reg        [7:0]    _zz_dataOut_payload_0_5976;
  reg        [7:0]    _zz_dataOut_payload_0_5977;
  reg        [7:0]    _zz_dataOut_payload_0_5978;
  reg        [7:0]    _zz_dataOut_payload_0_5979;
  wire                _zz_dataOut_payload_0_5980;
  wire       [7:0]    _zz_dataOut_payload_0_5981;
  wire       [7:0]    _zz_dataOut_payload_0_5982;
  wire                _zz_dataOut_payload_0_5983;
  wire       [7:0]    _zz_dataOut_payload_0_5984;
  wire       [7:0]    _zz_dataOut_payload_0_5985;
  wire                _zz_dataOut_payload_0_5986;
  wire                _zz_dataOut_payload_0_5987;
  reg        [7:0]    _zz_dataOut_payload_0_5988;
  reg        [7:0]    _zz_dataOut_payload_0_5989;
  reg        [7:0]    _zz_dataOut_payload_0_5990;
  reg        [7:0]    _zz_dataOut_payload_0_5991;
  reg        [7:0]    _zz_dataOut_payload_0_5992;
  reg        [7:0]    _zz_dataOut_payload_0_5993;
  reg        [7:0]    _zz_dataOut_payload_0_5994;
  reg        [7:0]    _zz_dataOut_payload_0_5995;
  reg        [7:0]    _zz_dataOut_payload_0_5996;
  reg        [7:0]    _zz_dataOut_payload_0_5997;
  reg        [7:0]    _zz_dataOut_payload_0_5998;
  reg        [7:0]    _zz_dataOut_payload_0_5999;
  reg        [7:0]    _zz_dataOut_payload_0_6000;
  reg        [7:0]    _zz_dataOut_payload_0_6001;
  reg        [7:0]    _zz_dataOut_payload_0_6002;
  reg        [7:0]    _zz_dataOut_payload_0_6003;
  reg        [7:0]    _zz_dataOut_payload_0_6004;
  reg        [7:0]    _zz_dataOut_payload_0_6005;
  reg        [7:0]    _zz_dataOut_payload_0_6006;
  reg        [7:0]    _zz_dataOut_payload_0_6007;
  reg        [7:0]    _zz_dataOut_payload_0_6008;
  reg        [7:0]    _zz_dataOut_payload_0_6009;
  reg        [7:0]    _zz_dataOut_payload_0_6010;
  reg        [7:0]    _zz_dataOut_payload_0_6011;
  reg        [7:0]    _zz_dataOut_payload_0_6012;
  reg        [7:0]    _zz_dataOut_payload_0_6013;
  reg        [7:0]    _zz_dataOut_payload_0_6014;
  reg        [7:0]    _zz_dataOut_payload_0_6015;
  reg        [7:0]    _zz_dataOut_payload_0_6016;
  reg        [7:0]    _zz_dataOut_payload_0_6017;
  reg        [7:0]    _zz_dataOut_payload_0_6018;
  reg        [7:0]    _zz_dataOut_payload_0_6019;
  reg        [7:0]    _zz_dataOut_payload_0_6020;
  reg        [7:0]    _zz_dataOut_payload_0_6021;
  reg        [7:0]    _zz_dataOut_payload_0_6022;
  reg        [7:0]    _zz_dataOut_payload_0_6023;
  reg        [7:0]    _zz_dataOut_payload_0_6024;
  reg        [7:0]    _zz_dataOut_payload_0_6025;
  reg        [7:0]    _zz_dataOut_payload_0_6026;
  reg        [7:0]    _zz_dataOut_payload_0_6027;
  reg        [7:0]    _zz_dataOut_payload_0_6028;
  reg        [7:0]    _zz_dataOut_payload_0_6029;
  reg        [7:0]    _zz_dataOut_payload_0_6030;
  reg        [7:0]    _zz_dataOut_payload_0_6031;
  reg        [7:0]    _zz_dataOut_payload_0_6032;
  reg        [7:0]    _zz_dataOut_payload_0_6033;
  reg        [7:0]    _zz_dataOut_payload_0_6034;
  reg        [7:0]    _zz_dataOut_payload_0_6035;
  reg        [7:0]    _zz_dataOut_payload_0_6036;
  reg        [7:0]    _zz_dataOut_payload_0_6037;
  reg        [7:0]    _zz_dataOut_payload_0_6038;
  reg        [7:0]    _zz_dataOut_payload_0_6039;
  reg        [7:0]    _zz_dataOut_payload_0_6040;
  reg        [7:0]    _zz_dataOut_payload_0_6041;
  reg        [7:0]    _zz_dataOut_payload_0_6042;
  reg        [7:0]    _zz_dataOut_payload_0_6043;
  reg        [7:0]    _zz_dataOut_payload_0_6044;
  reg        [7:0]    _zz_dataOut_payload_0_6045;
  reg        [7:0]    _zz_dataOut_payload_0_6046;
  reg        [7:0]    _zz_dataOut_payload_0_6047;
  wire                _zz_dataOut_payload_0_6048;
  wire       [7:0]    _zz_dataOut_payload_0_6049;
  wire       [7:0]    _zz_dataOut_payload_0_6050;
  wire                _zz_dataOut_payload_0_6051;
  wire       [7:0]    _zz_dataOut_payload_0_6052;
  wire       [7:0]    _zz_dataOut_payload_0_6053;
  wire                _zz_dataOut_payload_0_6054;
  wire       [7:0]    _zz_dataOut_payload_0_6055;
  wire       [7:0]    _zz_dataOut_payload_0_6056;
  wire                _zz_dataOut_payload_0_6057;
  wire       [7:0]    _zz_dataOut_payload_0_6058;
  wire       [7:0]    _zz_dataOut_payload_0_6059;
  wire                _zz_dataOut_payload_0_6060;
  wire       [7:0]    _zz_dataOut_payload_0_6061;
  wire       [7:0]    _zz_dataOut_payload_0_6062;
  wire                _zz_dataOut_payload_0_6063;
  wire       [7:0]    _zz_dataOut_payload_0_6064;
  wire       [7:0]    _zz_dataOut_payload_0_6065;
  wire                _zz_dataOut_payload_0_6066;
  wire       [7:0]    _zz_dataOut_payload_0_6067;
  wire       [7:0]    _zz_dataOut_payload_0_6068;
  wire                _zz_dataOut_payload_0_6069;
  wire       [7:0]    _zz_dataOut_payload_0_6070;
  wire       [7:0]    _zz_dataOut_payload_0_6071;
  wire                _zz_dataOut_payload_0_6072;
  wire       [7:0]    _zz_dataOut_payload_0_6073;
  wire       [7:0]    _zz_dataOut_payload_0_6074;
  wire                _zz_dataOut_payload_0_6075;
  wire       [7:0]    _zz_dataOut_payload_0_6076;
  wire       [7:0]    _zz_dataOut_payload_0_6077;
  wire                _zz_dataOut_payload_0_6078;
  wire       [7:0]    _zz_dataOut_payload_0_6079;
  wire       [7:0]    _zz_dataOut_payload_0_6080;
  wire                _zz_dataOut_payload_0_6081;
  wire       [7:0]    _zz_dataOut_payload_0_6082;
  wire       [7:0]    _zz_dataOut_payload_0_6083;
  wire                _zz_dataOut_payload_0_6084;
  wire       [7:0]    _zz_dataOut_payload_0_6085;
  wire       [7:0]    _zz_dataOut_payload_0_6086;
  wire                _zz_dataOut_payload_0_6087;
  wire       [7:0]    _zz_dataOut_payload_0_6088;
  wire       [7:0]    _zz_dataOut_payload_0_6089;
  wire                _zz_dataOut_payload_0_6090;
  wire       [7:0]    _zz_dataOut_payload_0_6091;
  wire       [7:0]    _zz_dataOut_payload_0_6092;
  wire                _zz_dataOut_payload_0_6093;
  wire       [7:0]    _zz_dataOut_payload_0_6094;
  wire       [7:0]    _zz_dataOut_payload_0_6095;
  wire                _zz_dataOut_payload_0_6096;
  wire       [7:0]    _zz_dataOut_payload_0_6097;
  wire       [7:0]    _zz_dataOut_payload_0_6098;
  wire                _zz_dataOut_payload_0_6099;
  wire       [7:0]    _zz_dataOut_payload_0_6100;
  wire       [7:0]    _zz_dataOut_payload_0_6101;
  wire                _zz_dataOut_payload_0_6102;
  wire       [7:0]    _zz_dataOut_payload_0_6103;
  wire       [7:0]    _zz_dataOut_payload_0_6104;
  wire                _zz_dataOut_payload_0_6105;
  wire       [7:0]    _zz_dataOut_payload_0_6106;
  wire       [7:0]    _zz_dataOut_payload_0_6107;
  wire                _zz_dataOut_payload_0_6108;
  wire       [7:0]    _zz_dataOut_payload_0_6109;
  wire       [7:0]    _zz_dataOut_payload_0_6110;
  wire                _zz_dataOut_payload_0_6111;
  wire       [7:0]    _zz_dataOut_payload_0_6112;
  wire       [7:0]    _zz_dataOut_payload_0_6113;
  wire                _zz_dataOut_payload_0_6114;
  wire       [7:0]    _zz_dataOut_payload_0_6115;
  wire       [7:0]    _zz_dataOut_payload_0_6116;
  wire                _zz_dataOut_payload_0_6117;
  wire       [7:0]    _zz_dataOut_payload_0_6118;
  wire       [7:0]    _zz_dataOut_payload_0_6119;
  wire                _zz_dataOut_payload_0_6120;
  wire       [7:0]    _zz_dataOut_payload_0_6121;
  wire       [7:0]    _zz_dataOut_payload_0_6122;
  wire                _zz_dataOut_payload_0_6123;
  wire       [7:0]    _zz_dataOut_payload_0_6124;
  wire       [7:0]    _zz_dataOut_payload_0_6125;
  wire                _zz_dataOut_payload_0_6126;
  wire       [7:0]    _zz_dataOut_payload_0_6127;
  wire       [7:0]    _zz_dataOut_payload_0_6128;
  wire                _zz_dataOut_payload_0_6129;
  wire       [7:0]    _zz_dataOut_payload_0_6130;
  wire       [7:0]    _zz_dataOut_payload_0_6131;
  wire                _zz_dataOut_payload_0_6132;
  wire       [7:0]    _zz_dataOut_payload_0_6133;
  wire       [7:0]    _zz_dataOut_payload_0_6134;
  wire                _zz_dataOut_payload_0_6135;
  wire       [7:0]    _zz_dataOut_payload_0_6136;
  wire       [7:0]    _zz_dataOut_payload_0_6137;
  wire                _zz_dataOut_payload_0_6138;
  wire                _zz_dataOut_payload_0_6139;
  reg        [7:0]    _zz_dataOut_payload_0_6140;
  reg        [7:0]    _zz_dataOut_payload_0_6141;
  reg        [7:0]    _zz_dataOut_payload_0_6142;
  reg        [7:0]    _zz_dataOut_payload_0_6143;
  wire                _zz_dataOut_payload_0_6144;
  wire       [7:0]    _zz_dataOut_payload_0_6145;
  wire       [7:0]    _zz_dataOut_payload_0_6146;
  wire                _zz_dataOut_payload_0_6147;
  wire       [7:0]    _zz_dataOut_payload_0_6148;
  wire       [7:0]    _zz_dataOut_payload_0_6149;
  wire                _zz_dataOut_payload_0_6150;
  wire                _zz_dataOut_payload_0_6151;
  reg        [7:0]    _zz_dataOut_payload_0_6152;
  reg        [7:0]    _zz_dataOut_payload_0_6153;
  reg        [7:0]    _zz_dataOut_payload_0_6154;
  reg        [7:0]    _zz_dataOut_payload_0_6155;
  reg        [7:0]    _zz_dataOut_payload_0_6156;
  reg        [7:0]    _zz_dataOut_payload_0_6157;
  reg        [7:0]    _zz_dataOut_payload_0_6158;
  reg        [7:0]    _zz_dataOut_payload_0_6159;
  reg        [7:0]    _zz_dataOut_payload_0_6160;
  reg        [7:0]    _zz_dataOut_payload_0_6161;
  reg        [7:0]    _zz_dataOut_payload_0_6162;
  reg        [7:0]    _zz_dataOut_payload_0_6163;
  wire                _zz_dataOut_payload_0_6164;
  wire       [7:0]    _zz_dataOut_payload_0_6165;
  wire       [7:0]    _zz_dataOut_payload_0_6166;
  wire                _zz_dataOut_payload_0_6167;
  wire       [7:0]    _zz_dataOut_payload_0_6168;
  wire       [7:0]    _zz_dataOut_payload_0_6169;
  wire                _zz_dataOut_payload_0_6170;
  wire       [7:0]    _zz_dataOut_payload_0_6171;
  wire       [7:0]    _zz_dataOut_payload_0_6172;
  wire                _zz_dataOut_payload_0_6173;
  wire       [7:0]    _zz_dataOut_payload_0_6174;
  wire       [7:0]    _zz_dataOut_payload_0_6175;
  wire                _zz_dataOut_payload_0_6176;
  wire       [7:0]    _zz_dataOut_payload_0_6177;
  wire       [7:0]    _zz_dataOut_payload_0_6178;
  wire                _zz_dataOut_payload_0_6179;
  wire       [7:0]    _zz_dataOut_payload_0_6180;
  wire       [7:0]    _zz_dataOut_payload_0_6181;
  wire                _zz_dataOut_payload_0_6182;
  wire                _zz_dataOut_payload_0_6183;
  reg        [7:0]    _zz_dataOut_payload_0_6184;
  reg        [7:0]    _zz_dataOut_payload_0_6185;
  reg        [7:0]    _zz_dataOut_payload_0_6186;
  reg        [7:0]    _zz_dataOut_payload_0_6187;
  wire                _zz_dataOut_payload_0_6188;
  wire       [7:0]    _zz_dataOut_payload_0_6189;
  wire       [7:0]    _zz_dataOut_payload_0_6190;
  wire                _zz_dataOut_payload_0_6191;
  wire       [7:0]    _zz_dataOut_payload_0_6192;
  wire       [7:0]    _zz_dataOut_payload_0_6193;
  wire                _zz_dataOut_payload_0_6194;
  wire                _zz_dataOut_payload_0_6195;
  reg        [7:0]    _zz_dataOut_payload_0_6196;
  reg        [7:0]    _zz_dataOut_payload_0_6197;
  reg        [7:0]    _zz_dataOut_payload_0_6198;
  reg        [7:0]    _zz_dataOut_payload_0_6199;
  reg        [7:0]    _zz_dataOut_payload_0_6200;
  reg        [7:0]    _zz_dataOut_payload_0_6201;
  reg        [7:0]    _zz_dataOut_payload_0_6202;
  reg        [7:0]    _zz_dataOut_payload_0_6203;
  reg        [7:0]    _zz_dataOut_payload_0_6204;
  reg        [7:0]    _zz_dataOut_payload_0_6205;
  reg        [7:0]    _zz_dataOut_payload_0_6206;
  reg        [7:0]    _zz_dataOut_payload_0_6207;
  reg        [7:0]    _zz_dataOut_payload_0_6208;
  reg        [7:0]    _zz_dataOut_payload_0_6209;
  reg        [7:0]    _zz_dataOut_payload_0_6210;
  reg        [7:0]    _zz_dataOut_payload_0_6211;
  reg        [7:0]    _zz_dataOut_payload_0_6212;
  reg        [7:0]    _zz_dataOut_payload_0_6213;
  reg        [7:0]    _zz_dataOut_payload_0_6214;
  reg        [7:0]    _zz_dataOut_payload_0_6215;
  reg        [7:0]    _zz_dataOut_payload_0_6216;
  reg        [7:0]    _zz_dataOut_payload_0_6217;
  reg        [7:0]    _zz_dataOut_payload_0_6218;
  reg        [7:0]    _zz_dataOut_payload_0_6219;
  reg        [7:0]    _zz_dataOut_payload_0_6220;
  reg        [7:0]    _zz_dataOut_payload_0_6221;
  reg        [7:0]    _zz_dataOut_payload_0_6222;
  reg        [7:0]    _zz_dataOut_payload_0_6223;
  wire                _zz_dataOut_payload_0_6224;
  wire       [7:0]    _zz_dataOut_payload_0_6225;
  wire       [7:0]    _zz_dataOut_payload_0_6226;
  wire                _zz_dataOut_payload_0_6227;
  wire       [7:0]    _zz_dataOut_payload_0_6228;
  wire       [7:0]    _zz_dataOut_payload_0_6229;
  wire                _zz_dataOut_payload_0_6230;
  wire       [7:0]    _zz_dataOut_payload_0_6231;
  wire       [7:0]    _zz_dataOut_payload_0_6232;
  wire                _zz_dataOut_payload_0_6233;
  wire       [7:0]    _zz_dataOut_payload_0_6234;
  wire       [7:0]    _zz_dataOut_payload_0_6235;
  wire                _zz_dataOut_payload_0_6236;
  wire       [7:0]    _zz_dataOut_payload_0_6237;
  wire       [7:0]    _zz_dataOut_payload_0_6238;
  wire                _zz_dataOut_payload_0_6239;
  wire       [7:0]    _zz_dataOut_payload_0_6240;
  wire       [7:0]    _zz_dataOut_payload_0_6241;
  wire                _zz_dataOut_payload_0_6242;
  wire       [7:0]    _zz_dataOut_payload_0_6243;
  wire       [7:0]    _zz_dataOut_payload_0_6244;
  wire                _zz_dataOut_payload_0_6245;
  wire       [7:0]    _zz_dataOut_payload_0_6246;
  wire       [7:0]    _zz_dataOut_payload_0_6247;
  wire                _zz_dataOut_payload_0_6248;
  wire       [7:0]    _zz_dataOut_payload_0_6249;
  wire       [7:0]    _zz_dataOut_payload_0_6250;
  wire                _zz_dataOut_payload_0_6251;
  wire       [7:0]    _zz_dataOut_payload_0_6252;
  wire       [7:0]    _zz_dataOut_payload_0_6253;
  wire                _zz_dataOut_payload_0_6254;
  wire       [7:0]    _zz_dataOut_payload_0_6255;
  wire       [7:0]    _zz_dataOut_payload_0_6256;
  wire                _zz_dataOut_payload_0_6257;
  wire       [7:0]    _zz_dataOut_payload_0_6258;
  wire       [7:0]    _zz_dataOut_payload_0_6259;
  wire                _zz_dataOut_payload_0_6260;
  wire       [7:0]    _zz_dataOut_payload_0_6261;
  wire       [7:0]    _zz_dataOut_payload_0_6262;
  wire                _zz_dataOut_payload_0_6263;
  wire       [7:0]    _zz_dataOut_payload_0_6264;
  wire       [7:0]    _zz_dataOut_payload_0_6265;
  wire                _zz_dataOut_payload_0_6266;
  wire                _zz_dataOut_payload_0_6267;
  reg        [7:0]    _zz_dataOut_payload_0_6268;
  reg        [7:0]    _zz_dataOut_payload_0_6269;
  reg        [7:0]    _zz_dataOut_payload_0_6270;
  reg        [7:0]    _zz_dataOut_payload_0_6271;
  wire                _zz_dataOut_payload_0_6272;
  wire       [7:0]    _zz_dataOut_payload_0_6273;
  wire       [7:0]    _zz_dataOut_payload_0_6274;
  wire                _zz_dataOut_payload_0_6275;
  wire       [7:0]    _zz_dataOut_payload_0_6276;
  wire       [7:0]    _zz_dataOut_payload_0_6277;
  wire                _zz_dataOut_payload_0_6278;
  wire                _zz_dataOut_payload_0_6279;
  reg        [7:0]    _zz_dataOut_payload_0_6280;
  reg        [7:0]    _zz_dataOut_payload_0_6281;
  reg        [7:0]    _zz_dataOut_payload_0_6282;
  reg        [7:0]    _zz_dataOut_payload_0_6283;
  reg        [7:0]    _zz_dataOut_payload_0_6284;
  reg        [7:0]    _zz_dataOut_payload_0_6285;
  reg        [7:0]    _zz_dataOut_payload_0_6286;
  reg        [7:0]    _zz_dataOut_payload_0_6287;
  reg        [7:0]    _zz_dataOut_payload_0_6288;
  reg        [7:0]    _zz_dataOut_payload_0_6289;
  reg        [7:0]    _zz_dataOut_payload_0_6290;
  reg        [7:0]    _zz_dataOut_payload_0_6291;
  wire                _zz_dataOut_payload_0_6292;
  wire       [7:0]    _zz_dataOut_payload_0_6293;
  wire       [7:0]    _zz_dataOut_payload_0_6294;
  wire                _zz_dataOut_payload_0_6295;
  wire       [7:0]    _zz_dataOut_payload_0_6296;
  wire       [7:0]    _zz_dataOut_payload_0_6297;
  wire                _zz_dataOut_payload_0_6298;
  wire       [7:0]    _zz_dataOut_payload_0_6299;
  wire       [7:0]    _zz_dataOut_payload_0_6300;
  wire                _zz_dataOut_payload_0_6301;
  wire       [7:0]    _zz_dataOut_payload_0_6302;
  wire       [7:0]    _zz_dataOut_payload_0_6303;
  wire                _zz_dataOut_payload_0_6304;
  wire       [7:0]    _zz_dataOut_payload_0_6305;
  wire       [7:0]    _zz_dataOut_payload_0_6306;
  wire                _zz_dataOut_payload_0_6307;
  wire       [7:0]    _zz_dataOut_payload_0_6308;
  wire       [7:0]    _zz_dataOut_payload_0_6309;
  wire                _zz_dataOut_payload_0_6310;
  wire                _zz_dataOut_payload_0_6311;
  reg        [7:0]    _zz_dataOut_payload_0_6312;
  reg        [7:0]    _zz_dataOut_payload_0_6313;
  reg        [7:0]    _zz_dataOut_payload_0_6314;
  reg        [7:0]    _zz_dataOut_payload_0_6315;
  wire                _zz_dataOut_payload_0_6316;
  wire       [7:0]    _zz_dataOut_payload_0_6317;
  wire       [7:0]    _zz_dataOut_payload_0_6318;
  wire                _zz_dataOut_payload_0_6319;
  wire       [7:0]    _zz_dataOut_payload_0_6320;
  wire       [7:0]    _zz_dataOut_payload_0_6321;
  wire                _zz_dataOut_payload_0_6322;
  wire                _zz_dataOut_payload_0_6323;
  reg        [7:0]    _zz_dataOut_payload_0_6324;
  reg        [7:0]    _zz_dataOut_payload_0_6325;
  reg        [7:0]    _zz_dataOut_payload_0_6326;
  reg        [7:0]    _zz_dataOut_payload_0_6327;
  reg        [7:0]    _zz_dataOut_payload_0_6328;
  reg        [7:0]    _zz_dataOut_payload_0_6329;
  reg        [7:0]    _zz_dataOut_payload_0_6330;
  reg        [7:0]    _zz_dataOut_payload_0_6331;
  reg        [7:0]    _zz_dataOut_payload_0_6332;
  reg        [7:0]    _zz_dataOut_payload_0_6333;
  reg        [7:0]    _zz_dataOut_payload_0_6334;
  reg        [7:0]    _zz_dataOut_payload_0_6335;
  reg        [7:0]    _zz_dataOut_payload_0_6336;
  reg        [7:0]    _zz_dataOut_payload_0_6337;
  reg        [7:0]    _zz_dataOut_payload_0_6338;
  reg        [7:0]    _zz_dataOut_payload_0_6339;
  reg        [7:0]    _zz_dataOut_payload_0_6340;
  reg        [7:0]    _zz_dataOut_payload_0_6341;
  reg        [7:0]    _zz_dataOut_payload_0_6342;
  reg        [7:0]    _zz_dataOut_payload_0_6343;
  reg        [7:0]    _zz_dataOut_payload_0_6344;
  reg        [7:0]    _zz_dataOut_payload_0_6345;
  reg        [7:0]    _zz_dataOut_payload_0_6346;
  reg        [7:0]    _zz_dataOut_payload_0_6347;
  reg        [7:0]    _zz_dataOut_payload_0_6348;
  reg        [7:0]    _zz_dataOut_payload_0_6349;
  reg        [7:0]    _zz_dataOut_payload_0_6350;
  reg        [7:0]    _zz_dataOut_payload_0_6351;
  reg        [7:0]    _zz_dataOut_payload_0_6352;
  reg        [7:0]    _zz_dataOut_payload_0_6353;
  reg        [7:0]    _zz_dataOut_payload_0_6354;
  reg        [7:0]    _zz_dataOut_payload_0_6355;
  reg        [7:0]    _zz_dataOut_payload_0_6356;
  reg        [7:0]    _zz_dataOut_payload_0_6357;
  reg        [7:0]    _zz_dataOut_payload_0_6358;
  reg        [7:0]    _zz_dataOut_payload_0_6359;
  reg        [7:0]    _zz_dataOut_payload_0_6360;
  reg        [7:0]    _zz_dataOut_payload_0_6361;
  reg        [7:0]    _zz_dataOut_payload_0_6362;
  reg        [7:0]    _zz_dataOut_payload_0_6363;
  reg        [7:0]    _zz_dataOut_payload_0_6364;
  reg        [7:0]    _zz_dataOut_payload_0_6365;
  reg        [7:0]    _zz_dataOut_payload_0_6366;
  reg        [7:0]    _zz_dataOut_payload_0_6367;
  reg        [7:0]    _zz_dataOut_payload_0_6368;
  reg        [7:0]    _zz_dataOut_payload_0_6369;
  reg        [7:0]    _zz_dataOut_payload_0_6370;
  reg        [7:0]    _zz_dataOut_payload_0_6371;
  reg        [7:0]    _zz_dataOut_payload_0_6372;
  reg        [7:0]    _zz_dataOut_payload_0_6373;
  reg        [7:0]    _zz_dataOut_payload_0_6374;
  reg        [7:0]    _zz_dataOut_payload_0_6375;
  reg        [7:0]    _zz_dataOut_payload_0_6376;
  reg        [7:0]    _zz_dataOut_payload_0_6377;
  reg        [7:0]    _zz_dataOut_payload_0_6378;
  reg        [7:0]    _zz_dataOut_payload_0_6379;
  reg        [7:0]    _zz_dataOut_payload_0_6380;
  reg        [7:0]    _zz_dataOut_payload_0_6381;
  reg        [7:0]    _zz_dataOut_payload_0_6382;
  reg        [7:0]    _zz_dataOut_payload_0_6383;
  wire                _zz_dataOut_payload_0_6384;
  wire       [7:0]    _zz_dataOut_payload_0_6385;
  wire       [7:0]    _zz_dataOut_payload_0_6386;
  wire                _zz_dataOut_payload_0_6387;
  wire       [7:0]    _zz_dataOut_payload_0_6388;
  wire       [7:0]    _zz_dataOut_payload_0_6389;
  wire                _zz_dataOut_payload_0_6390;
  wire       [7:0]    _zz_dataOut_payload_0_6391;
  wire       [7:0]    _zz_dataOut_payload_0_6392;
  wire                _zz_dataOut_payload_0_6393;
  wire       [7:0]    _zz_dataOut_payload_0_6394;
  wire       [7:0]    _zz_dataOut_payload_0_6395;
  wire                _zz_dataOut_payload_0_6396;
  wire       [7:0]    _zz_dataOut_payload_0_6397;
  wire       [7:0]    _zz_dataOut_payload_0_6398;
  wire                _zz_dataOut_payload_0_6399;
  wire       [7:0]    _zz_dataOut_payload_0_6400;
  wire       [7:0]    _zz_dataOut_payload_0_6401;
  wire                _zz_dataOut_payload_0_6402;
  wire       [7:0]    _zz_dataOut_payload_0_6403;
  wire       [7:0]    _zz_dataOut_payload_0_6404;
  wire                _zz_dataOut_payload_0_6405;
  wire       [7:0]    _zz_dataOut_payload_0_6406;
  wire       [7:0]    _zz_dataOut_payload_0_6407;
  wire                _zz_dataOut_payload_0_6408;
  wire       [7:0]    _zz_dataOut_payload_0_6409;
  wire       [7:0]    _zz_dataOut_payload_0_6410;
  wire                _zz_dataOut_payload_0_6411;
  wire       [7:0]    _zz_dataOut_payload_0_6412;
  wire       [7:0]    _zz_dataOut_payload_0_6413;
  wire                _zz_dataOut_payload_0_6414;
  wire       [7:0]    _zz_dataOut_payload_0_6415;
  wire       [7:0]    _zz_dataOut_payload_0_6416;
  wire                _zz_dataOut_payload_0_6417;
  wire       [7:0]    _zz_dataOut_payload_0_6418;
  wire       [7:0]    _zz_dataOut_payload_0_6419;
  wire                _zz_dataOut_payload_0_6420;
  wire       [7:0]    _zz_dataOut_payload_0_6421;
  wire       [7:0]    _zz_dataOut_payload_0_6422;
  wire                _zz_dataOut_payload_0_6423;
  wire       [7:0]    _zz_dataOut_payload_0_6424;
  wire       [7:0]    _zz_dataOut_payload_0_6425;
  wire                _zz_dataOut_payload_0_6426;
  wire       [7:0]    _zz_dataOut_payload_0_6427;
  wire       [7:0]    _zz_dataOut_payload_0_6428;
  wire                _zz_dataOut_payload_0_6429;
  wire       [7:0]    _zz_dataOut_payload_0_6430;
  wire       [7:0]    _zz_dataOut_payload_0_6431;
  wire                _zz_dataOut_payload_0_6432;
  wire       [7:0]    _zz_dataOut_payload_0_6433;
  wire       [7:0]    _zz_dataOut_payload_0_6434;
  wire                _zz_dataOut_payload_0_6435;
  wire       [7:0]    _zz_dataOut_payload_0_6436;
  wire       [7:0]    _zz_dataOut_payload_0_6437;
  wire                _zz_dataOut_payload_0_6438;
  wire       [7:0]    _zz_dataOut_payload_0_6439;
  wire       [7:0]    _zz_dataOut_payload_0_6440;
  wire                _zz_dataOut_payload_0_6441;
  wire       [7:0]    _zz_dataOut_payload_0_6442;
  wire       [7:0]    _zz_dataOut_payload_0_6443;
  wire                _zz_dataOut_payload_0_6444;
  wire       [7:0]    _zz_dataOut_payload_0_6445;
  wire       [7:0]    _zz_dataOut_payload_0_6446;
  wire                _zz_dataOut_payload_0_6447;
  wire       [7:0]    _zz_dataOut_payload_0_6448;
  wire       [7:0]    _zz_dataOut_payload_0_6449;
  wire                _zz_dataOut_payload_0_6450;
  wire       [7:0]    _zz_dataOut_payload_0_6451;
  wire       [7:0]    _zz_dataOut_payload_0_6452;
  wire                _zz_dataOut_payload_0_6453;
  wire       [7:0]    _zz_dataOut_payload_0_6454;
  wire       [7:0]    _zz_dataOut_payload_0_6455;
  wire                _zz_dataOut_payload_0_6456;
  wire       [7:0]    _zz_dataOut_payload_0_6457;
  wire       [7:0]    _zz_dataOut_payload_0_6458;
  wire                _zz_dataOut_payload_0_6459;
  wire       [7:0]    _zz_dataOut_payload_0_6460;
  wire       [7:0]    _zz_dataOut_payload_0_6461;
  wire                _zz_dataOut_payload_0_6462;
  wire       [7:0]    _zz_dataOut_payload_0_6463;
  wire       [7:0]    _zz_dataOut_payload_0_6464;
  wire                _zz_dataOut_payload_0_6465;
  wire       [7:0]    _zz_dataOut_payload_0_6466;
  wire       [7:0]    _zz_dataOut_payload_0_6467;
  wire                _zz_dataOut_payload_0_6468;
  wire       [7:0]    _zz_dataOut_payload_0_6469;
  wire       [7:0]    _zz_dataOut_payload_0_6470;
  wire                _zz_dataOut_payload_0_6471;
  wire       [7:0]    _zz_dataOut_payload_0_6472;
  wire       [7:0]    _zz_dataOut_payload_0_6473;
  wire                _zz_dataOut_payload_0_6474;
  wire                _zz_dataOut_payload_0_6475;
  reg        [7:0]    _zz_dataOut_payload_0_6476;
  reg        [7:0]    _zz_dataOut_payload_0_6477;
  reg        [7:0]    _zz_dataOut_payload_0_6478;
  reg        [7:0]    _zz_dataOut_payload_0_6479;
  wire                _zz_dataOut_payload_0_6480;
  wire       [7:0]    _zz_dataOut_payload_0_6481;
  wire       [7:0]    _zz_dataOut_payload_0_6482;
  wire                _zz_dataOut_payload_0_6483;
  wire       [7:0]    _zz_dataOut_payload_0_6484;
  wire       [7:0]    _zz_dataOut_payload_0_6485;
  wire                _zz_dataOut_payload_0_6486;
  wire                _zz_dataOut_payload_0_6487;
  reg        [7:0]    _zz_dataOut_payload_0_6488;
  reg        [7:0]    _zz_dataOut_payload_0_6489;
  reg        [7:0]    _zz_dataOut_payload_0_6490;
  reg        [7:0]    _zz_dataOut_payload_0_6491;
  reg        [7:0]    _zz_dataOut_payload_0_6492;
  reg        [7:0]    _zz_dataOut_payload_0_6493;
  reg        [7:0]    _zz_dataOut_payload_0_6494;
  reg        [7:0]    _zz_dataOut_payload_0_6495;
  reg        [7:0]    _zz_dataOut_payload_0_6496;
  reg        [7:0]    _zz_dataOut_payload_0_6497;
  reg        [7:0]    _zz_dataOut_payload_0_6498;
  reg        [7:0]    _zz_dataOut_payload_0_6499;
  wire                _zz_dataOut_payload_0_6500;
  wire       [7:0]    _zz_dataOut_payload_0_6501;
  wire       [7:0]    _zz_dataOut_payload_0_6502;
  wire                _zz_dataOut_payload_0_6503;
  wire       [7:0]    _zz_dataOut_payload_0_6504;
  wire       [7:0]    _zz_dataOut_payload_0_6505;
  wire                _zz_dataOut_payload_0_6506;
  wire       [7:0]    _zz_dataOut_payload_0_6507;
  wire       [7:0]    _zz_dataOut_payload_0_6508;
  wire                _zz_dataOut_payload_0_6509;
  wire       [7:0]    _zz_dataOut_payload_0_6510;
  wire       [7:0]    _zz_dataOut_payload_0_6511;
  wire                _zz_dataOut_payload_0_6512;
  wire       [7:0]    _zz_dataOut_payload_0_6513;
  wire       [7:0]    _zz_dataOut_payload_0_6514;
  wire                _zz_dataOut_payload_0_6515;
  wire       [7:0]    _zz_dataOut_payload_0_6516;
  wire       [7:0]    _zz_dataOut_payload_0_6517;
  wire                _zz_dataOut_payload_0_6518;
  wire                _zz_dataOut_payload_0_6519;
  reg        [7:0]    _zz_dataOut_payload_0_6520;
  reg        [7:0]    _zz_dataOut_payload_0_6521;
  reg        [7:0]    _zz_dataOut_payload_0_6522;
  reg        [7:0]    _zz_dataOut_payload_0_6523;
  wire                _zz_dataOut_payload_0_6524;
  wire       [7:0]    _zz_dataOut_payload_0_6525;
  wire       [7:0]    _zz_dataOut_payload_0_6526;
  wire                _zz_dataOut_payload_0_6527;
  wire       [7:0]    _zz_dataOut_payload_0_6528;
  wire       [7:0]    _zz_dataOut_payload_0_6529;
  wire                _zz_dataOut_payload_0_6530;
  wire                _zz_dataOut_payload_0_6531;
  reg        [7:0]    _zz_dataOut_payload_0_6532;
  reg        [7:0]    _zz_dataOut_payload_0_6533;
  reg        [7:0]    _zz_dataOut_payload_0_6534;
  reg        [7:0]    _zz_dataOut_payload_0_6535;
  reg        [7:0]    _zz_dataOut_payload_0_6536;
  reg        [7:0]    _zz_dataOut_payload_0_6537;
  reg        [7:0]    _zz_dataOut_payload_0_6538;
  reg        [7:0]    _zz_dataOut_payload_0_6539;
  reg        [7:0]    _zz_dataOut_payload_0_6540;
  reg        [7:0]    _zz_dataOut_payload_0_6541;
  reg        [7:0]    _zz_dataOut_payload_0_6542;
  reg        [7:0]    _zz_dataOut_payload_0_6543;
  reg        [7:0]    _zz_dataOut_payload_0_6544;
  reg        [7:0]    _zz_dataOut_payload_0_6545;
  reg        [7:0]    _zz_dataOut_payload_0_6546;
  reg        [7:0]    _zz_dataOut_payload_0_6547;
  reg        [7:0]    _zz_dataOut_payload_0_6548;
  reg        [7:0]    _zz_dataOut_payload_0_6549;
  reg        [7:0]    _zz_dataOut_payload_0_6550;
  reg        [7:0]    _zz_dataOut_payload_0_6551;
  reg        [7:0]    _zz_dataOut_payload_0_6552;
  reg        [7:0]    _zz_dataOut_payload_0_6553;
  reg        [7:0]    _zz_dataOut_payload_0_6554;
  reg        [7:0]    _zz_dataOut_payload_0_6555;
  reg        [7:0]    _zz_dataOut_payload_0_6556;
  reg        [7:0]    _zz_dataOut_payload_0_6557;
  reg        [7:0]    _zz_dataOut_payload_0_6558;
  reg        [7:0]    _zz_dataOut_payload_0_6559;
  wire                _zz_dataOut_payload_0_6560;
  wire       [7:0]    _zz_dataOut_payload_0_6561;
  wire       [7:0]    _zz_dataOut_payload_0_6562;
  wire                _zz_dataOut_payload_0_6563;
  wire       [7:0]    _zz_dataOut_payload_0_6564;
  wire       [7:0]    _zz_dataOut_payload_0_6565;
  wire                _zz_dataOut_payload_0_6566;
  wire       [7:0]    _zz_dataOut_payload_0_6567;
  wire       [7:0]    _zz_dataOut_payload_0_6568;
  wire                _zz_dataOut_payload_0_6569;
  wire       [7:0]    _zz_dataOut_payload_0_6570;
  wire       [7:0]    _zz_dataOut_payload_0_6571;
  wire                _zz_dataOut_payload_0_6572;
  wire       [7:0]    _zz_dataOut_payload_0_6573;
  wire       [7:0]    _zz_dataOut_payload_0_6574;
  wire                _zz_dataOut_payload_0_6575;
  wire       [7:0]    _zz_dataOut_payload_0_6576;
  wire       [7:0]    _zz_dataOut_payload_0_6577;
  wire                _zz_dataOut_payload_0_6578;
  wire       [7:0]    _zz_dataOut_payload_0_6579;
  wire       [7:0]    _zz_dataOut_payload_0_6580;
  wire                _zz_dataOut_payload_0_6581;
  wire       [7:0]    _zz_dataOut_payload_0_6582;
  wire       [7:0]    _zz_dataOut_payload_0_6583;
  wire                _zz_dataOut_payload_0_6584;
  wire       [7:0]    _zz_dataOut_payload_0_6585;
  wire       [7:0]    _zz_dataOut_payload_0_6586;
  wire                _zz_dataOut_payload_0_6587;
  wire       [7:0]    _zz_dataOut_payload_0_6588;
  wire       [7:0]    _zz_dataOut_payload_0_6589;
  wire                _zz_dataOut_payload_0_6590;
  wire       [7:0]    _zz_dataOut_payload_0_6591;
  wire       [7:0]    _zz_dataOut_payload_0_6592;
  wire                _zz_dataOut_payload_0_6593;
  wire       [7:0]    _zz_dataOut_payload_0_6594;
  wire       [7:0]    _zz_dataOut_payload_0_6595;
  wire                _zz_dataOut_payload_0_6596;
  wire       [7:0]    _zz_dataOut_payload_0_6597;
  wire       [7:0]    _zz_dataOut_payload_0_6598;
  wire                _zz_dataOut_payload_0_6599;
  wire       [7:0]    _zz_dataOut_payload_0_6600;
  wire       [7:0]    _zz_dataOut_payload_0_6601;
  wire                _zz_dataOut_payload_0_6602;
  wire                _zz_dataOut_payload_0_6603;
  reg        [7:0]    _zz_dataOut_payload_0_6604;
  reg        [7:0]    _zz_dataOut_payload_0_6605;
  reg        [7:0]    _zz_dataOut_payload_0_6606;
  reg        [7:0]    _zz_dataOut_payload_0_6607;
  wire                _zz_dataOut_payload_0_6608;
  wire       [7:0]    _zz_dataOut_payload_0_6609;
  wire       [7:0]    _zz_dataOut_payload_0_6610;
  wire                _zz_dataOut_payload_0_6611;
  wire       [7:0]    _zz_dataOut_payload_0_6612;
  wire       [7:0]    _zz_dataOut_payload_0_6613;
  wire                _zz_dataOut_payload_0_6614;
  wire                _zz_dataOut_payload_0_6615;
  reg        [7:0]    _zz_dataOut_payload_0_6616;
  reg        [7:0]    _zz_dataOut_payload_0_6617;
  reg        [7:0]    _zz_dataOut_payload_0_6618;
  reg        [7:0]    _zz_dataOut_payload_0_6619;
  reg        [7:0]    _zz_dataOut_payload_0_6620;
  reg        [7:0]    _zz_dataOut_payload_0_6621;
  reg        [7:0]    _zz_dataOut_payload_0_6622;
  reg        [7:0]    _zz_dataOut_payload_0_6623;
  reg        [7:0]    _zz_dataOut_payload_0_6624;
  reg        [7:0]    _zz_dataOut_payload_0_6625;
  reg        [7:0]    _zz_dataOut_payload_0_6626;
  reg        [7:0]    _zz_dataOut_payload_0_6627;
  wire                _zz_dataOut_payload_0_6628;
  wire       [7:0]    _zz_dataOut_payload_0_6629;
  wire       [7:0]    _zz_dataOut_payload_0_6630;
  wire                _zz_dataOut_payload_0_6631;
  wire       [7:0]    _zz_dataOut_payload_0_6632;
  wire       [7:0]    _zz_dataOut_payload_0_6633;
  wire                _zz_dataOut_payload_0_6634;
  wire       [7:0]    _zz_dataOut_payload_0_6635;
  wire       [7:0]    _zz_dataOut_payload_0_6636;
  wire                _zz_dataOut_payload_0_6637;
  wire       [7:0]    _zz_dataOut_payload_0_6638;
  wire       [7:0]    _zz_dataOut_payload_0_6639;
  wire                _zz_dataOut_payload_0_6640;
  wire       [7:0]    _zz_dataOut_payload_0_6641;
  wire       [7:0]    _zz_dataOut_payload_0_6642;
  wire                _zz_dataOut_payload_0_6643;
  wire       [7:0]    _zz_dataOut_payload_0_6644;
  wire       [7:0]    _zz_dataOut_payload_0_6645;
  wire                _zz_dataOut_payload_0_6646;
  wire                _zz_dataOut_payload_0_6647;
  reg        [7:0]    _zz_dataOut_payload_0_6648;
  reg        [7:0]    _zz_dataOut_payload_0_6649;
  reg        [7:0]    _zz_dataOut_payload_0_6650;
  reg        [7:0]    _zz_dataOut_payload_0_6651;
  wire                _zz_dataOut_payload_0_6652;
  wire       [7:0]    _zz_dataOut_payload_0_6653;
  wire       [7:0]    _zz_dataOut_payload_0_6654;
  wire                _zz_dataOut_payload_0_6655;
  wire       [7:0]    _zz_dataOut_payload_0_6656;
  wire       [7:0]    _zz_dataOut_payload_0_6657;
  wire                _zz_dataOut_payload_0_6658;
  wire                _zz_dataOut_payload_0_6659;
  reg        [7:0]    _zz_dataOut_payload_0_6660;
  reg        [7:0]    _zz_dataOut_payload_0_6661;
  reg        [7:0]    _zz_dataOut_payload_0_6662;
  reg        [7:0]    _zz_dataOut_payload_0_6663;
  reg        [7:0]    _zz_dataOut_payload_0_6664;
  reg        [7:0]    _zz_dataOut_payload_0_6665;
  reg        [7:0]    _zz_dataOut_payload_0_6666;
  reg        [7:0]    _zz_dataOut_payload_0_6667;
  reg        [7:0]    _zz_dataOut_payload_0_6668;
  reg        [7:0]    _zz_dataOut_payload_0_6669;
  reg        [7:0]    _zz_dataOut_payload_0_6670;
  reg        [7:0]    _zz_dataOut_payload_0_6671;
  reg        [7:0]    _zz_dataOut_payload_0_6672;
  reg        [7:0]    _zz_dataOut_payload_0_6673;
  reg        [7:0]    _zz_dataOut_payload_0_6674;
  reg        [7:0]    _zz_dataOut_payload_0_6675;
  reg        [7:0]    _zz_dataOut_payload_0_6676;
  reg        [7:0]    _zz_dataOut_payload_0_6677;
  reg        [7:0]    _zz_dataOut_payload_0_6678;
  reg        [7:0]    _zz_dataOut_payload_0_6679;
  reg        [7:0]    _zz_dataOut_payload_0_6680;
  reg        [7:0]    _zz_dataOut_payload_0_6681;
  reg        [7:0]    _zz_dataOut_payload_0_6682;
  reg        [7:0]    _zz_dataOut_payload_0_6683;
  reg        [7:0]    _zz_dataOut_payload_0_6684;
  reg        [7:0]    _zz_dataOut_payload_0_6685;
  reg        [7:0]    _zz_dataOut_payload_0_6686;
  reg        [7:0]    _zz_dataOut_payload_0_6687;
  reg        [7:0]    _zz_dataOut_payload_0_6688;
  reg        [7:0]    _zz_dataOut_payload_0_6689;
  reg        [7:0]    _zz_dataOut_payload_0_6690;
  reg        [7:0]    _zz_dataOut_payload_0_6691;
  reg        [7:0]    _zz_dataOut_payload_0_6692;
  reg        [7:0]    _zz_dataOut_payload_0_6693;
  reg        [7:0]    _zz_dataOut_payload_0_6694;
  reg        [7:0]    _zz_dataOut_payload_0_6695;
  reg        [7:0]    _zz_dataOut_payload_0_6696;
  reg        [7:0]    _zz_dataOut_payload_0_6697;
  reg        [7:0]    _zz_dataOut_payload_0_6698;
  reg        [7:0]    _zz_dataOut_payload_0_6699;
  reg        [7:0]    _zz_dataOut_payload_0_6700;
  reg        [7:0]    _zz_dataOut_payload_0_6701;
  reg        [7:0]    _zz_dataOut_payload_0_6702;
  reg        [7:0]    _zz_dataOut_payload_0_6703;
  reg        [7:0]    _zz_dataOut_payload_0_6704;
  reg        [7:0]    _zz_dataOut_payload_0_6705;
  reg        [7:0]    _zz_dataOut_payload_0_6706;
  reg        [7:0]    _zz_dataOut_payload_0_6707;
  reg        [7:0]    _zz_dataOut_payload_0_6708;
  reg        [7:0]    _zz_dataOut_payload_0_6709;
  reg        [7:0]    _zz_dataOut_payload_0_6710;
  reg        [7:0]    _zz_dataOut_payload_0_6711;
  reg        [7:0]    _zz_dataOut_payload_0_6712;
  reg        [7:0]    _zz_dataOut_payload_0_6713;
  reg        [7:0]    _zz_dataOut_payload_0_6714;
  reg        [7:0]    _zz_dataOut_payload_0_6715;
  reg        [7:0]    _zz_dataOut_payload_0_6716;
  reg        [7:0]    _zz_dataOut_payload_0_6717;
  reg        [7:0]    _zz_dataOut_payload_0_6718;
  reg        [7:0]    _zz_dataOut_payload_0_6719;
  wire                _zz_dataOut_payload_0_6720;
  wire       [7:0]    _zz_dataOut_payload_0_6721;
  wire       [7:0]    _zz_dataOut_payload_0_6722;
  wire                _zz_dataOut_payload_0_6723;
  wire       [7:0]    _zz_dataOut_payload_0_6724;
  wire       [7:0]    _zz_dataOut_payload_0_6725;
  wire                _zz_dataOut_payload_0_6726;
  wire       [7:0]    _zz_dataOut_payload_0_6727;
  wire       [7:0]    _zz_dataOut_payload_0_6728;
  wire                _zz_dataOut_payload_0_6729;
  wire       [7:0]    _zz_dataOut_payload_0_6730;
  wire       [7:0]    _zz_dataOut_payload_0_6731;
  wire                _zz_dataOut_payload_0_6732;
  wire       [7:0]    _zz_dataOut_payload_0_6733;
  wire       [7:0]    _zz_dataOut_payload_0_6734;
  wire                _zz_dataOut_payload_0_6735;
  wire       [7:0]    _zz_dataOut_payload_0_6736;
  wire       [7:0]    _zz_dataOut_payload_0_6737;
  wire                _zz_dataOut_payload_0_6738;
  wire       [7:0]    _zz_dataOut_payload_0_6739;
  wire       [7:0]    _zz_dataOut_payload_0_6740;
  wire                _zz_dataOut_payload_0_6741;
  wire       [7:0]    _zz_dataOut_payload_0_6742;
  wire       [7:0]    _zz_dataOut_payload_0_6743;
  wire                _zz_dataOut_payload_0_6744;
  wire       [7:0]    _zz_dataOut_payload_0_6745;
  wire       [7:0]    _zz_dataOut_payload_0_6746;
  wire                _zz_dataOut_payload_0_6747;
  wire       [7:0]    _zz_dataOut_payload_0_6748;
  wire       [7:0]    _zz_dataOut_payload_0_6749;
  wire                _zz_dataOut_payload_0_6750;
  wire       [7:0]    _zz_dataOut_payload_0_6751;
  wire       [7:0]    _zz_dataOut_payload_0_6752;
  wire                _zz_dataOut_payload_0_6753;
  wire       [7:0]    _zz_dataOut_payload_0_6754;
  wire       [7:0]    _zz_dataOut_payload_0_6755;
  wire                _zz_dataOut_payload_0_6756;
  wire       [7:0]    _zz_dataOut_payload_0_6757;
  wire       [7:0]    _zz_dataOut_payload_0_6758;
  wire                _zz_dataOut_payload_0_6759;
  wire       [7:0]    _zz_dataOut_payload_0_6760;
  wire       [7:0]    _zz_dataOut_payload_0_6761;
  wire                _zz_dataOut_payload_0_6762;
  wire       [7:0]    _zz_dataOut_payload_0_6763;
  wire       [7:0]    _zz_dataOut_payload_0_6764;
  wire                _zz_dataOut_payload_0_6765;
  wire       [7:0]    _zz_dataOut_payload_0_6766;
  wire       [7:0]    _zz_dataOut_payload_0_6767;
  wire                _zz_dataOut_payload_0_6768;
  wire       [7:0]    _zz_dataOut_payload_0_6769;
  wire       [7:0]    _zz_dataOut_payload_0_6770;
  wire                _zz_dataOut_payload_0_6771;
  wire       [7:0]    _zz_dataOut_payload_0_6772;
  wire       [7:0]    _zz_dataOut_payload_0_6773;
  wire                _zz_dataOut_payload_0_6774;
  wire       [7:0]    _zz_dataOut_payload_0_6775;
  wire       [7:0]    _zz_dataOut_payload_0_6776;
  wire                _zz_dataOut_payload_0_6777;
  wire       [7:0]    _zz_dataOut_payload_0_6778;
  wire       [7:0]    _zz_dataOut_payload_0_6779;
  wire                _zz_dataOut_payload_0_6780;
  wire       [7:0]    _zz_dataOut_payload_0_6781;
  wire       [7:0]    _zz_dataOut_payload_0_6782;
  wire                _zz_dataOut_payload_0_6783;
  wire       [7:0]    _zz_dataOut_payload_0_6784;
  wire       [7:0]    _zz_dataOut_payload_0_6785;
  wire                _zz_dataOut_payload_0_6786;
  wire       [7:0]    _zz_dataOut_payload_0_6787;
  wire       [7:0]    _zz_dataOut_payload_0_6788;
  wire                _zz_dataOut_payload_0_6789;
  wire       [7:0]    _zz_dataOut_payload_0_6790;
  wire       [7:0]    _zz_dataOut_payload_0_6791;
  wire                _zz_dataOut_payload_0_6792;
  wire       [7:0]    _zz_dataOut_payload_0_6793;
  wire       [7:0]    _zz_dataOut_payload_0_6794;
  wire                _zz_dataOut_payload_0_6795;
  wire       [7:0]    _zz_dataOut_payload_0_6796;
  wire       [7:0]    _zz_dataOut_payload_0_6797;
  wire                _zz_dataOut_payload_0_6798;
  wire       [7:0]    _zz_dataOut_payload_0_6799;
  wire       [7:0]    _zz_dataOut_payload_0_6800;
  wire                _zz_dataOut_payload_0_6801;
  wire       [7:0]    _zz_dataOut_payload_0_6802;
  wire       [7:0]    _zz_dataOut_payload_0_6803;
  wire                _zz_dataOut_payload_0_6804;
  wire       [7:0]    _zz_dataOut_payload_0_6805;
  wire       [7:0]    _zz_dataOut_payload_0_6806;
  wire                _zz_dataOut_payload_0_6807;
  wire       [7:0]    _zz_dataOut_payload_0_6808;
  wire       [7:0]    _zz_dataOut_payload_0_6809;
  wire                _zz_dataOut_payload_0_6810;
  wire                _zz_dataOut_payload_0_6811;
  reg        [7:0]    _zz_dataOut_payload_0_6812;
  reg        [7:0]    _zz_dataOut_payload_0_6813;
  reg        [7:0]    _zz_dataOut_payload_0_6814;
  reg        [7:0]    _zz_dataOut_payload_0_6815;
  wire                _zz_dataOut_payload_0_6816;
  wire       [7:0]    _zz_dataOut_payload_0_6817;
  wire       [7:0]    _zz_dataOut_payload_0_6818;
  wire                _zz_dataOut_payload_0_6819;
  wire       [7:0]    _zz_dataOut_payload_0_6820;
  wire       [7:0]    _zz_dataOut_payload_0_6821;
  wire                _zz_dataOut_payload_0_6822;
  wire                _zz_dataOut_payload_0_6823;
  reg        [7:0]    _zz_dataOut_payload_0_6824;
  reg        [7:0]    _zz_dataOut_payload_0_6825;
  reg        [7:0]    _zz_dataOut_payload_0_6826;
  reg        [7:0]    _zz_dataOut_payload_0_6827;
  reg        [7:0]    _zz_dataOut_payload_0_6828;
  reg        [7:0]    _zz_dataOut_payload_0_6829;
  reg        [7:0]    _zz_dataOut_payload_0_6830;
  reg        [7:0]    _zz_dataOut_payload_0_6831;
  reg        [7:0]    _zz_dataOut_payload_0_6832;
  reg        [7:0]    _zz_dataOut_payload_0_6833;
  reg        [7:0]    _zz_dataOut_payload_0_6834;
  reg        [7:0]    _zz_dataOut_payload_0_6835;
  wire                _zz_dataOut_payload_0_6836;
  wire       [7:0]    _zz_dataOut_payload_0_6837;
  wire       [7:0]    _zz_dataOut_payload_0_6838;
  wire                _zz_dataOut_payload_0_6839;
  wire       [7:0]    _zz_dataOut_payload_0_6840;
  wire       [7:0]    _zz_dataOut_payload_0_6841;
  wire                _zz_dataOut_payload_0_6842;
  wire       [7:0]    _zz_dataOut_payload_0_6843;
  wire       [7:0]    _zz_dataOut_payload_0_6844;
  wire                _zz_dataOut_payload_0_6845;
  wire       [7:0]    _zz_dataOut_payload_0_6846;
  wire       [7:0]    _zz_dataOut_payload_0_6847;
  wire                _zz_dataOut_payload_0_6848;
  wire       [7:0]    _zz_dataOut_payload_0_6849;
  wire       [7:0]    _zz_dataOut_payload_0_6850;
  wire                _zz_dataOut_payload_0_6851;
  wire       [7:0]    _zz_dataOut_payload_0_6852;
  wire       [7:0]    _zz_dataOut_payload_0_6853;
  wire                _zz_dataOut_payload_0_6854;
  wire                _zz_dataOut_payload_0_6855;
  reg        [7:0]    _zz_dataOut_payload_0_6856;
  reg        [7:0]    _zz_dataOut_payload_0_6857;
  reg        [7:0]    _zz_dataOut_payload_0_6858;
  reg        [7:0]    _zz_dataOut_payload_0_6859;
  wire                _zz_dataOut_payload_0_6860;
  wire       [7:0]    _zz_dataOut_payload_0_6861;
  wire       [7:0]    _zz_dataOut_payload_0_6862;
  wire                _zz_dataOut_payload_0_6863;
  wire       [7:0]    _zz_dataOut_payload_0_6864;
  wire       [7:0]    _zz_dataOut_payload_0_6865;
  wire                _zz_dataOut_payload_0_6866;
  wire                _zz_dataOut_payload_0_6867;
  reg        [7:0]    _zz_dataOut_payload_0_6868;
  reg        [7:0]    _zz_dataOut_payload_0_6869;
  reg        [7:0]    _zz_dataOut_payload_0_6870;
  reg        [7:0]    _zz_dataOut_payload_0_6871;
  reg        [7:0]    _zz_dataOut_payload_0_6872;
  reg        [7:0]    _zz_dataOut_payload_0_6873;
  reg        [7:0]    _zz_dataOut_payload_0_6874;
  reg        [7:0]    _zz_dataOut_payload_0_6875;
  reg        [7:0]    _zz_dataOut_payload_0_6876;
  reg        [7:0]    _zz_dataOut_payload_0_6877;
  reg        [7:0]    _zz_dataOut_payload_0_6878;
  reg        [7:0]    _zz_dataOut_payload_0_6879;
  reg        [7:0]    _zz_dataOut_payload_0_6880;
  reg        [7:0]    _zz_dataOut_payload_0_6881;
  reg        [7:0]    _zz_dataOut_payload_0_6882;
  reg        [7:0]    _zz_dataOut_payload_0_6883;
  reg        [7:0]    _zz_dataOut_payload_0_6884;
  reg        [7:0]    _zz_dataOut_payload_0_6885;
  reg        [7:0]    _zz_dataOut_payload_0_6886;
  reg        [7:0]    _zz_dataOut_payload_0_6887;
  reg        [7:0]    _zz_dataOut_payload_0_6888;
  reg        [7:0]    _zz_dataOut_payload_0_6889;
  reg        [7:0]    _zz_dataOut_payload_0_6890;
  reg        [7:0]    _zz_dataOut_payload_0_6891;
  reg        [7:0]    _zz_dataOut_payload_0_6892;
  reg        [7:0]    _zz_dataOut_payload_0_6893;
  reg        [7:0]    _zz_dataOut_payload_0_6894;
  reg        [7:0]    _zz_dataOut_payload_0_6895;
  wire                _zz_dataOut_payload_0_6896;
  wire       [7:0]    _zz_dataOut_payload_0_6897;
  wire       [7:0]    _zz_dataOut_payload_0_6898;
  wire                _zz_dataOut_payload_0_6899;
  wire       [7:0]    _zz_dataOut_payload_0_6900;
  wire       [7:0]    _zz_dataOut_payload_0_6901;
  wire                _zz_dataOut_payload_0_6902;
  wire       [7:0]    _zz_dataOut_payload_0_6903;
  wire       [7:0]    _zz_dataOut_payload_0_6904;
  wire                _zz_dataOut_payload_0_6905;
  wire       [7:0]    _zz_dataOut_payload_0_6906;
  wire       [7:0]    _zz_dataOut_payload_0_6907;
  wire                _zz_dataOut_payload_0_6908;
  wire       [7:0]    _zz_dataOut_payload_0_6909;
  wire       [7:0]    _zz_dataOut_payload_0_6910;
  wire                _zz_dataOut_payload_0_6911;
  wire       [7:0]    _zz_dataOut_payload_0_6912;
  wire       [7:0]    _zz_dataOut_payload_0_6913;
  wire                _zz_dataOut_payload_0_6914;
  wire       [7:0]    _zz_dataOut_payload_0_6915;
  wire       [7:0]    _zz_dataOut_payload_0_6916;
  wire                _zz_dataOut_payload_0_6917;
  wire       [7:0]    _zz_dataOut_payload_0_6918;
  wire       [7:0]    _zz_dataOut_payload_0_6919;
  wire                _zz_dataOut_payload_0_6920;
  wire       [7:0]    _zz_dataOut_payload_0_6921;
  wire       [7:0]    _zz_dataOut_payload_0_6922;
  wire                _zz_dataOut_payload_0_6923;
  wire       [7:0]    _zz_dataOut_payload_0_6924;
  wire       [7:0]    _zz_dataOut_payload_0_6925;
  wire                _zz_dataOut_payload_0_6926;
  wire       [7:0]    _zz_dataOut_payload_0_6927;
  wire       [7:0]    _zz_dataOut_payload_0_6928;
  wire                _zz_dataOut_payload_0_6929;
  wire       [7:0]    _zz_dataOut_payload_0_6930;
  wire       [7:0]    _zz_dataOut_payload_0_6931;
  wire                _zz_dataOut_payload_0_6932;
  wire       [7:0]    _zz_dataOut_payload_0_6933;
  wire       [7:0]    _zz_dataOut_payload_0_6934;
  wire                _zz_dataOut_payload_0_6935;
  wire       [7:0]    _zz_dataOut_payload_0_6936;
  wire       [7:0]    _zz_dataOut_payload_0_6937;
  wire                _zz_dataOut_payload_0_6938;
  wire                _zz_dataOut_payload_0_6939;
  reg        [7:0]    _zz_dataOut_payload_0_6940;
  reg        [7:0]    _zz_dataOut_payload_0_6941;
  reg        [7:0]    _zz_dataOut_payload_0_6942;
  reg        [7:0]    _zz_dataOut_payload_0_6943;
  wire                _zz_dataOut_payload_0_6944;
  wire       [7:0]    _zz_dataOut_payload_0_6945;
  wire       [7:0]    _zz_dataOut_payload_0_6946;
  wire                _zz_dataOut_payload_0_6947;
  wire       [7:0]    _zz_dataOut_payload_0_6948;
  wire       [7:0]    _zz_dataOut_payload_0_6949;
  wire                _zz_dataOut_payload_0_6950;
  wire                _zz_dataOut_payload_0_6951;
  reg        [7:0]    _zz_dataOut_payload_0_6952;
  reg        [7:0]    _zz_dataOut_payload_0_6953;
  reg        [7:0]    _zz_dataOut_payload_0_6954;
  reg        [7:0]    _zz_dataOut_payload_0_6955;
  reg        [7:0]    _zz_dataOut_payload_0_6956;
  reg        [7:0]    _zz_dataOut_payload_0_6957;
  reg        [7:0]    _zz_dataOut_payload_0_6958;
  reg        [7:0]    _zz_dataOut_payload_0_6959;
  reg        [7:0]    _zz_dataOut_payload_0_6960;
  reg        [7:0]    _zz_dataOut_payload_0_6961;
  reg        [7:0]    _zz_dataOut_payload_0_6962;
  reg        [7:0]    _zz_dataOut_payload_0_6963;
  wire                _zz_dataOut_payload_0_6964;
  wire       [7:0]    _zz_dataOut_payload_0_6965;
  wire       [7:0]    _zz_dataOut_payload_0_6966;
  wire                _zz_dataOut_payload_0_6967;
  wire       [7:0]    _zz_dataOut_payload_0_6968;
  wire       [7:0]    _zz_dataOut_payload_0_6969;
  wire                _zz_dataOut_payload_0_6970;
  wire       [7:0]    _zz_dataOut_payload_0_6971;
  wire       [7:0]    _zz_dataOut_payload_0_6972;
  wire                _zz_dataOut_payload_0_6973;
  wire       [7:0]    _zz_dataOut_payload_0_6974;
  wire       [7:0]    _zz_dataOut_payload_0_6975;
  wire                _zz_dataOut_payload_0_6976;
  wire       [7:0]    _zz_dataOut_payload_0_6977;
  wire       [7:0]    _zz_dataOut_payload_0_6978;
  wire                _zz_dataOut_payload_0_6979;
  wire       [7:0]    _zz_dataOut_payload_0_6980;
  wire       [7:0]    _zz_dataOut_payload_0_6981;
  wire                _zz_dataOut_payload_0_6982;
  wire                _zz_dataOut_payload_0_6983;
  reg        [7:0]    _zz_dataOut_payload_0_6984;
  reg        [7:0]    _zz_dataOut_payload_0_6985;
  reg        [7:0]    _zz_dataOut_payload_0_6986;
  reg        [7:0]    _zz_dataOut_payload_0_6987;
  wire                _zz_dataOut_payload_0_6988;
  wire       [7:0]    _zz_dataOut_payload_0_6989;
  wire       [7:0]    _zz_dataOut_payload_0_6990;
  wire                _zz_dataOut_payload_0_6991;
  wire       [7:0]    _zz_dataOut_payload_0_6992;
  wire       [7:0]    _zz_dataOut_payload_0_6993;
  wire                _zz_dataOut_payload_0_6994;
  wire                _zz_dataOut_payload_0_6995;
  reg        [7:0]    _zz_dataOut_payload_0_6996;
  reg        [7:0]    _zz_dataOut_payload_0_6997;
  reg        [7:0]    _zz_dataOut_payload_0_6998;
  reg        [7:0]    _zz_dataOut_payload_0_6999;
  reg        [7:0]    _zz_dataOut_payload_0_7000;
  reg        [7:0]    _zz_dataOut_payload_0_7001;
  reg        [7:0]    _zz_dataOut_payload_0_7002;
  reg        [7:0]    _zz_dataOut_payload_0_7003;
  reg        [7:0]    _zz_dataOut_payload_0_7004;
  reg        [7:0]    _zz_dataOut_payload_0_7005;
  reg        [7:0]    _zz_dataOut_payload_0_7006;
  reg        [7:0]    _zz_dataOut_payload_0_7007;
  reg        [7:0]    _zz_dataOut_payload_0_7008;
  reg        [7:0]    _zz_dataOut_payload_0_7009;
  reg        [7:0]    _zz_dataOut_payload_0_7010;
  reg        [7:0]    _zz_dataOut_payload_0_7011;
  reg        [7:0]    _zz_dataOut_payload_0_7012;
  reg        [7:0]    _zz_dataOut_payload_0_7013;
  reg        [7:0]    _zz_dataOut_payload_0_7014;
  reg        [7:0]    _zz_dataOut_payload_0_7015;
  reg        [7:0]    _zz_dataOut_payload_0_7016;
  reg        [7:0]    _zz_dataOut_payload_0_7017;
  reg        [7:0]    _zz_dataOut_payload_0_7018;
  reg        [7:0]    _zz_dataOut_payload_0_7019;
  reg        [7:0]    _zz_dataOut_payload_0_7020;
  reg        [7:0]    _zz_dataOut_payload_0_7021;
  reg        [7:0]    _zz_dataOut_payload_0_7022;
  reg        [7:0]    _zz_dataOut_payload_0_7023;
  reg        [7:0]    _zz_dataOut_payload_0_7024;
  reg        [7:0]    _zz_dataOut_payload_0_7025;
  reg        [7:0]    _zz_dataOut_payload_0_7026;
  reg        [7:0]    _zz_dataOut_payload_0_7027;
  reg        [7:0]    _zz_dataOut_payload_0_7028;
  reg        [7:0]    _zz_dataOut_payload_0_7029;
  reg        [7:0]    _zz_dataOut_payload_0_7030;
  reg        [7:0]    _zz_dataOut_payload_0_7031;
  reg        [7:0]    _zz_dataOut_payload_0_7032;
  reg        [7:0]    _zz_dataOut_payload_0_7033;
  reg        [7:0]    _zz_dataOut_payload_0_7034;
  reg        [7:0]    _zz_dataOut_payload_0_7035;
  reg        [7:0]    _zz_dataOut_payload_0_7036;
  reg        [7:0]    _zz_dataOut_payload_0_7037;
  reg        [7:0]    _zz_dataOut_payload_0_7038;
  reg        [7:0]    _zz_dataOut_payload_0_7039;
  reg        [7:0]    _zz_dataOut_payload_0_7040;
  reg        [7:0]    _zz_dataOut_payload_0_7041;
  reg        [7:0]    _zz_dataOut_payload_0_7042;
  reg        [7:0]    _zz_dataOut_payload_0_7043;
  reg        [7:0]    _zz_dataOut_payload_0_7044;
  reg        [7:0]    _zz_dataOut_payload_0_7045;
  reg        [7:0]    _zz_dataOut_payload_0_7046;
  reg        [7:0]    _zz_dataOut_payload_0_7047;
  reg        [7:0]    _zz_dataOut_payload_0_7048;
  reg        [7:0]    _zz_dataOut_payload_0_7049;
  reg        [7:0]    _zz_dataOut_payload_0_7050;
  reg        [7:0]    _zz_dataOut_payload_0_7051;
  reg        [7:0]    _zz_dataOut_payload_0_7052;
  reg        [7:0]    _zz_dataOut_payload_0_7053;
  reg        [7:0]    _zz_dataOut_payload_0_7054;
  reg        [7:0]    _zz_dataOut_payload_0_7055;
  wire                _zz_dataOut_payload_0_7056;
  wire       [7:0]    _zz_dataOut_payload_0_7057;
  wire       [7:0]    _zz_dataOut_payload_0_7058;
  wire                _zz_dataOut_payload_0_7059;
  wire       [7:0]    _zz_dataOut_payload_0_7060;
  wire       [7:0]    _zz_dataOut_payload_0_7061;
  wire                _zz_dataOut_payload_0_7062;
  wire       [7:0]    _zz_dataOut_payload_0_7063;
  wire       [7:0]    _zz_dataOut_payload_0_7064;
  wire                _zz_dataOut_payload_0_7065;
  wire       [7:0]    _zz_dataOut_payload_0_7066;
  wire       [7:0]    _zz_dataOut_payload_0_7067;
  wire                _zz_dataOut_payload_0_7068;
  wire       [7:0]    _zz_dataOut_payload_0_7069;
  wire       [7:0]    _zz_dataOut_payload_0_7070;
  wire                _zz_dataOut_payload_0_7071;
  wire       [7:0]    _zz_dataOut_payload_0_7072;
  wire       [7:0]    _zz_dataOut_payload_0_7073;
  wire                _zz_dataOut_payload_0_7074;
  wire       [7:0]    _zz_dataOut_payload_0_7075;
  wire       [7:0]    _zz_dataOut_payload_0_7076;
  wire                _zz_dataOut_payload_0_7077;
  wire       [7:0]    _zz_dataOut_payload_0_7078;
  wire       [7:0]    _zz_dataOut_payload_0_7079;
  wire                _zz_dataOut_payload_0_7080;
  wire       [7:0]    _zz_dataOut_payload_0_7081;
  wire       [7:0]    _zz_dataOut_payload_0_7082;
  wire                _zz_dataOut_payload_0_7083;
  wire       [7:0]    _zz_dataOut_payload_0_7084;
  wire       [7:0]    _zz_dataOut_payload_0_7085;
  wire                _zz_dataOut_payload_0_7086;
  wire       [7:0]    _zz_dataOut_payload_0_7087;
  wire       [7:0]    _zz_dataOut_payload_0_7088;
  wire                _zz_dataOut_payload_0_7089;
  wire       [7:0]    _zz_dataOut_payload_0_7090;
  wire       [7:0]    _zz_dataOut_payload_0_7091;
  wire                _zz_dataOut_payload_0_7092;
  wire       [7:0]    _zz_dataOut_payload_0_7093;
  wire       [7:0]    _zz_dataOut_payload_0_7094;
  wire                _zz_dataOut_payload_0_7095;
  wire       [7:0]    _zz_dataOut_payload_0_7096;
  wire       [7:0]    _zz_dataOut_payload_0_7097;
  wire                _zz_dataOut_payload_0_7098;
  wire       [7:0]    _zz_dataOut_payload_0_7099;
  wire       [7:0]    _zz_dataOut_payload_0_7100;
  wire                _zz_dataOut_payload_0_7101;
  wire       [7:0]    _zz_dataOut_payload_0_7102;
  wire       [7:0]    _zz_dataOut_payload_0_7103;
  wire                _zz_dataOut_payload_0_7104;
  wire       [7:0]    _zz_dataOut_payload_0_7105;
  wire       [7:0]    _zz_dataOut_payload_0_7106;
  wire                _zz_dataOut_payload_0_7107;
  wire       [7:0]    _zz_dataOut_payload_0_7108;
  wire       [7:0]    _zz_dataOut_payload_0_7109;
  wire                _zz_dataOut_payload_0_7110;
  wire       [7:0]    _zz_dataOut_payload_0_7111;
  wire       [7:0]    _zz_dataOut_payload_0_7112;
  wire                _zz_dataOut_payload_0_7113;
  wire       [7:0]    _zz_dataOut_payload_0_7114;
  wire       [7:0]    _zz_dataOut_payload_0_7115;
  wire                _zz_dataOut_payload_0_7116;
  wire       [7:0]    _zz_dataOut_payload_0_7117;
  wire       [7:0]    _zz_dataOut_payload_0_7118;
  wire                _zz_dataOut_payload_0_7119;
  wire       [7:0]    _zz_dataOut_payload_0_7120;
  wire       [7:0]    _zz_dataOut_payload_0_7121;
  wire                _zz_dataOut_payload_0_7122;
  wire       [7:0]    _zz_dataOut_payload_0_7123;
  wire       [7:0]    _zz_dataOut_payload_0_7124;
  wire                _zz_dataOut_payload_0_7125;
  wire       [7:0]    _zz_dataOut_payload_0_7126;
  wire       [7:0]    _zz_dataOut_payload_0_7127;
  wire                _zz_dataOut_payload_0_7128;
  wire       [7:0]    _zz_dataOut_payload_0_7129;
  wire       [7:0]    _zz_dataOut_payload_0_7130;
  wire                _zz_dataOut_payload_0_7131;
  wire       [7:0]    _zz_dataOut_payload_0_7132;
  wire       [7:0]    _zz_dataOut_payload_0_7133;
  wire                _zz_dataOut_payload_0_7134;
  wire       [7:0]    _zz_dataOut_payload_0_7135;
  wire       [7:0]    _zz_dataOut_payload_0_7136;
  wire                _zz_dataOut_payload_0_7137;
  wire       [7:0]    _zz_dataOut_payload_0_7138;
  wire       [7:0]    _zz_dataOut_payload_0_7139;
  wire                _zz_dataOut_payload_0_7140;
  wire       [7:0]    _zz_dataOut_payload_0_7141;
  wire       [7:0]    _zz_dataOut_payload_0_7142;
  wire                _zz_dataOut_payload_0_7143;
  wire       [7:0]    _zz_dataOut_payload_0_7144;
  wire       [7:0]    _zz_dataOut_payload_0_7145;
  wire                _zz_dataOut_payload_0_7146;
  wire                _zz_dataOut_payload_0_7147;
  reg        [7:0]    _zz_dataOut_payload_0_7148;
  reg        [7:0]    _zz_dataOut_payload_0_7149;
  reg        [7:0]    _zz_dataOut_payload_0_7150;
  reg        [7:0]    _zz_dataOut_payload_0_7151;
  wire                _zz_dataOut_payload_0_7152;
  wire       [7:0]    _zz_dataOut_payload_0_7153;
  wire       [7:0]    _zz_dataOut_payload_0_7154;
  wire                _zz_dataOut_payload_0_7155;
  wire       [7:0]    _zz_dataOut_payload_0_7156;
  wire       [7:0]    _zz_dataOut_payload_0_7157;
  wire                _zz_dataOut_payload_0_7158;
  wire                _zz_dataOut_payload_0_7159;
  reg        [7:0]    _zz_dataOut_payload_0_7160;
  reg        [7:0]    _zz_dataOut_payload_0_7161;
  reg        [7:0]    _zz_dataOut_payload_0_7162;
  reg        [7:0]    _zz_dataOut_payload_0_7163;
  reg        [7:0]    _zz_dataOut_payload_0_7164;
  reg        [7:0]    _zz_dataOut_payload_0_7165;
  reg        [7:0]    _zz_dataOut_payload_0_7166;
  reg        [7:0]    _zz_dataOut_payload_0_7167;
  reg        [7:0]    _zz_dataOut_payload_0_7168;
  reg        [7:0]    _zz_dataOut_payload_0_7169;
  reg        [7:0]    _zz_dataOut_payload_0_7170;
  reg        [7:0]    _zz_dataOut_payload_0_7171;
  wire                _zz_dataOut_payload_0_7172;
  wire       [7:0]    _zz_dataOut_payload_0_7173;
  wire       [7:0]    _zz_dataOut_payload_0_7174;
  wire                _zz_dataOut_payload_0_7175;
  wire       [7:0]    _zz_dataOut_payload_0_7176;
  wire       [7:0]    _zz_dataOut_payload_0_7177;
  wire                _zz_dataOut_payload_0_7178;
  wire       [7:0]    _zz_dataOut_payload_0_7179;
  wire       [7:0]    _zz_dataOut_payload_0_7180;
  wire                _zz_dataOut_payload_0_7181;
  wire       [7:0]    _zz_dataOut_payload_0_7182;
  wire       [7:0]    _zz_dataOut_payload_0_7183;
  wire                _zz_dataOut_payload_0_7184;
  wire       [7:0]    _zz_dataOut_payload_0_7185;
  wire       [7:0]    _zz_dataOut_payload_0_7186;
  wire                _zz_dataOut_payload_0_7187;
  wire       [7:0]    _zz_dataOut_payload_0_7188;
  wire       [7:0]    _zz_dataOut_payload_0_7189;
  wire                _zz_dataOut_payload_0_7190;
  wire                _zz_dataOut_payload_0_7191;
  reg        [7:0]    _zz_dataOut_payload_0_7192;
  reg        [7:0]    _zz_dataOut_payload_0_7193;
  reg        [7:0]    _zz_dataOut_payload_0_7194;
  reg        [7:0]    _zz_dataOut_payload_0_7195;
  wire                _zz_dataOut_payload_0_7196;
  wire       [7:0]    _zz_dataOut_payload_0_7197;
  wire       [7:0]    _zz_dataOut_payload_0_7198;
  wire                _zz_dataOut_payload_0_7199;
  wire       [7:0]    _zz_dataOut_payload_0_7200;
  wire       [7:0]    _zz_dataOut_payload_0_7201;
  wire                _zz_dataOut_payload_0_7202;
  wire                _zz_dataOut_payload_0_7203;
  reg        [7:0]    _zz_dataOut_payload_0_7204;
  reg        [7:0]    _zz_dataOut_payload_0_7205;
  reg        [7:0]    _zz_dataOut_payload_0_7206;
  reg        [7:0]    _zz_dataOut_payload_0_7207;
  reg        [7:0]    _zz_dataOut_payload_0_7208;
  reg        [7:0]    _zz_dataOut_payload_0_7209;
  reg        [7:0]    _zz_dataOut_payload_0_7210;
  reg        [7:0]    _zz_dataOut_payload_0_7211;
  reg        [7:0]    _zz_dataOut_payload_0_7212;
  reg        [7:0]    _zz_dataOut_payload_0_7213;
  reg        [7:0]    _zz_dataOut_payload_0_7214;
  reg        [7:0]    _zz_dataOut_payload_0_7215;
  reg        [7:0]    _zz_dataOut_payload_0_7216;
  reg        [7:0]    _zz_dataOut_payload_0_7217;
  reg        [7:0]    _zz_dataOut_payload_0_7218;
  reg        [7:0]    _zz_dataOut_payload_0_7219;
  reg        [7:0]    _zz_dataOut_payload_0_7220;
  reg        [7:0]    _zz_dataOut_payload_0_7221;
  reg        [7:0]    _zz_dataOut_payload_0_7222;
  reg        [7:0]    _zz_dataOut_payload_0_7223;
  reg        [7:0]    _zz_dataOut_payload_0_7224;
  reg        [7:0]    _zz_dataOut_payload_0_7225;
  reg        [7:0]    _zz_dataOut_payload_0_7226;
  reg        [7:0]    _zz_dataOut_payload_0_7227;
  reg        [7:0]    _zz_dataOut_payload_0_7228;
  reg        [7:0]    _zz_dataOut_payload_0_7229;
  reg        [7:0]    _zz_dataOut_payload_0_7230;
  reg        [7:0]    _zz_dataOut_payload_0_7231;
  wire                _zz_dataOut_payload_0_7232;
  wire       [7:0]    _zz_dataOut_payload_0_7233;
  wire       [7:0]    _zz_dataOut_payload_0_7234;
  wire                _zz_dataOut_payload_0_7235;
  wire       [7:0]    _zz_dataOut_payload_0_7236;
  wire       [7:0]    _zz_dataOut_payload_0_7237;
  wire                _zz_dataOut_payload_0_7238;
  wire       [7:0]    _zz_dataOut_payload_0_7239;
  wire       [7:0]    _zz_dataOut_payload_0_7240;
  wire                _zz_dataOut_payload_0_7241;
  wire       [7:0]    _zz_dataOut_payload_0_7242;
  wire       [7:0]    _zz_dataOut_payload_0_7243;
  wire                _zz_dataOut_payload_0_7244;
  wire       [7:0]    _zz_dataOut_payload_0_7245;
  wire       [7:0]    _zz_dataOut_payload_0_7246;
  wire                _zz_dataOut_payload_0_7247;
  wire       [7:0]    _zz_dataOut_payload_0_7248;
  wire       [7:0]    _zz_dataOut_payload_0_7249;
  wire                _zz_dataOut_payload_0_7250;
  wire       [7:0]    _zz_dataOut_payload_0_7251;
  wire       [7:0]    _zz_dataOut_payload_0_7252;
  wire                _zz_dataOut_payload_0_7253;
  wire       [7:0]    _zz_dataOut_payload_0_7254;
  wire       [7:0]    _zz_dataOut_payload_0_7255;
  wire                _zz_dataOut_payload_0_7256;
  wire       [7:0]    _zz_dataOut_payload_0_7257;
  wire       [7:0]    _zz_dataOut_payload_0_7258;
  wire                _zz_dataOut_payload_0_7259;
  wire       [7:0]    _zz_dataOut_payload_0_7260;
  wire       [7:0]    _zz_dataOut_payload_0_7261;
  wire                _zz_dataOut_payload_0_7262;
  wire       [7:0]    _zz_dataOut_payload_0_7263;
  wire       [7:0]    _zz_dataOut_payload_0_7264;
  wire                _zz_dataOut_payload_0_7265;
  wire       [7:0]    _zz_dataOut_payload_0_7266;
  wire       [7:0]    _zz_dataOut_payload_0_7267;
  wire                _zz_dataOut_payload_0_7268;
  wire       [7:0]    _zz_dataOut_payload_0_7269;
  wire       [7:0]    _zz_dataOut_payload_0_7270;
  wire                _zz_dataOut_payload_0_7271;
  wire       [7:0]    _zz_dataOut_payload_0_7272;
  wire       [7:0]    _zz_dataOut_payload_0_7273;
  wire                _zz_dataOut_payload_0_7274;
  wire                _zz_dataOut_payload_0_7275;
  reg        [7:0]    _zz_dataOut_payload_0_7276;
  reg        [7:0]    _zz_dataOut_payload_0_7277;
  reg        [7:0]    _zz_dataOut_payload_0_7278;
  reg        [7:0]    _zz_dataOut_payload_0_7279;
  wire                _zz_dataOut_payload_0_7280;
  wire       [7:0]    _zz_dataOut_payload_0_7281;
  wire       [7:0]    _zz_dataOut_payload_0_7282;
  wire                _zz_dataOut_payload_0_7283;
  wire       [7:0]    _zz_dataOut_payload_0_7284;
  wire       [7:0]    _zz_dataOut_payload_0_7285;
  wire                _zz_dataOut_payload_0_7286;
  wire                _zz_dataOut_payload_0_7287;
  reg        [7:0]    _zz_dataOut_payload_0_7288;
  reg        [7:0]    _zz_dataOut_payload_0_7289;
  reg        [7:0]    _zz_dataOut_payload_0_7290;
  reg        [7:0]    _zz_dataOut_payload_0_7291;
  reg        [7:0]    _zz_dataOut_payload_0_7292;
  reg        [7:0]    _zz_dataOut_payload_0_7293;
  reg        [7:0]    _zz_dataOut_payload_0_7294;
  reg        [7:0]    _zz_dataOut_payload_0_7295;
  reg        [7:0]    _zz_dataOut_payload_0_7296;
  reg        [7:0]    _zz_dataOut_payload_0_7297;
  reg        [7:0]    _zz_dataOut_payload_0_7298;
  reg        [7:0]    _zz_dataOut_payload_0_7299;
  wire                _zz_dataOut_payload_0_7300;
  wire       [7:0]    _zz_dataOut_payload_0_7301;
  wire       [7:0]    _zz_dataOut_payload_0_7302;
  wire                _zz_dataOut_payload_0_7303;
  wire       [7:0]    _zz_dataOut_payload_0_7304;
  wire       [7:0]    _zz_dataOut_payload_0_7305;
  wire                _zz_dataOut_payload_0_7306;
  wire       [7:0]    _zz_dataOut_payload_0_7307;
  wire       [7:0]    _zz_dataOut_payload_0_7308;
  wire                _zz_dataOut_payload_0_7309;
  wire       [7:0]    _zz_dataOut_payload_0_7310;
  wire       [7:0]    _zz_dataOut_payload_0_7311;
  wire                _zz_dataOut_payload_0_7312;
  wire       [7:0]    _zz_dataOut_payload_0_7313;
  wire       [7:0]    _zz_dataOut_payload_0_7314;
  wire                _zz_dataOut_payload_0_7315;
  wire       [7:0]    _zz_dataOut_payload_0_7316;
  wire       [7:0]    _zz_dataOut_payload_0_7317;
  wire                _zz_dataOut_payload_0_7318;
  wire                _zz_dataOut_payload_0_7319;
  reg        [7:0]    _zz_dataOut_payload_0_7320;
  reg        [7:0]    _zz_dataOut_payload_0_7321;
  reg        [7:0]    _zz_dataOut_payload_0_7322;
  reg        [7:0]    _zz_dataOut_payload_0_7323;
  wire                _zz_dataOut_payload_0_7324;
  wire       [7:0]    _zz_dataOut_payload_0_7325;
  wire       [7:0]    _zz_dataOut_payload_0_7326;
  wire                _zz_dataOut_payload_0_7327;
  wire       [7:0]    _zz_dataOut_payload_0_7328;
  wire       [7:0]    _zz_dataOut_payload_0_7329;
  wire                _zz_dataOut_payload_0_7330;
  wire                _zz_dataOut_payload_0_7331;
  reg        [7:0]    _zz_dataOut_payload_0_7332;
  reg        [7:0]    _zz_dataOut_payload_0_7333;
  reg        [7:0]    _zz_dataOut_payload_0_7334;
  reg        [7:0]    _zz_dataOut_payload_0_7335;
  reg        [7:0]    _zz_dataOut_payload_0_7336;
  reg        [7:0]    _zz_dataOut_payload_0_7337;
  reg        [7:0]    _zz_dataOut_payload_0_7338;
  reg        [7:0]    _zz_dataOut_payload_0_7339;
  reg        [7:0]    _zz_dataOut_payload_0_7340;
  reg        [7:0]    _zz_dataOut_payload_0_7341;
  reg        [7:0]    _zz_dataOut_payload_0_7342;
  reg        [7:0]    _zz_dataOut_payload_0_7343;
  reg        [7:0]    _zz_dataOut_payload_0_7344;
  reg        [7:0]    _zz_dataOut_payload_0_7345;
  reg        [7:0]    _zz_dataOut_payload_0_7346;
  reg        [7:0]    _zz_dataOut_payload_0_7347;
  reg        [7:0]    _zz_dataOut_payload_0_7348;
  reg        [7:0]    _zz_dataOut_payload_0_7349;
  reg        [7:0]    _zz_dataOut_payload_0_7350;
  reg        [7:0]    _zz_dataOut_payload_0_7351;
  reg        [7:0]    _zz_dataOut_payload_0_7352;
  reg        [7:0]    _zz_dataOut_payload_0_7353;
  reg        [7:0]    _zz_dataOut_payload_0_7354;
  reg        [7:0]    _zz_dataOut_payload_0_7355;
  reg        [7:0]    _zz_dataOut_payload_0_7356;
  reg        [7:0]    _zz_dataOut_payload_0_7357;
  reg        [7:0]    _zz_dataOut_payload_0_7358;
  reg        [7:0]    _zz_dataOut_payload_0_7359;
  reg        [7:0]    _zz_dataOut_payload_0_7360;
  reg        [7:0]    _zz_dataOut_payload_0_7361;
  reg        [7:0]    _zz_dataOut_payload_0_7362;
  reg        [7:0]    _zz_dataOut_payload_0_7363;
  reg        [7:0]    _zz_dataOut_payload_0_7364;
  reg        [7:0]    _zz_dataOut_payload_0_7365;
  reg        [7:0]    _zz_dataOut_payload_0_7366;
  reg        [7:0]    _zz_dataOut_payload_0_7367;
  reg        [7:0]    _zz_dataOut_payload_0_7368;
  reg        [7:0]    _zz_dataOut_payload_0_7369;
  reg        [7:0]    _zz_dataOut_payload_0_7370;
  reg        [7:0]    _zz_dataOut_payload_0_7371;
  reg        [7:0]    _zz_dataOut_payload_0_7372;
  reg        [7:0]    _zz_dataOut_payload_0_7373;
  reg        [7:0]    _zz_dataOut_payload_0_7374;
  reg        [7:0]    _zz_dataOut_payload_0_7375;
  reg        [7:0]    _zz_dataOut_payload_0_7376;
  reg        [7:0]    _zz_dataOut_payload_0_7377;
  reg        [7:0]    _zz_dataOut_payload_0_7378;
  reg        [7:0]    _zz_dataOut_payload_0_7379;
  reg        [7:0]    _zz_dataOut_payload_0_7380;
  reg        [7:0]    _zz_dataOut_payload_0_7381;
  reg        [7:0]    _zz_dataOut_payload_0_7382;
  reg        [7:0]    _zz_dataOut_payload_0_7383;
  reg        [7:0]    _zz_dataOut_payload_0_7384;
  reg        [7:0]    _zz_dataOut_payload_0_7385;
  reg        [7:0]    _zz_dataOut_payload_0_7386;
  reg        [7:0]    _zz_dataOut_payload_0_7387;
  reg        [7:0]    _zz_dataOut_payload_0_7388;
  reg        [7:0]    _zz_dataOut_payload_0_7389;
  reg        [7:0]    _zz_dataOut_payload_0_7390;
  reg        [7:0]    _zz_dataOut_payload_0_7391;
  wire                _zz_dataOut_payload_0_7392;
  wire       [7:0]    _zz_dataOut_payload_0_7393;
  wire       [7:0]    _zz_dataOut_payload_0_7394;
  wire                _zz_dataOut_payload_0_7395;
  wire       [7:0]    _zz_dataOut_payload_0_7396;
  wire       [7:0]    _zz_dataOut_payload_0_7397;
  wire                _zz_dataOut_payload_0_7398;
  wire       [7:0]    _zz_dataOut_payload_0_7399;
  wire       [7:0]    _zz_dataOut_payload_0_7400;
  wire                _zz_dataOut_payload_0_7401;
  wire       [7:0]    _zz_dataOut_payload_0_7402;
  wire       [7:0]    _zz_dataOut_payload_0_7403;
  wire                _zz_dataOut_payload_0_7404;
  wire       [7:0]    _zz_dataOut_payload_0_7405;
  wire       [7:0]    _zz_dataOut_payload_0_7406;
  wire                _zz_dataOut_payload_0_7407;
  wire       [7:0]    _zz_dataOut_payload_0_7408;
  wire       [7:0]    _zz_dataOut_payload_0_7409;
  wire                _zz_dataOut_payload_0_7410;
  wire       [7:0]    _zz_dataOut_payload_0_7411;
  wire       [7:0]    _zz_dataOut_payload_0_7412;
  wire                _zz_dataOut_payload_0_7413;
  wire       [7:0]    _zz_dataOut_payload_0_7414;
  wire       [7:0]    _zz_dataOut_payload_0_7415;
  wire                _zz_dataOut_payload_0_7416;
  wire       [7:0]    _zz_dataOut_payload_0_7417;
  wire       [7:0]    _zz_dataOut_payload_0_7418;
  wire                _zz_dataOut_payload_0_7419;
  wire       [7:0]    _zz_dataOut_payload_0_7420;
  wire       [7:0]    _zz_dataOut_payload_0_7421;
  wire                _zz_dataOut_payload_0_7422;
  wire       [7:0]    _zz_dataOut_payload_0_7423;
  wire       [7:0]    _zz_dataOut_payload_0_7424;
  wire                _zz_dataOut_payload_0_7425;
  wire       [7:0]    _zz_dataOut_payload_0_7426;
  wire       [7:0]    _zz_dataOut_payload_0_7427;
  wire                _zz_dataOut_payload_0_7428;
  wire       [7:0]    _zz_dataOut_payload_0_7429;
  wire       [7:0]    _zz_dataOut_payload_0_7430;
  wire                _zz_dataOut_payload_0_7431;
  wire       [7:0]    _zz_dataOut_payload_0_7432;
  wire       [7:0]    _zz_dataOut_payload_0_7433;
  wire                _zz_dataOut_payload_0_7434;
  wire       [7:0]    _zz_dataOut_payload_0_7435;
  wire       [7:0]    _zz_dataOut_payload_0_7436;
  wire                _zz_dataOut_payload_0_7437;
  wire       [7:0]    _zz_dataOut_payload_0_7438;
  wire       [7:0]    _zz_dataOut_payload_0_7439;
  wire                _zz_dataOut_payload_0_7440;
  wire       [7:0]    _zz_dataOut_payload_0_7441;
  wire       [7:0]    _zz_dataOut_payload_0_7442;
  wire                _zz_dataOut_payload_0_7443;
  wire       [7:0]    _zz_dataOut_payload_0_7444;
  wire       [7:0]    _zz_dataOut_payload_0_7445;
  wire                _zz_dataOut_payload_0_7446;
  wire       [7:0]    _zz_dataOut_payload_0_7447;
  wire       [7:0]    _zz_dataOut_payload_0_7448;
  wire                _zz_dataOut_payload_0_7449;
  wire       [7:0]    _zz_dataOut_payload_0_7450;
  wire       [7:0]    _zz_dataOut_payload_0_7451;
  wire                _zz_dataOut_payload_0_7452;
  wire       [7:0]    _zz_dataOut_payload_0_7453;
  wire       [7:0]    _zz_dataOut_payload_0_7454;
  wire                _zz_dataOut_payload_0_7455;
  wire       [7:0]    _zz_dataOut_payload_0_7456;
  wire       [7:0]    _zz_dataOut_payload_0_7457;
  wire                _zz_dataOut_payload_0_7458;
  wire       [7:0]    _zz_dataOut_payload_0_7459;
  wire       [7:0]    _zz_dataOut_payload_0_7460;
  wire                _zz_dataOut_payload_0_7461;
  wire       [7:0]    _zz_dataOut_payload_0_7462;
  wire       [7:0]    _zz_dataOut_payload_0_7463;
  wire                _zz_dataOut_payload_0_7464;
  wire       [7:0]    _zz_dataOut_payload_0_7465;
  wire       [7:0]    _zz_dataOut_payload_0_7466;
  wire                _zz_dataOut_payload_0_7467;
  wire       [7:0]    _zz_dataOut_payload_0_7468;
  wire       [7:0]    _zz_dataOut_payload_0_7469;
  wire                _zz_dataOut_payload_0_7470;
  wire       [7:0]    _zz_dataOut_payload_0_7471;
  wire       [7:0]    _zz_dataOut_payload_0_7472;
  wire                _zz_dataOut_payload_0_7473;
  wire       [7:0]    _zz_dataOut_payload_0_7474;
  wire       [7:0]    _zz_dataOut_payload_0_7475;
  wire                _zz_dataOut_payload_0_7476;
  wire       [7:0]    _zz_dataOut_payload_0_7477;
  wire       [7:0]    _zz_dataOut_payload_0_7478;
  wire                _zz_dataOut_payload_0_7479;
  wire       [7:0]    _zz_dataOut_payload_0_7480;
  wire       [7:0]    _zz_dataOut_payload_0_7481;
  wire                _zz_dataOut_payload_0_7482;
  wire                _zz_dataOut_payload_0_7483;
  reg        [7:0]    _zz_dataOut_payload_0_7484;
  reg        [7:0]    _zz_dataOut_payload_0_7485;
  reg        [7:0]    _zz_dataOut_payload_0_7486;
  reg        [7:0]    _zz_dataOut_payload_0_7487;
  wire                _zz_dataOut_payload_0_7488;
  wire       [7:0]    _zz_dataOut_payload_0_7489;
  wire       [7:0]    _zz_dataOut_payload_0_7490;
  wire                _zz_dataOut_payload_0_7491;
  wire       [7:0]    _zz_dataOut_payload_0_7492;
  wire       [7:0]    _zz_dataOut_payload_0_7493;
  wire                _zz_dataOut_payload_0_7494;
  wire                _zz_dataOut_payload_0_7495;
  reg        [7:0]    _zz_dataOut_payload_0_7496;
  reg        [7:0]    _zz_dataOut_payload_0_7497;
  reg        [7:0]    _zz_dataOut_payload_0_7498;
  reg        [7:0]    _zz_dataOut_payload_0_7499;
  reg        [7:0]    _zz_dataOut_payload_0_7500;
  reg        [7:0]    _zz_dataOut_payload_0_7501;
  reg        [7:0]    _zz_dataOut_payload_0_7502;
  reg        [7:0]    _zz_dataOut_payload_0_7503;
  reg        [7:0]    _zz_dataOut_payload_0_7504;
  reg        [7:0]    _zz_dataOut_payload_0_7505;
  reg        [7:0]    _zz_dataOut_payload_0_7506;
  reg        [7:0]    _zz_dataOut_payload_0_7507;
  wire                _zz_dataOut_payload_0_7508;
  wire       [7:0]    _zz_dataOut_payload_0_7509;
  wire       [7:0]    _zz_dataOut_payload_0_7510;
  wire                _zz_dataOut_payload_0_7511;
  wire       [7:0]    _zz_dataOut_payload_0_7512;
  wire       [7:0]    _zz_dataOut_payload_0_7513;
  wire                _zz_dataOut_payload_0_7514;
  wire       [7:0]    _zz_dataOut_payload_0_7515;
  wire       [7:0]    _zz_dataOut_payload_0_7516;
  wire                _zz_dataOut_payload_0_7517;
  wire       [7:0]    _zz_dataOut_payload_0_7518;
  wire       [7:0]    _zz_dataOut_payload_0_7519;
  wire                _zz_dataOut_payload_0_7520;
  wire       [7:0]    _zz_dataOut_payload_0_7521;
  wire       [7:0]    _zz_dataOut_payload_0_7522;
  wire                _zz_dataOut_payload_0_7523;
  wire       [7:0]    _zz_dataOut_payload_0_7524;
  wire       [7:0]    _zz_dataOut_payload_0_7525;
  wire                _zz_dataOut_payload_0_7526;
  wire                _zz_dataOut_payload_0_7527;
  reg        [7:0]    _zz_dataOut_payload_0_7528;
  reg        [7:0]    _zz_dataOut_payload_0_7529;
  reg        [7:0]    _zz_dataOut_payload_0_7530;
  reg        [7:0]    _zz_dataOut_payload_0_7531;
  wire                _zz_dataOut_payload_0_7532;
  wire       [7:0]    _zz_dataOut_payload_0_7533;
  wire       [7:0]    _zz_dataOut_payload_0_7534;
  wire                _zz_dataOut_payload_0_7535;
  wire       [7:0]    _zz_dataOut_payload_0_7536;
  wire       [7:0]    _zz_dataOut_payload_0_7537;
  wire                _zz_dataOut_payload_0_7538;
  wire                _zz_dataOut_payload_0_7539;
  reg        [7:0]    _zz_dataOut_payload_0_7540;
  reg        [7:0]    _zz_dataOut_payload_0_7541;
  reg        [7:0]    _zz_dataOut_payload_0_7542;
  reg        [7:0]    _zz_dataOut_payload_0_7543;
  reg        [7:0]    _zz_dataOut_payload_0_7544;
  reg        [7:0]    _zz_dataOut_payload_0_7545;
  reg        [7:0]    _zz_dataOut_payload_0_7546;
  reg        [7:0]    _zz_dataOut_payload_0_7547;
  reg        [7:0]    _zz_dataOut_payload_0_7548;
  reg        [7:0]    _zz_dataOut_payload_0_7549;
  reg        [7:0]    _zz_dataOut_payload_0_7550;
  reg        [7:0]    _zz_dataOut_payload_0_7551;
  reg        [7:0]    _zz_dataOut_payload_0_7552;
  reg        [7:0]    _zz_dataOut_payload_0_7553;
  reg        [7:0]    _zz_dataOut_payload_0_7554;
  reg        [7:0]    _zz_dataOut_payload_0_7555;
  reg        [7:0]    _zz_dataOut_payload_0_7556;
  reg        [7:0]    _zz_dataOut_payload_0_7557;
  reg        [7:0]    _zz_dataOut_payload_0_7558;
  reg        [7:0]    _zz_dataOut_payload_0_7559;
  reg        [7:0]    _zz_dataOut_payload_0_7560;
  reg        [7:0]    _zz_dataOut_payload_0_7561;
  reg        [7:0]    _zz_dataOut_payload_0_7562;
  reg        [7:0]    _zz_dataOut_payload_0_7563;
  reg        [7:0]    _zz_dataOut_payload_0_7564;
  reg        [7:0]    _zz_dataOut_payload_0_7565;
  reg        [7:0]    _zz_dataOut_payload_0_7566;
  reg        [7:0]    _zz_dataOut_payload_0_7567;
  wire                _zz_dataOut_payload_0_7568;
  wire       [7:0]    _zz_dataOut_payload_0_7569;
  wire       [7:0]    _zz_dataOut_payload_0_7570;
  wire                _zz_dataOut_payload_0_7571;
  wire       [7:0]    _zz_dataOut_payload_0_7572;
  wire       [7:0]    _zz_dataOut_payload_0_7573;
  wire                _zz_dataOut_payload_0_7574;
  wire       [7:0]    _zz_dataOut_payload_0_7575;
  wire       [7:0]    _zz_dataOut_payload_0_7576;
  wire                _zz_dataOut_payload_0_7577;
  wire       [7:0]    _zz_dataOut_payload_0_7578;
  wire       [7:0]    _zz_dataOut_payload_0_7579;
  wire                _zz_dataOut_payload_0_7580;
  wire       [7:0]    _zz_dataOut_payload_0_7581;
  wire       [7:0]    _zz_dataOut_payload_0_7582;
  wire                _zz_dataOut_payload_0_7583;
  wire       [7:0]    _zz_dataOut_payload_0_7584;
  wire       [7:0]    _zz_dataOut_payload_0_7585;
  wire                _zz_dataOut_payload_0_7586;
  wire       [7:0]    _zz_dataOut_payload_0_7587;
  wire       [7:0]    _zz_dataOut_payload_0_7588;
  wire                _zz_dataOut_payload_0_7589;
  wire       [7:0]    _zz_dataOut_payload_0_7590;
  wire       [7:0]    _zz_dataOut_payload_0_7591;
  wire                _zz_dataOut_payload_0_7592;
  wire       [7:0]    _zz_dataOut_payload_0_7593;
  wire       [7:0]    _zz_dataOut_payload_0_7594;
  wire                _zz_dataOut_payload_0_7595;
  wire       [7:0]    _zz_dataOut_payload_0_7596;
  wire       [7:0]    _zz_dataOut_payload_0_7597;
  wire                _zz_dataOut_payload_0_7598;
  wire       [7:0]    _zz_dataOut_payload_0_7599;
  wire       [7:0]    _zz_dataOut_payload_0_7600;
  wire                _zz_dataOut_payload_0_7601;
  wire       [7:0]    _zz_dataOut_payload_0_7602;
  wire       [7:0]    _zz_dataOut_payload_0_7603;
  wire                _zz_dataOut_payload_0_7604;
  wire       [7:0]    _zz_dataOut_payload_0_7605;
  wire       [7:0]    _zz_dataOut_payload_0_7606;
  wire                _zz_dataOut_payload_0_7607;
  wire       [7:0]    _zz_dataOut_payload_0_7608;
  wire       [7:0]    _zz_dataOut_payload_0_7609;
  wire                _zz_dataOut_payload_0_7610;
  wire                _zz_dataOut_payload_0_7611;
  reg        [7:0]    _zz_dataOut_payload_0_7612;
  reg        [7:0]    _zz_dataOut_payload_0_7613;
  reg        [7:0]    _zz_dataOut_payload_0_7614;
  reg        [7:0]    _zz_dataOut_payload_0_7615;
  wire                _zz_dataOut_payload_0_7616;
  wire       [7:0]    _zz_dataOut_payload_0_7617;
  wire       [7:0]    _zz_dataOut_payload_0_7618;
  wire                _zz_dataOut_payload_0_7619;
  wire       [7:0]    _zz_dataOut_payload_0_7620;
  wire       [7:0]    _zz_dataOut_payload_0_7621;
  wire                _zz_dataOut_payload_0_7622;
  wire                _zz_dataOut_payload_0_7623;
  reg        [7:0]    _zz_dataOut_payload_0_7624;
  reg        [7:0]    _zz_dataOut_payload_0_7625;
  reg        [7:0]    _zz_dataOut_payload_0_7626;
  reg        [7:0]    _zz_dataOut_payload_0_7627;
  reg        [7:0]    _zz_dataOut_payload_0_7628;
  reg        [7:0]    _zz_dataOut_payload_0_7629;
  reg        [7:0]    _zz_dataOut_payload_0_7630;
  reg        [7:0]    _zz_dataOut_payload_0_7631;
  reg        [7:0]    _zz_dataOut_payload_0_7632;
  reg        [7:0]    _zz_dataOut_payload_0_7633;
  reg        [7:0]    _zz_dataOut_payload_0_7634;
  reg        [7:0]    _zz_dataOut_payload_0_7635;
  wire                _zz_dataOut_payload_0_7636;
  wire       [7:0]    _zz_dataOut_payload_0_7637;
  wire       [7:0]    _zz_dataOut_payload_0_7638;
  wire                _zz_dataOut_payload_0_7639;
  wire       [7:0]    _zz_dataOut_payload_0_7640;
  wire       [7:0]    _zz_dataOut_payload_0_7641;
  wire                _zz_dataOut_payload_0_7642;
  wire       [7:0]    _zz_dataOut_payload_0_7643;
  wire       [7:0]    _zz_dataOut_payload_0_7644;
  wire                _zz_dataOut_payload_0_7645;
  wire       [7:0]    _zz_dataOut_payload_0_7646;
  wire       [7:0]    _zz_dataOut_payload_0_7647;
  wire                _zz_dataOut_payload_0_7648;
  wire       [7:0]    _zz_dataOut_payload_0_7649;
  wire       [7:0]    _zz_dataOut_payload_0_7650;
  wire                _zz_dataOut_payload_0_7651;
  wire       [7:0]    _zz_dataOut_payload_0_7652;
  wire       [7:0]    _zz_dataOut_payload_0_7653;
  wire                _zz_dataOut_payload_0_7654;
  wire                _zz_dataOut_payload_0_7655;
  reg        [7:0]    _zz_dataOut_payload_0_7656;
  reg        [7:0]    _zz_dataOut_payload_0_7657;
  reg        [7:0]    _zz_dataOut_payload_0_7658;
  reg        [7:0]    _zz_dataOut_payload_0_7659;
  wire                _zz_dataOut_payload_0_7660;
  wire       [7:0]    _zz_dataOut_payload_0_7661;
  wire       [7:0]    _zz_dataOut_payload_0_7662;
  wire                _zz_dataOut_payload_0_7663;
  wire       [7:0]    _zz_dataOut_payload_0_7664;
  wire       [7:0]    _zz_dataOut_payload_0_7665;
  wire                _zz_dataOut_payload_0_7666;
  wire                _zz_dataOut_payload_0_7667;
  reg        [7:0]    _zz_dataOut_payload_0_7668;
  reg        [7:0]    _zz_dataOut_payload_0_7669;
  reg        [7:0]    _zz_dataOut_payload_0_7670;
  reg        [7:0]    _zz_dataOut_payload_0_7671;
  reg        [7:0]    _zz_dataOut_payload_0_7672;
  reg        [7:0]    _zz_dataOut_payload_0_7673;
  reg        [7:0]    _zz_dataOut_payload_0_7674;
  reg        [7:0]    _zz_dataOut_payload_0_7675;
  reg        [7:0]    _zz_dataOut_payload_0_7676;
  reg        [7:0]    _zz_dataOut_payload_0_7677;
  reg        [7:0]    _zz_dataOut_payload_0_7678;
  reg        [7:0]    _zz_dataOut_payload_0_7679;
  reg        [7:0]    _zz_dataOut_payload_0_7680;
  reg        [7:0]    _zz_dataOut_payload_0_7681;
  reg        [7:0]    _zz_dataOut_payload_0_7682;
  reg        [7:0]    _zz_dataOut_payload_0_7683;
  reg        [7:0]    _zz_dataOut_payload_0_7684;
  reg        [7:0]    _zz_dataOut_payload_0_7685;
  reg        [7:0]    _zz_dataOut_payload_0_7686;
  reg        [7:0]    _zz_dataOut_payload_0_7687;
  reg        [7:0]    _zz_dataOut_payload_0_7688;
  reg        [7:0]    _zz_dataOut_payload_0_7689;
  reg        [7:0]    _zz_dataOut_payload_0_7690;
  reg        [7:0]    _zz_dataOut_payload_0_7691;
  reg        [7:0]    _zz_dataOut_payload_0_7692;
  reg        [7:0]    _zz_dataOut_payload_0_7693;
  reg        [7:0]    _zz_dataOut_payload_0_7694;
  reg        [7:0]    _zz_dataOut_payload_0_7695;
  reg        [7:0]    _zz_dataOut_payload_0_7696;
  reg        [7:0]    _zz_dataOut_payload_0_7697;
  reg        [7:0]    _zz_dataOut_payload_0_7698;
  reg        [7:0]    _zz_dataOut_payload_0_7699;
  reg        [7:0]    _zz_dataOut_payload_0_7700;
  reg        [7:0]    _zz_dataOut_payload_0_7701;
  reg        [7:0]    _zz_dataOut_payload_0_7702;
  reg        [7:0]    _zz_dataOut_payload_0_7703;
  reg        [7:0]    _zz_dataOut_payload_0_7704;
  reg        [7:0]    _zz_dataOut_payload_0_7705;
  reg        [7:0]    _zz_dataOut_payload_0_7706;
  reg        [7:0]    _zz_dataOut_payload_0_7707;
  reg        [7:0]    _zz_dataOut_payload_0_7708;
  reg        [7:0]    _zz_dataOut_payload_0_7709;
  reg        [7:0]    _zz_dataOut_payload_0_7710;
  reg        [7:0]    _zz_dataOut_payload_0_7711;
  reg        [7:0]    _zz_dataOut_payload_0_7712;
  reg        [7:0]    _zz_dataOut_payload_0_7713;
  reg        [7:0]    _zz_dataOut_payload_0_7714;
  reg        [7:0]    _zz_dataOut_payload_0_7715;
  reg        [7:0]    _zz_dataOut_payload_0_7716;
  reg        [7:0]    _zz_dataOut_payload_0_7717;
  reg        [7:0]    _zz_dataOut_payload_0_7718;
  reg        [7:0]    _zz_dataOut_payload_0_7719;
  reg        [7:0]    _zz_dataOut_payload_0_7720;
  reg        [7:0]    _zz_dataOut_payload_0_7721;
  reg        [7:0]    _zz_dataOut_payload_0_7722;
  reg        [7:0]    _zz_dataOut_payload_0_7723;
  reg        [7:0]    _zz_dataOut_payload_0_7724;
  reg        [7:0]    _zz_dataOut_payload_0_7725;
  reg        [7:0]    _zz_dataOut_payload_0_7726;
  reg        [7:0]    _zz_dataOut_payload_0_7727;
  wire                _zz_dataOut_payload_0_7728;
  wire       [7:0]    _zz_dataOut_payload_0_7729;
  wire       [7:0]    _zz_dataOut_payload_0_7730;
  wire                _zz_dataOut_payload_0_7731;
  wire       [7:0]    _zz_dataOut_payload_0_7732;
  wire       [7:0]    _zz_dataOut_payload_0_7733;
  wire                _zz_dataOut_payload_0_7734;
  wire       [7:0]    _zz_dataOut_payload_0_7735;
  wire       [7:0]    _zz_dataOut_payload_0_7736;
  wire                _zz_dataOut_payload_0_7737;
  wire       [7:0]    _zz_dataOut_payload_0_7738;
  wire       [7:0]    _zz_dataOut_payload_0_7739;
  wire                _zz_dataOut_payload_0_7740;
  wire       [7:0]    _zz_dataOut_payload_0_7741;
  wire       [7:0]    _zz_dataOut_payload_0_7742;
  wire                _zz_dataOut_payload_0_7743;
  wire       [7:0]    _zz_dataOut_payload_0_7744;
  wire       [7:0]    _zz_dataOut_payload_0_7745;
  wire                _zz_dataOut_payload_0_7746;
  wire       [7:0]    _zz_dataOut_payload_0_7747;
  wire       [7:0]    _zz_dataOut_payload_0_7748;
  wire                _zz_dataOut_payload_0_7749;
  wire       [7:0]    _zz_dataOut_payload_0_7750;
  wire       [7:0]    _zz_dataOut_payload_0_7751;
  wire                _zz_dataOut_payload_0_7752;
  wire       [7:0]    _zz_dataOut_payload_0_7753;
  wire       [7:0]    _zz_dataOut_payload_0_7754;
  wire                _zz_dataOut_payload_0_7755;
  wire       [7:0]    _zz_dataOut_payload_0_7756;
  wire       [7:0]    _zz_dataOut_payload_0_7757;
  wire                _zz_dataOut_payload_0_7758;
  wire       [7:0]    _zz_dataOut_payload_0_7759;
  wire       [7:0]    _zz_dataOut_payload_0_7760;
  wire                _zz_dataOut_payload_0_7761;
  wire       [7:0]    _zz_dataOut_payload_0_7762;
  wire       [7:0]    _zz_dataOut_payload_0_7763;
  wire                _zz_dataOut_payload_0_7764;
  wire       [7:0]    _zz_dataOut_payload_0_7765;
  wire       [7:0]    _zz_dataOut_payload_0_7766;
  wire                _zz_dataOut_payload_0_7767;
  wire       [7:0]    _zz_dataOut_payload_0_7768;
  wire       [7:0]    _zz_dataOut_payload_0_7769;
  wire                _zz_dataOut_payload_0_7770;
  wire       [7:0]    _zz_dataOut_payload_0_7771;
  wire       [7:0]    _zz_dataOut_payload_0_7772;
  wire                _zz_dataOut_payload_0_7773;
  wire       [7:0]    _zz_dataOut_payload_0_7774;
  wire       [7:0]    _zz_dataOut_payload_0_7775;
  wire                _zz_dataOut_payload_0_7776;
  wire       [7:0]    _zz_dataOut_payload_0_7777;
  wire       [7:0]    _zz_dataOut_payload_0_7778;
  wire                _zz_dataOut_payload_0_7779;
  wire       [7:0]    _zz_dataOut_payload_0_7780;
  wire       [7:0]    _zz_dataOut_payload_0_7781;
  wire                _zz_dataOut_payload_0_7782;
  wire       [7:0]    _zz_dataOut_payload_0_7783;
  wire       [7:0]    _zz_dataOut_payload_0_7784;
  wire                _zz_dataOut_payload_0_7785;
  wire       [7:0]    _zz_dataOut_payload_0_7786;
  wire       [7:0]    _zz_dataOut_payload_0_7787;
  wire                _zz_dataOut_payload_0_7788;
  wire       [7:0]    _zz_dataOut_payload_0_7789;
  wire       [7:0]    _zz_dataOut_payload_0_7790;
  wire                _zz_dataOut_payload_0_7791;
  wire       [7:0]    _zz_dataOut_payload_0_7792;
  wire       [7:0]    _zz_dataOut_payload_0_7793;
  wire                _zz_dataOut_payload_0_7794;
  wire       [7:0]    _zz_dataOut_payload_0_7795;
  wire       [7:0]    _zz_dataOut_payload_0_7796;
  wire                _zz_dataOut_payload_0_7797;
  wire       [7:0]    _zz_dataOut_payload_0_7798;
  wire       [7:0]    _zz_dataOut_payload_0_7799;
  wire                _zz_dataOut_payload_0_7800;
  wire       [7:0]    _zz_dataOut_payload_0_7801;
  wire       [7:0]    _zz_dataOut_payload_0_7802;
  wire                _zz_dataOut_payload_0_7803;
  wire       [7:0]    _zz_dataOut_payload_0_7804;
  wire       [7:0]    _zz_dataOut_payload_0_7805;
  wire                _zz_dataOut_payload_0_7806;
  wire       [7:0]    _zz_dataOut_payload_0_7807;
  wire       [7:0]    _zz_dataOut_payload_0_7808;
  wire                _zz_dataOut_payload_0_7809;
  wire       [7:0]    _zz_dataOut_payload_0_7810;
  wire       [7:0]    _zz_dataOut_payload_0_7811;
  wire                _zz_dataOut_payload_0_7812;
  wire       [7:0]    _zz_dataOut_payload_0_7813;
  wire       [7:0]    _zz_dataOut_payload_0_7814;
  wire                _zz_dataOut_payload_0_7815;
  wire       [7:0]    _zz_dataOut_payload_0_7816;
  wire       [7:0]    _zz_dataOut_payload_0_7817;
  wire                _zz_dataOut_payload_0_7818;
  wire                _zz_dataOut_payload_0_7819;
  reg        [7:0]    _zz_dataOut_payload_0_7820;
  reg        [7:0]    _zz_dataOut_payload_0_7821;
  reg        [7:0]    _zz_dataOut_payload_0_7822;
  reg        [7:0]    _zz_dataOut_payload_0_7823;
  wire                _zz_dataOut_payload_0_7824;
  wire       [7:0]    _zz_dataOut_payload_0_7825;
  wire       [7:0]    _zz_dataOut_payload_0_7826;
  wire                _zz_dataOut_payload_0_7827;
  wire       [7:0]    _zz_dataOut_payload_0_7828;
  wire       [7:0]    _zz_dataOut_payload_0_7829;
  wire                _zz_dataOut_payload_0_7830;
  wire                _zz_dataOut_payload_0_7831;
  reg        [7:0]    _zz_dataOut_payload_0_7832;
  reg        [7:0]    _zz_dataOut_payload_0_7833;
  reg        [7:0]    _zz_dataOut_payload_0_7834;
  reg        [7:0]    _zz_dataOut_payload_0_7835;
  reg        [7:0]    _zz_dataOut_payload_0_7836;
  reg        [7:0]    _zz_dataOut_payload_0_7837;
  reg        [7:0]    _zz_dataOut_payload_0_7838;
  reg        [7:0]    _zz_dataOut_payload_0_7839;
  reg        [7:0]    _zz_dataOut_payload_0_7840;
  reg        [7:0]    _zz_dataOut_payload_0_7841;
  reg        [7:0]    _zz_dataOut_payload_0_7842;
  reg        [7:0]    _zz_dataOut_payload_0_7843;
  wire                _zz_dataOut_payload_0_7844;
  wire       [7:0]    _zz_dataOut_payload_0_7845;
  wire       [7:0]    _zz_dataOut_payload_0_7846;
  wire                _zz_dataOut_payload_0_7847;
  wire       [7:0]    _zz_dataOut_payload_0_7848;
  wire       [7:0]    _zz_dataOut_payload_0_7849;
  wire                _zz_dataOut_payload_0_7850;
  wire       [7:0]    _zz_dataOut_payload_0_7851;
  wire       [7:0]    _zz_dataOut_payload_0_7852;
  wire                _zz_dataOut_payload_0_7853;
  wire       [7:0]    _zz_dataOut_payload_0_7854;
  wire       [7:0]    _zz_dataOut_payload_0_7855;
  wire                _zz_dataOut_payload_0_7856;
  wire       [7:0]    _zz_dataOut_payload_0_7857;
  wire       [7:0]    _zz_dataOut_payload_0_7858;
  wire                _zz_dataOut_payload_0_7859;
  wire       [7:0]    _zz_dataOut_payload_0_7860;
  wire       [7:0]    _zz_dataOut_payload_0_7861;
  wire                _zz_dataOut_payload_0_7862;
  wire                _zz_dataOut_payload_0_7863;
  reg        [7:0]    _zz_dataOut_payload_0_7864;
  reg        [7:0]    _zz_dataOut_payload_0_7865;
  reg        [7:0]    _zz_dataOut_payload_0_7866;
  reg        [7:0]    _zz_dataOut_payload_0_7867;
  wire                _zz_dataOut_payload_0_7868;
  wire       [7:0]    _zz_dataOut_payload_0_7869;
  wire       [7:0]    _zz_dataOut_payload_0_7870;
  wire                _zz_dataOut_payload_0_7871;
  wire       [7:0]    _zz_dataOut_payload_0_7872;
  wire       [7:0]    _zz_dataOut_payload_0_7873;
  wire                _zz_dataOut_payload_0_7874;
  wire                _zz_dataOut_payload_0_7875;
  reg        [7:0]    _zz_dataOut_payload_0_7876;
  reg        [7:0]    _zz_dataOut_payload_0_7877;
  reg        [7:0]    _zz_dataOut_payload_0_7878;
  reg        [7:0]    _zz_dataOut_payload_0_7879;
  reg        [7:0]    _zz_dataOut_payload_0_7880;
  reg        [7:0]    _zz_dataOut_payload_0_7881;
  reg        [7:0]    _zz_dataOut_payload_0_7882;
  reg        [7:0]    _zz_dataOut_payload_0_7883;
  reg        [7:0]    _zz_dataOut_payload_0_7884;
  reg        [7:0]    _zz_dataOut_payload_0_7885;
  reg        [7:0]    _zz_dataOut_payload_0_7886;
  reg        [7:0]    _zz_dataOut_payload_0_7887;
  reg        [7:0]    _zz_dataOut_payload_0_7888;
  reg        [7:0]    _zz_dataOut_payload_0_7889;
  reg        [7:0]    _zz_dataOut_payload_0_7890;
  reg        [7:0]    _zz_dataOut_payload_0_7891;
  reg        [7:0]    _zz_dataOut_payload_0_7892;
  reg        [7:0]    _zz_dataOut_payload_0_7893;
  reg        [7:0]    _zz_dataOut_payload_0_7894;
  reg        [7:0]    _zz_dataOut_payload_0_7895;
  reg        [7:0]    _zz_dataOut_payload_0_7896;
  reg        [7:0]    _zz_dataOut_payload_0_7897;
  reg        [7:0]    _zz_dataOut_payload_0_7898;
  reg        [7:0]    _zz_dataOut_payload_0_7899;
  reg        [7:0]    _zz_dataOut_payload_0_7900;
  reg        [7:0]    _zz_dataOut_payload_0_7901;
  reg        [7:0]    _zz_dataOut_payload_0_7902;
  reg        [7:0]    _zz_dataOut_payload_0_7903;
  wire                _zz_dataOut_payload_0_7904;
  wire       [7:0]    _zz_dataOut_payload_0_7905;
  wire       [7:0]    _zz_dataOut_payload_0_7906;
  wire                _zz_dataOut_payload_0_7907;
  wire       [7:0]    _zz_dataOut_payload_0_7908;
  wire       [7:0]    _zz_dataOut_payload_0_7909;
  wire                _zz_dataOut_payload_0_7910;
  wire       [7:0]    _zz_dataOut_payload_0_7911;
  wire       [7:0]    _zz_dataOut_payload_0_7912;
  wire                _zz_dataOut_payload_0_7913;
  wire       [7:0]    _zz_dataOut_payload_0_7914;
  wire       [7:0]    _zz_dataOut_payload_0_7915;
  wire                _zz_dataOut_payload_0_7916;
  wire       [7:0]    _zz_dataOut_payload_0_7917;
  wire       [7:0]    _zz_dataOut_payload_0_7918;
  wire                _zz_dataOut_payload_0_7919;
  wire       [7:0]    _zz_dataOut_payload_0_7920;
  wire       [7:0]    _zz_dataOut_payload_0_7921;
  wire                _zz_dataOut_payload_0_7922;
  wire       [7:0]    _zz_dataOut_payload_0_7923;
  wire       [7:0]    _zz_dataOut_payload_0_7924;
  wire                _zz_dataOut_payload_0_7925;
  wire       [7:0]    _zz_dataOut_payload_0_7926;
  wire       [7:0]    _zz_dataOut_payload_0_7927;
  wire                _zz_dataOut_payload_0_7928;
  wire       [7:0]    _zz_dataOut_payload_0_7929;
  wire       [7:0]    _zz_dataOut_payload_0_7930;
  wire                _zz_dataOut_payload_0_7931;
  wire       [7:0]    _zz_dataOut_payload_0_7932;
  wire       [7:0]    _zz_dataOut_payload_0_7933;
  wire                _zz_dataOut_payload_0_7934;
  wire       [7:0]    _zz_dataOut_payload_0_7935;
  wire       [7:0]    _zz_dataOut_payload_0_7936;
  wire                _zz_dataOut_payload_0_7937;
  wire       [7:0]    _zz_dataOut_payload_0_7938;
  wire       [7:0]    _zz_dataOut_payload_0_7939;
  wire                _zz_dataOut_payload_0_7940;
  wire       [7:0]    _zz_dataOut_payload_0_7941;
  wire       [7:0]    _zz_dataOut_payload_0_7942;
  wire                _zz_dataOut_payload_0_7943;
  wire       [7:0]    _zz_dataOut_payload_0_7944;
  wire       [7:0]    _zz_dataOut_payload_0_7945;
  wire                _zz_dataOut_payload_0_7946;
  wire                _zz_dataOut_payload_0_7947;
  reg        [7:0]    _zz_dataOut_payload_0_7948;
  reg        [7:0]    _zz_dataOut_payload_0_7949;
  reg        [7:0]    _zz_dataOut_payload_0_7950;
  reg        [7:0]    _zz_dataOut_payload_0_7951;
  wire                _zz_dataOut_payload_0_7952;
  wire       [7:0]    _zz_dataOut_payload_0_7953;
  wire       [7:0]    _zz_dataOut_payload_0_7954;
  wire                _zz_dataOut_payload_0_7955;
  wire       [7:0]    _zz_dataOut_payload_0_7956;
  wire       [7:0]    _zz_dataOut_payload_0_7957;
  wire                _zz_dataOut_payload_0_7958;
  wire                _zz_dataOut_payload_0_7959;
  reg        [7:0]    _zz_dataOut_payload_0_7960;
  reg        [7:0]    _zz_dataOut_payload_0_7961;
  reg        [7:0]    _zz_dataOut_payload_0_7962;
  reg        [7:0]    _zz_dataOut_payload_0_7963;
  reg        [7:0]    _zz_dataOut_payload_0_7964;
  reg        [7:0]    _zz_dataOut_payload_0_7965;
  reg        [7:0]    _zz_dataOut_payload_0_7966;
  reg        [7:0]    _zz_dataOut_payload_0_7967;
  reg        [7:0]    _zz_dataOut_payload_0_7968;
  reg        [7:0]    _zz_dataOut_payload_0_7969;
  reg        [7:0]    _zz_dataOut_payload_0_7970;
  reg        [7:0]    _zz_dataOut_payload_0_7971;
  wire                _zz_dataOut_payload_0_7972;
  wire       [7:0]    _zz_dataOut_payload_0_7973;
  wire       [7:0]    _zz_dataOut_payload_0_7974;
  wire                _zz_dataOut_payload_0_7975;
  wire       [7:0]    _zz_dataOut_payload_0_7976;
  wire       [7:0]    _zz_dataOut_payload_0_7977;
  wire                _zz_dataOut_payload_0_7978;
  wire       [7:0]    _zz_dataOut_payload_0_7979;
  wire       [7:0]    _zz_dataOut_payload_0_7980;
  wire                _zz_dataOut_payload_0_7981;
  wire       [7:0]    _zz_dataOut_payload_0_7982;
  wire       [7:0]    _zz_dataOut_payload_0_7983;
  wire                _zz_dataOut_payload_0_7984;
  wire       [7:0]    _zz_dataOut_payload_0_7985;
  wire       [7:0]    _zz_dataOut_payload_0_7986;
  wire                _zz_dataOut_payload_0_7987;
  wire       [7:0]    _zz_dataOut_payload_0_7988;
  wire       [7:0]    _zz_dataOut_payload_0_7989;
  wire                _zz_dataOut_payload_0_7990;
  wire                _zz_dataOut_payload_0_7991;
  reg        [7:0]    _zz_dataOut_payload_0_7992;
  reg        [7:0]    _zz_dataOut_payload_0_7993;
  reg        [7:0]    _zz_dataOut_payload_0_7994;
  reg        [7:0]    _zz_dataOut_payload_0_7995;
  wire                _zz_dataOut_payload_0_7996;
  wire       [7:0]    _zz_dataOut_payload_0_7997;
  wire       [7:0]    _zz_dataOut_payload_0_7998;
  wire                _zz_dataOut_payload_0_7999;
  wire       [7:0]    _zz_dataOut_payload_0_8000;
  wire       [7:0]    _zz_dataOut_payload_0_8001;
  wire                _zz_dataOut_payload_0_8002;
  wire                _zz_dataOut_payload_0_8003;
  reg        [7:0]    _zz_dataOut_payload_0_8004;
  reg        [7:0]    _zz_dataOut_payload_0_8005;
  reg        [7:0]    _zz_dataOut_payload_0_8006;
  reg        [7:0]    _zz_dataOut_payload_0_8007;
  reg        [7:0]    _zz_dataOut_payload_0_8008;
  reg        [7:0]    _zz_dataOut_payload_0_8009;
  reg        [7:0]    _zz_dataOut_payload_0_8010;
  reg        [7:0]    _zz_dataOut_payload_0_8011;
  reg        [7:0]    _zz_dataOut_payload_0_8012;
  reg        [7:0]    _zz_dataOut_payload_0_8013;
  reg        [7:0]    _zz_dataOut_payload_0_8014;
  reg        [7:0]    _zz_dataOut_payload_0_8015;
  reg        [7:0]    _zz_dataOut_payload_0_8016;
  reg        [7:0]    _zz_dataOut_payload_0_8017;
  reg        [7:0]    _zz_dataOut_payload_0_8018;
  reg        [7:0]    _zz_dataOut_payload_0_8019;
  reg        [7:0]    _zz_dataOut_payload_0_8020;
  reg        [7:0]    _zz_dataOut_payload_0_8021;
  reg        [7:0]    _zz_dataOut_payload_0_8022;
  reg        [7:0]    _zz_dataOut_payload_0_8023;
  reg        [7:0]    _zz_dataOut_payload_0_8024;
  reg        [7:0]    _zz_dataOut_payload_0_8025;
  reg        [7:0]    _zz_dataOut_payload_0_8026;
  reg        [7:0]    _zz_dataOut_payload_0_8027;
  reg        [7:0]    _zz_dataOut_payload_0_8028;
  reg        [7:0]    _zz_dataOut_payload_0_8029;
  reg        [7:0]    _zz_dataOut_payload_0_8030;
  reg        [7:0]    _zz_dataOut_payload_0_8031;
  reg        [7:0]    _zz_dataOut_payload_0_8032;
  reg        [7:0]    _zz_dataOut_payload_0_8033;
  reg        [7:0]    _zz_dataOut_payload_0_8034;
  reg        [7:0]    _zz_dataOut_payload_0_8035;
  reg        [7:0]    _zz_dataOut_payload_0_8036;
  reg        [7:0]    _zz_dataOut_payload_0_8037;
  reg        [7:0]    _zz_dataOut_payload_0_8038;
  reg        [7:0]    _zz_dataOut_payload_0_8039;
  reg        [7:0]    _zz_dataOut_payload_0_8040;
  reg        [7:0]    _zz_dataOut_payload_0_8041;
  reg        [7:0]    _zz_dataOut_payload_0_8042;
  reg        [7:0]    _zz_dataOut_payload_0_8043;
  reg        [7:0]    _zz_dataOut_payload_0_8044;
  reg        [7:0]    _zz_dataOut_payload_0_8045;
  reg        [7:0]    _zz_dataOut_payload_0_8046;
  reg        [7:0]    _zz_dataOut_payload_0_8047;
  reg        [7:0]    _zz_dataOut_payload_0_8048;
  reg        [7:0]    _zz_dataOut_payload_0_8049;
  reg        [7:0]    _zz_dataOut_payload_0_8050;
  reg        [7:0]    _zz_dataOut_payload_0_8051;
  reg        [7:0]    _zz_dataOut_payload_0_8052;
  reg        [7:0]    _zz_dataOut_payload_0_8053;
  reg        [7:0]    _zz_dataOut_payload_0_8054;
  reg        [7:0]    _zz_dataOut_payload_0_8055;
  reg        [7:0]    _zz_dataOut_payload_0_8056;
  reg        [7:0]    _zz_dataOut_payload_0_8057;
  reg        [7:0]    _zz_dataOut_payload_0_8058;
  reg        [7:0]    _zz_dataOut_payload_0_8059;
  reg        [7:0]    _zz_dataOut_payload_0_8060;
  reg        [7:0]    _zz_dataOut_payload_0_8061;
  reg        [7:0]    _zz_dataOut_payload_0_8062;
  reg        [7:0]    _zz_dataOut_payload_0_8063;
  reg        [7:0]    _zz_dataOut_payload_0_8064;
  reg        [7:0]    _zz_dataOut_payload_0_8065;
  reg        [7:0]    _zz_dataOut_payload_0_8066;
  reg        [7:0]    _zz_dataOut_payload_0_8067;
  reg        [7:0]    _zz_dataOut_payload_0_8068;
  reg        [7:0]    _zz_dataOut_payload_0_8069;
  reg        [7:0]    _zz_dataOut_payload_0_8070;
  reg        [7:0]    _zz_dataOut_payload_0_8071;
  reg        [7:0]    _zz_dataOut_payload_0_8072;
  reg        [7:0]    _zz_dataOut_payload_0_8073;
  reg        [7:0]    _zz_dataOut_payload_0_8074;
  reg        [7:0]    _zz_dataOut_payload_0_8075;
  reg        [7:0]    _zz_dataOut_payload_0_8076;
  reg        [7:0]    _zz_dataOut_payload_0_8077;
  reg        [7:0]    _zz_dataOut_payload_0_8078;
  reg        [7:0]    _zz_dataOut_payload_0_8079;
  reg        [7:0]    _zz_dataOut_payload_0_8080;
  reg        [7:0]    _zz_dataOut_payload_0_8081;
  reg        [7:0]    _zz_dataOut_payload_0_8082;
  reg        [7:0]    _zz_dataOut_payload_0_8083;
  reg        [7:0]    _zz_dataOut_payload_0_8084;
  reg        [7:0]    _zz_dataOut_payload_0_8085;
  reg        [7:0]    _zz_dataOut_payload_0_8086;
  reg        [7:0]    _zz_dataOut_payload_0_8087;
  reg        [7:0]    _zz_dataOut_payload_0_8088;
  reg        [7:0]    _zz_dataOut_payload_0_8089;
  reg        [7:0]    _zz_dataOut_payload_0_8090;
  reg        [7:0]    _zz_dataOut_payload_0_8091;
  reg        [7:0]    _zz_dataOut_payload_0_8092;
  reg        [7:0]    _zz_dataOut_payload_0_8093;
  reg        [7:0]    _zz_dataOut_payload_0_8094;
  reg        [7:0]    _zz_dataOut_payload_0_8095;
  reg        [7:0]    _zz_dataOut_payload_0_8096;
  reg        [7:0]    _zz_dataOut_payload_0_8097;
  reg        [7:0]    _zz_dataOut_payload_0_8098;
  reg        [7:0]    _zz_dataOut_payload_0_8099;
  reg        [7:0]    _zz_dataOut_payload_0_8100;
  reg        [7:0]    _zz_dataOut_payload_0_8101;
  reg        [7:0]    _zz_dataOut_payload_0_8102;
  reg        [7:0]    _zz_dataOut_payload_0_8103;
  reg        [7:0]    _zz_dataOut_payload_0_8104;
  reg        [7:0]    _zz_dataOut_payload_0_8105;
  reg        [7:0]    _zz_dataOut_payload_0_8106;
  reg        [7:0]    _zz_dataOut_payload_0_8107;
  reg        [7:0]    _zz_dataOut_payload_0_8108;
  reg        [7:0]    _zz_dataOut_payload_0_8109;
  reg        [7:0]    _zz_dataOut_payload_0_8110;
  reg        [7:0]    _zz_dataOut_payload_0_8111;
  reg        [7:0]    _zz_dataOut_payload_0_8112;
  reg        [7:0]    _zz_dataOut_payload_0_8113;
  reg        [7:0]    _zz_dataOut_payload_0_8114;
  reg        [7:0]    _zz_dataOut_payload_0_8115;
  reg        [7:0]    _zz_dataOut_payload_0_8116;
  reg        [7:0]    _zz_dataOut_payload_0_8117;
  reg        [7:0]    _zz_dataOut_payload_0_8118;
  reg        [7:0]    _zz_dataOut_payload_0_8119;
  reg        [7:0]    _zz_dataOut_payload_0_8120;
  reg        [7:0]    _zz_dataOut_payload_0_8121;
  reg        [7:0]    _zz_dataOut_payload_0_8122;
  reg        [7:0]    _zz_dataOut_payload_0_8123;
  reg        [7:0]    _zz_dataOut_payload_0_8124;
  reg        [7:0]    _zz_dataOut_payload_0_8125;
  reg        [7:0]    _zz_dataOut_payload_0_8126;
  reg        [7:0]    _zz_dataOut_payload_0_8127;
  reg        [7:0]    _zz_dataOut_payload_0_8128;
  reg        [7:0]    _zz_dataOut_payload_0_8129;
  reg        [7:0]    _zz_dataOut_payload_0_8130;
  reg        [7:0]    _zz_dataOut_payload_0_8131;
  reg        [7:0]    _zz_dataOut_payload_0_8132;
  reg        [7:0]    _zz_dataOut_payload_0_8133;
  reg        [7:0]    _zz_dataOut_payload_0_8134;
  reg        [7:0]    _zz_dataOut_payload_0_8135;
  reg        [7:0]    _zz_dataOut_payload_0_8136;
  reg        [7:0]    _zz_dataOut_payload_0_8137;
  reg        [7:0]    _zz_dataOut_payload_0_8138;
  reg        [7:0]    _zz_dataOut_payload_0_8139;
  reg        [7:0]    _zz_dataOut_payload_0_8140;
  reg        [7:0]    _zz_dataOut_payload_0_8141;
  reg        [7:0]    _zz_dataOut_payload_0_8142;
  reg        [7:0]    _zz_dataOut_payload_0_8143;
  reg        [7:0]    _zz_dataOut_payload_0_8144;
  reg        [7:0]    _zz_dataOut_payload_0_8145;
  reg        [7:0]    _zz_dataOut_payload_0_8146;
  reg        [7:0]    _zz_dataOut_payload_0_8147;
  reg        [7:0]    _zz_dataOut_payload_0_8148;
  reg        [7:0]    _zz_dataOut_payload_0_8149;
  reg        [7:0]    _zz_dataOut_payload_0_8150;
  reg        [7:0]    _zz_dataOut_payload_0_8151;
  reg        [7:0]    _zz_dataOut_payload_0_8152;
  reg        [7:0]    _zz_dataOut_payload_0_8153;
  reg        [7:0]    _zz_dataOut_payload_0_8154;
  reg        [7:0]    _zz_dataOut_payload_0_8155;
  reg        [7:0]    _zz_dataOut_payload_0_8156;
  reg        [7:0]    _zz_dataOut_payload_0_8157;
  reg        [7:0]    _zz_dataOut_payload_0_8158;
  reg        [7:0]    _zz_dataOut_payload_0_8159;
  reg        [7:0]    _zz_dataOut_payload_0_8160;
  reg        [7:0]    _zz_dataOut_payload_0_8161;
  reg        [7:0]    _zz_dataOut_payload_0_8162;
  reg        [7:0]    _zz_dataOut_payload_0_8163;
  reg        [7:0]    _zz_dataOut_payload_0_8164;
  reg        [7:0]    _zz_dataOut_payload_0_8165;
  reg        [7:0]    _zz_dataOut_payload_0_8166;
  reg        [7:0]    _zz_dataOut_payload_0_8167;
  reg        [7:0]    _zz_dataOut_payload_0_8168;
  reg        [7:0]    _zz_dataOut_payload_0_8169;
  reg        [7:0]    _zz_dataOut_payload_0_8170;
  reg        [7:0]    _zz_dataOut_payload_0_8171;
  reg        [7:0]    _zz_dataOut_payload_0_8172;
  reg        [7:0]    _zz_dataOut_payload_0_8173;
  reg        [7:0]    _zz_dataOut_payload_0_8174;
  reg        [7:0]    _zz_dataOut_payload_0_8175;
  reg        [7:0]    _zz_dataOut_payload_0_8176;
  reg        [7:0]    _zz_dataOut_payload_0_8177;
  reg        [7:0]    _zz_dataOut_payload_0_8178;
  reg        [7:0]    _zz_dataOut_payload_0_8179;
  reg        [7:0]    _zz_dataOut_payload_0_8180;
  reg        [7:0]    _zz_dataOut_payload_0_8181;
  reg        [7:0]    _zz_dataOut_payload_0_8182;
  reg        [7:0]    _zz_dataOut_payload_0_8183;
  reg        [7:0]    _zz_dataOut_payload_0_8184;
  reg        [7:0]    _zz_dataOut_payload_0_8185;
  reg        [7:0]    _zz_dataOut_payload_0_8186;
  reg        [7:0]    _zz_dataOut_payload_0_8187;
  reg        [7:0]    _zz_dataOut_payload_0_8188;
  reg        [7:0]    _zz_dataOut_payload_0_8189;
  reg        [7:0]    _zz_dataOut_payload_0_8190;
  reg        [7:0]    _zz_dataOut_payload_0_8191;
  reg        [7:0]    _zz_dataOut_payload_0_8192;
  reg        [7:0]    _zz_dataOut_payload_0_8193;
  reg        [7:0]    _zz_dataOut_payload_0_8194;
  reg        [7:0]    _zz_dataOut_payload_0_8195;
  reg        [7:0]    _zz_dataOut_payload_0_8196;
  reg        [7:0]    _zz_dataOut_payload_0_8197;
  reg        [7:0]    _zz_dataOut_payload_0_8198;
  reg        [7:0]    _zz_dataOut_payload_0_8199;
  reg        [7:0]    _zz_dataOut_payload_0_8200;
  reg        [7:0]    _zz_dataOut_payload_0_8201;
  reg        [7:0]    _zz_dataOut_payload_0_8202;
  reg        [7:0]    _zz_dataOut_payload_0_8203;
  reg        [7:0]    _zz_dataOut_payload_0_8204;
  reg        [7:0]    _zz_dataOut_payload_0_8205;
  reg        [7:0]    _zz_dataOut_payload_0_8206;
  reg        [7:0]    _zz_dataOut_payload_0_8207;
  reg        [7:0]    _zz_dataOut_payload_0_8208;
  reg        [7:0]    _zz_dataOut_payload_0_8209;
  reg        [7:0]    _zz_dataOut_payload_0_8210;
  reg        [7:0]    _zz_dataOut_payload_0_8211;
  reg        [7:0]    _zz_dataOut_payload_0_8212;
  reg        [7:0]    _zz_dataOut_payload_0_8213;
  reg        [7:0]    _zz_dataOut_payload_0_8214;
  reg        [7:0]    _zz_dataOut_payload_0_8215;
  reg        [7:0]    _zz_dataOut_payload_0_8216;
  reg        [7:0]    _zz_dataOut_payload_0_8217;
  reg        [7:0]    _zz_dataOut_payload_0_8218;
  reg        [7:0]    _zz_dataOut_payload_0_8219;
  reg        [7:0]    _zz_dataOut_payload_0_8220;
  reg        [7:0]    _zz_dataOut_payload_0_8221;
  reg        [7:0]    _zz_dataOut_payload_0_8222;
  reg        [7:0]    _zz_dataOut_payload_0_8223;
  reg        [7:0]    _zz_dataOut_payload_0_8224;
  reg        [7:0]    _zz_dataOut_payload_0_8225;
  reg        [7:0]    _zz_dataOut_payload_0_8226;
  reg        [7:0]    _zz_dataOut_payload_0_8227;
  reg        [7:0]    _zz_dataOut_payload_0_8228;
  reg        [7:0]    _zz_dataOut_payload_0_8229;
  reg        [7:0]    _zz_dataOut_payload_0_8230;
  reg        [7:0]    _zz_dataOut_payload_0_8231;
  reg        [7:0]    _zz_dataOut_payload_0_8232;
  reg        [7:0]    _zz_dataOut_payload_0_8233;
  reg        [7:0]    _zz_dataOut_payload_0_8234;
  reg        [7:0]    _zz_dataOut_payload_0_8235;
  reg        [7:0]    _zz_dataOut_payload_0_8236;
  reg        [7:0]    _zz_dataOut_payload_0_8237;
  reg        [7:0]    _zz_dataOut_payload_0_8238;
  reg        [7:0]    _zz_dataOut_payload_0_8239;
  reg        [7:0]    _zz_dataOut_payload_0_8240;
  reg        [7:0]    _zz_dataOut_payload_0_8241;
  reg        [7:0]    _zz_dataOut_payload_0_8242;
  reg        [7:0]    _zz_dataOut_payload_0_8243;
  reg        [7:0]    _zz_dataOut_payload_0_8244;
  reg        [7:0]    _zz_dataOut_payload_0_8245;
  reg        [7:0]    _zz_dataOut_payload_0_8246;
  reg        [7:0]    _zz_dataOut_payload_0_8247;
  reg        [7:0]    _zz_dataOut_payload_0_8248;
  reg        [7:0]    _zz_dataOut_payload_0_8249;
  reg        [7:0]    _zz_dataOut_payload_0_8250;
  reg        [7:0]    _zz_dataOut_payload_0_8251;
  reg        [7:0]    _zz_dataOut_payload_0_8252;
  reg        [7:0]    _zz_dataOut_payload_0_8253;
  reg        [7:0]    _zz_dataOut_payload_0_8254;
  reg        [7:0]    _zz_dataOut_payload_0_8255;
  reg        [7:0]    _zz_dataOut_payload_0_8256;
  reg        [7:0]    _zz_dataOut_payload_0_8257;
  reg        [7:0]    _zz_dataOut_payload_0_8258;
  reg        [7:0]    _zz_dataOut_payload_0_8259;
  reg        [7:0]    _zz_dataOut_payload_0_8260;
  reg        [7:0]    _zz_dataOut_payload_0_8261;
  reg        [7:0]    _zz_dataOut_payload_0_8262;
  reg        [7:0]    _zz_dataOut_payload_0_8263;
  reg        [7:0]    _zz_dataOut_payload_0_8264;
  reg        [7:0]    _zz_dataOut_payload_0_8265;
  reg        [7:0]    _zz_dataOut_payload_0_8266;
  reg        [7:0]    _zz_dataOut_payload_0_8267;
  reg        [7:0]    _zz_dataOut_payload_0_8268;
  reg        [7:0]    _zz_dataOut_payload_0_8269;
  reg        [7:0]    _zz_dataOut_payload_0_8270;
  reg        [7:0]    _zz_dataOut_payload_0_8271;
  reg        [7:0]    _zz_dataOut_payload_0_8272;
  reg        [7:0]    _zz_dataOut_payload_0_8273;
  reg        [7:0]    _zz_dataOut_payload_0_8274;
  reg        [7:0]    _zz_dataOut_payload_0_8275;
  reg        [7:0]    _zz_dataOut_payload_0_8276;
  reg        [7:0]    _zz_dataOut_payload_0_8277;
  reg        [7:0]    _zz_dataOut_payload_0_8278;
  reg        [7:0]    _zz_dataOut_payload_0_8279;
  reg        [7:0]    _zz_dataOut_payload_0_8280;
  reg        [7:0]    _zz_dataOut_payload_0_8281;
  reg        [7:0]    _zz_dataOut_payload_0_8282;
  reg        [7:0]    _zz_dataOut_payload_0_8283;
  reg        [7:0]    _zz_dataOut_payload_0_8284;
  reg        [7:0]    _zz_dataOut_payload_0_8285;
  reg        [7:0]    _zz_dataOut_payload_0_8286;
  reg        [7:0]    _zz_dataOut_payload_0_8287;
  reg        [7:0]    _zz_dataOut_payload_0_8288;
  reg        [7:0]    _zz_dataOut_payload_0_8289;
  reg        [7:0]    _zz_dataOut_payload_0_8290;
  reg        [7:0]    _zz_dataOut_payload_0_8291;
  reg        [7:0]    _zz_dataOut_payload_0_8292;
  reg        [7:0]    _zz_dataOut_payload_0_8293;
  reg        [7:0]    _zz_dataOut_payload_0_8294;
  reg        [7:0]    _zz_dataOut_payload_0_8295;
  reg        [7:0]    _zz_dataOut_payload_0_8296;
  reg        [7:0]    _zz_dataOut_payload_0_8297;
  reg        [7:0]    _zz_dataOut_payload_0_8298;
  reg        [7:0]    _zz_dataOut_payload_0_8299;
  reg        [7:0]    _zz_dataOut_payload_0_8300;
  reg        [7:0]    _zz_dataOut_payload_0_8301;
  reg        [7:0]    _zz_dataOut_payload_0_8302;
  reg        [7:0]    _zz_dataOut_payload_0_8303;
  reg        [7:0]    _zz_dataOut_payload_0_8304;
  reg        [7:0]    _zz_dataOut_payload_0_8305;
  reg        [7:0]    _zz_dataOut_payload_0_8306;
  reg        [7:0]    _zz_dataOut_payload_0_8307;
  reg        [7:0]    _zz_dataOut_payload_0_8308;
  reg        [7:0]    _zz_dataOut_payload_0_8309;
  reg        [7:0]    _zz_dataOut_payload_0_8310;
  reg        [7:0]    _zz_dataOut_payload_0_8311;
  reg        [7:0]    _zz_dataOut_payload_0_8312;
  reg        [7:0]    _zz_dataOut_payload_0_8313;
  reg        [7:0]    _zz_dataOut_payload_0_8314;
  reg        [7:0]    _zz_dataOut_payload_0_8315;
  reg        [7:0]    _zz_dataOut_payload_0_8316;
  reg        [7:0]    _zz_dataOut_payload_0_8317;
  reg        [7:0]    _zz_dataOut_payload_0_8318;
  reg        [7:0]    _zz_dataOut_payload_0_8319;
  wire                _zz_dataOut_payload_0_8320;
  wire       [7:0]    _zz_dataOut_payload_0_8321;
  wire       [7:0]    _zz_dataOut_payload_0_8322;
  wire                _zz_dataOut_payload_0_8323;
  wire       [7:0]    _zz_dataOut_payload_0_8324;
  wire       [7:0]    _zz_dataOut_payload_0_8325;
  wire                _zz_dataOut_payload_0_8326;
  wire       [7:0]    _zz_dataOut_payload_0_8327;
  wire       [7:0]    _zz_dataOut_payload_0_8328;
  wire                _zz_dataOut_payload_0_8329;
  wire       [7:0]    _zz_dataOut_payload_0_8330;
  wire       [7:0]    _zz_dataOut_payload_0_8331;
  wire                _zz_dataOut_payload_0_8332;
  wire       [7:0]    _zz_dataOut_payload_0_8333;
  wire       [7:0]    _zz_dataOut_payload_0_8334;
  wire                _zz_dataOut_payload_0_8335;
  wire       [7:0]    _zz_dataOut_payload_0_8336;
  wire       [7:0]    _zz_dataOut_payload_0_8337;
  wire                _zz_dataOut_payload_0_8338;
  wire       [7:0]    _zz_dataOut_payload_0_8339;
  wire       [7:0]    _zz_dataOut_payload_0_8340;
  wire                _zz_dataOut_payload_0_8341;
  wire       [7:0]    _zz_dataOut_payload_0_8342;
  wire       [7:0]    _zz_dataOut_payload_0_8343;
  wire                _zz_dataOut_payload_0_8344;
  wire       [7:0]    _zz_dataOut_payload_0_8345;
  wire       [7:0]    _zz_dataOut_payload_0_8346;
  wire                _zz_dataOut_payload_0_8347;
  wire       [7:0]    _zz_dataOut_payload_0_8348;
  wire       [7:0]    _zz_dataOut_payload_0_8349;
  wire                _zz_dataOut_payload_0_8350;
  wire       [7:0]    _zz_dataOut_payload_0_8351;
  wire       [7:0]    _zz_dataOut_payload_0_8352;
  wire                _zz_dataOut_payload_0_8353;
  wire       [7:0]    _zz_dataOut_payload_0_8354;
  wire       [7:0]    _zz_dataOut_payload_0_8355;
  wire                _zz_dataOut_payload_0_8356;
  wire       [7:0]    _zz_dataOut_payload_0_8357;
  wire       [7:0]    _zz_dataOut_payload_0_8358;
  wire                _zz_dataOut_payload_0_8359;
  wire       [7:0]    _zz_dataOut_payload_0_8360;
  wire       [7:0]    _zz_dataOut_payload_0_8361;
  wire                _zz_dataOut_payload_0_8362;
  wire       [7:0]    _zz_dataOut_payload_0_8363;
  wire       [7:0]    _zz_dataOut_payload_0_8364;
  wire                _zz_dataOut_payload_0_8365;
  wire       [7:0]    _zz_dataOut_payload_0_8366;
  wire       [7:0]    _zz_dataOut_payload_0_8367;
  wire                _zz_dataOut_payload_0_8368;
  wire       [7:0]    _zz_dataOut_payload_0_8369;
  wire       [7:0]    _zz_dataOut_payload_0_8370;
  wire                _zz_dataOut_payload_0_8371;
  wire       [7:0]    _zz_dataOut_payload_0_8372;
  wire       [7:0]    _zz_dataOut_payload_0_8373;
  wire                _zz_dataOut_payload_0_8374;
  wire       [7:0]    _zz_dataOut_payload_0_8375;
  wire       [7:0]    _zz_dataOut_payload_0_8376;
  wire                _zz_dataOut_payload_0_8377;
  wire       [7:0]    _zz_dataOut_payload_0_8378;
  wire       [7:0]    _zz_dataOut_payload_0_8379;
  wire                _zz_dataOut_payload_0_8380;
  wire       [7:0]    _zz_dataOut_payload_0_8381;
  wire       [7:0]    _zz_dataOut_payload_0_8382;
  wire                _zz_dataOut_payload_0_8383;
  wire       [7:0]    _zz_dataOut_payload_0_8384;
  wire       [7:0]    _zz_dataOut_payload_0_8385;
  wire                _zz_dataOut_payload_0_8386;
  wire       [7:0]    _zz_dataOut_payload_0_8387;
  wire       [7:0]    _zz_dataOut_payload_0_8388;
  wire                _zz_dataOut_payload_0_8389;
  wire       [7:0]    _zz_dataOut_payload_0_8390;
  wire       [7:0]    _zz_dataOut_payload_0_8391;
  wire                _zz_dataOut_payload_0_8392;
  wire       [7:0]    _zz_dataOut_payload_0_8393;
  wire       [7:0]    _zz_dataOut_payload_0_8394;
  wire                _zz_dataOut_payload_0_8395;
  wire       [7:0]    _zz_dataOut_payload_0_8396;
  wire       [7:0]    _zz_dataOut_payload_0_8397;
  wire                _zz_dataOut_payload_0_8398;
  wire       [7:0]    _zz_dataOut_payload_0_8399;
  wire       [7:0]    _zz_dataOut_payload_0_8400;
  wire                _zz_dataOut_payload_0_8401;
  wire       [7:0]    _zz_dataOut_payload_0_8402;
  wire       [7:0]    _zz_dataOut_payload_0_8403;
  wire                _zz_dataOut_payload_0_8404;
  wire       [7:0]    _zz_dataOut_payload_0_8405;
  wire       [7:0]    _zz_dataOut_payload_0_8406;
  wire                _zz_dataOut_payload_0_8407;
  wire       [7:0]    _zz_dataOut_payload_0_8408;
  wire       [7:0]    _zz_dataOut_payload_0_8409;
  wire                _zz_dataOut_payload_0_8410;
  wire       [7:0]    _zz_dataOut_payload_0_8411;
  wire       [7:0]    _zz_dataOut_payload_0_8412;
  wire                _zz_dataOut_payload_0_8413;
  wire       [7:0]    _zz_dataOut_payload_0_8414;
  wire       [7:0]    _zz_dataOut_payload_0_8415;
  wire                _zz_dataOut_payload_0_8416;
  wire       [7:0]    _zz_dataOut_payload_0_8417;
  wire       [7:0]    _zz_dataOut_payload_0_8418;
  wire                _zz_dataOut_payload_0_8419;
  wire       [7:0]    _zz_dataOut_payload_0_8420;
  wire       [7:0]    _zz_dataOut_payload_0_8421;
  wire                _zz_dataOut_payload_0_8422;
  wire       [7:0]    _zz_dataOut_payload_0_8423;
  wire       [7:0]    _zz_dataOut_payload_0_8424;
  wire                _zz_dataOut_payload_0_8425;
  wire       [7:0]    _zz_dataOut_payload_0_8426;
  wire       [7:0]    _zz_dataOut_payload_0_8427;
  wire                _zz_dataOut_payload_0_8428;
  wire       [7:0]    _zz_dataOut_payload_0_8429;
  wire       [7:0]    _zz_dataOut_payload_0_8430;
  wire                _zz_dataOut_payload_0_8431;
  wire       [7:0]    _zz_dataOut_payload_0_8432;
  wire       [7:0]    _zz_dataOut_payload_0_8433;
  wire                _zz_dataOut_payload_0_8434;
  wire       [7:0]    _zz_dataOut_payload_0_8435;
  wire       [7:0]    _zz_dataOut_payload_0_8436;
  wire                _zz_dataOut_payload_0_8437;
  wire       [7:0]    _zz_dataOut_payload_0_8438;
  wire       [7:0]    _zz_dataOut_payload_0_8439;
  wire                _zz_dataOut_payload_0_8440;
  wire       [7:0]    _zz_dataOut_payload_0_8441;
  wire       [7:0]    _zz_dataOut_payload_0_8442;
  wire                _zz_dataOut_payload_0_8443;
  wire       [7:0]    _zz_dataOut_payload_0_8444;
  wire       [7:0]    _zz_dataOut_payload_0_8445;
  wire                _zz_dataOut_payload_0_8446;
  wire       [7:0]    _zz_dataOut_payload_0_8447;
  wire       [7:0]    _zz_dataOut_payload_0_8448;
  wire                _zz_dataOut_payload_0_8449;
  wire       [7:0]    _zz_dataOut_payload_0_8450;
  wire       [7:0]    _zz_dataOut_payload_0_8451;
  wire                _zz_dataOut_payload_0_8452;
  wire       [7:0]    _zz_dataOut_payload_0_8453;
  wire       [7:0]    _zz_dataOut_payload_0_8454;
  wire                _zz_dataOut_payload_0_8455;
  wire       [7:0]    _zz_dataOut_payload_0_8456;
  wire       [7:0]    _zz_dataOut_payload_0_8457;
  wire                _zz_dataOut_payload_0_8458;
  wire       [7:0]    _zz_dataOut_payload_0_8459;
  wire       [7:0]    _zz_dataOut_payload_0_8460;
  wire                _zz_dataOut_payload_0_8461;
  wire       [7:0]    _zz_dataOut_payload_0_8462;
  wire       [7:0]    _zz_dataOut_payload_0_8463;
  wire                _zz_dataOut_payload_0_8464;
  wire       [7:0]    _zz_dataOut_payload_0_8465;
  wire       [7:0]    _zz_dataOut_payload_0_8466;
  wire                _zz_dataOut_payload_0_8467;
  wire       [7:0]    _zz_dataOut_payload_0_8468;
  wire       [7:0]    _zz_dataOut_payload_0_8469;
  wire                _zz_dataOut_payload_0_8470;
  wire       [7:0]    _zz_dataOut_payload_0_8471;
  wire       [7:0]    _zz_dataOut_payload_0_8472;
  wire                _zz_dataOut_payload_0_8473;
  wire       [7:0]    _zz_dataOut_payload_0_8474;
  wire       [7:0]    _zz_dataOut_payload_0_8475;
  wire                _zz_dataOut_payload_0_8476;
  wire       [7:0]    _zz_dataOut_payload_0_8477;
  wire       [7:0]    _zz_dataOut_payload_0_8478;
  wire                _zz_dataOut_payload_0_8479;
  wire       [7:0]    _zz_dataOut_payload_0_8480;
  wire       [7:0]    _zz_dataOut_payload_0_8481;
  wire                _zz_dataOut_payload_0_8482;
  wire       [7:0]    _zz_dataOut_payload_0_8483;
  wire       [7:0]    _zz_dataOut_payload_0_8484;
  wire                _zz_dataOut_payload_0_8485;
  wire       [7:0]    _zz_dataOut_payload_0_8486;
  wire       [7:0]    _zz_dataOut_payload_0_8487;
  wire                _zz_dataOut_payload_0_8488;
  wire       [7:0]    _zz_dataOut_payload_0_8489;
  wire       [7:0]    _zz_dataOut_payload_0_8490;
  wire                _zz_dataOut_payload_0_8491;
  wire       [7:0]    _zz_dataOut_payload_0_8492;
  wire       [7:0]    _zz_dataOut_payload_0_8493;
  wire                _zz_dataOut_payload_0_8494;
  wire       [7:0]    _zz_dataOut_payload_0_8495;
  wire       [7:0]    _zz_dataOut_payload_0_8496;
  wire                _zz_dataOut_payload_0_8497;
  wire       [7:0]    _zz_dataOut_payload_0_8498;
  wire       [7:0]    _zz_dataOut_payload_0_8499;
  wire                _zz_dataOut_payload_0_8500;
  wire       [7:0]    _zz_dataOut_payload_0_8501;
  wire       [7:0]    _zz_dataOut_payload_0_8502;
  wire                _zz_dataOut_payload_0_8503;
  wire       [7:0]    _zz_dataOut_payload_0_8504;
  wire       [7:0]    _zz_dataOut_payload_0_8505;
  wire                _zz_dataOut_payload_0_8506;
  wire                _zz_dataOut_payload_0_8507;
  reg        [7:0]    _zz_dataOut_payload_0_8508;
  reg        [7:0]    _zz_dataOut_payload_0_8509;
  reg        [7:0]    _zz_dataOut_payload_0_8510;
  reg        [7:0]    _zz_dataOut_payload_0_8511;
  wire                _zz_dataOut_payload_0_8512;
  wire       [7:0]    _zz_dataOut_payload_0_8513;
  wire       [7:0]    _zz_dataOut_payload_0_8514;
  wire                _zz_dataOut_payload_0_8515;
  wire       [7:0]    _zz_dataOut_payload_0_8516;
  wire       [7:0]    _zz_dataOut_payload_0_8517;
  wire                _zz_dataOut_payload_0_8518;
  wire                _zz_dataOut_payload_0_8519;
  reg        [7:0]    _zz_dataOut_payload_0_8520;
  reg        [7:0]    _zz_dataOut_payload_0_8521;
  reg        [7:0]    _zz_dataOut_payload_0_8522;
  reg        [7:0]    _zz_dataOut_payload_0_8523;
  reg        [7:0]    _zz_dataOut_payload_0_8524;
  reg        [7:0]    _zz_dataOut_payload_0_8525;
  reg        [7:0]    _zz_dataOut_payload_0_8526;
  reg        [7:0]    _zz_dataOut_payload_0_8527;
  reg        [7:0]    _zz_dataOut_payload_0_8528;
  reg        [7:0]    _zz_dataOut_payload_0_8529;
  reg        [7:0]    _zz_dataOut_payload_0_8530;
  reg        [7:0]    _zz_dataOut_payload_0_8531;
  wire                _zz_dataOut_payload_0_8532;
  wire       [7:0]    _zz_dataOut_payload_0_8533;
  wire       [7:0]    _zz_dataOut_payload_0_8534;
  wire                _zz_dataOut_payload_0_8535;
  wire       [7:0]    _zz_dataOut_payload_0_8536;
  wire       [7:0]    _zz_dataOut_payload_0_8537;
  wire                _zz_dataOut_payload_0_8538;
  wire       [7:0]    _zz_dataOut_payload_0_8539;
  wire       [7:0]    _zz_dataOut_payload_0_8540;
  wire                _zz_dataOut_payload_0_8541;
  wire       [7:0]    _zz_dataOut_payload_0_8542;
  wire       [7:0]    _zz_dataOut_payload_0_8543;
  wire                _zz_dataOut_payload_0_8544;
  wire       [7:0]    _zz_dataOut_payload_0_8545;
  wire       [7:0]    _zz_dataOut_payload_0_8546;
  wire                _zz_dataOut_payload_0_8547;
  wire       [7:0]    _zz_dataOut_payload_0_8548;
  wire       [7:0]    _zz_dataOut_payload_0_8549;
  wire                _zz_dataOut_payload_0_8550;
  wire                _zz_dataOut_payload_0_8551;
  reg        [7:0]    _zz_dataOut_payload_0_8552;
  reg        [7:0]    _zz_dataOut_payload_0_8553;
  reg        [7:0]    _zz_dataOut_payload_0_8554;
  reg        [7:0]    _zz_dataOut_payload_0_8555;
  wire                _zz_dataOut_payload_0_8556;
  wire       [7:0]    _zz_dataOut_payload_0_8557;
  wire       [7:0]    _zz_dataOut_payload_0_8558;
  wire                _zz_dataOut_payload_0_8559;
  wire       [7:0]    _zz_dataOut_payload_0_8560;
  wire       [7:0]    _zz_dataOut_payload_0_8561;
  wire                _zz_dataOut_payload_0_8562;
  wire                _zz_dataOut_payload_0_8563;
  reg        [7:0]    _zz_dataOut_payload_0_8564;
  reg        [7:0]    _zz_dataOut_payload_0_8565;
  reg        [7:0]    _zz_dataOut_payload_0_8566;
  reg        [7:0]    _zz_dataOut_payload_0_8567;
  reg        [7:0]    _zz_dataOut_payload_0_8568;
  reg        [7:0]    _zz_dataOut_payload_0_8569;
  reg        [7:0]    _zz_dataOut_payload_0_8570;
  reg        [7:0]    _zz_dataOut_payload_0_8571;
  reg        [7:0]    _zz_dataOut_payload_0_8572;
  reg        [7:0]    _zz_dataOut_payload_0_8573;
  reg        [7:0]    _zz_dataOut_payload_0_8574;
  reg        [7:0]    _zz_dataOut_payload_0_8575;
  reg        [7:0]    _zz_dataOut_payload_0_8576;
  reg        [7:0]    _zz_dataOut_payload_0_8577;
  reg        [7:0]    _zz_dataOut_payload_0_8578;
  reg        [7:0]    _zz_dataOut_payload_0_8579;
  reg        [7:0]    _zz_dataOut_payload_0_8580;
  reg        [7:0]    _zz_dataOut_payload_0_8581;
  reg        [7:0]    _zz_dataOut_payload_0_8582;
  reg        [7:0]    _zz_dataOut_payload_0_8583;
  reg        [7:0]    _zz_dataOut_payload_0_8584;
  reg        [7:0]    _zz_dataOut_payload_0_8585;
  reg        [7:0]    _zz_dataOut_payload_0_8586;
  reg        [7:0]    _zz_dataOut_payload_0_8587;
  reg        [7:0]    _zz_dataOut_payload_0_8588;
  reg        [7:0]    _zz_dataOut_payload_0_8589;
  reg        [7:0]    _zz_dataOut_payload_0_8590;
  reg        [7:0]    _zz_dataOut_payload_0_8591;
  wire                _zz_dataOut_payload_0_8592;
  wire       [7:0]    _zz_dataOut_payload_0_8593;
  wire       [7:0]    _zz_dataOut_payload_0_8594;
  wire                _zz_dataOut_payload_0_8595;
  wire       [7:0]    _zz_dataOut_payload_0_8596;
  wire       [7:0]    _zz_dataOut_payload_0_8597;
  wire                _zz_dataOut_payload_0_8598;
  wire       [7:0]    _zz_dataOut_payload_0_8599;
  wire       [7:0]    _zz_dataOut_payload_0_8600;
  wire                _zz_dataOut_payload_0_8601;
  wire       [7:0]    _zz_dataOut_payload_0_8602;
  wire       [7:0]    _zz_dataOut_payload_0_8603;
  wire                _zz_dataOut_payload_0_8604;
  wire       [7:0]    _zz_dataOut_payload_0_8605;
  wire       [7:0]    _zz_dataOut_payload_0_8606;
  wire                _zz_dataOut_payload_0_8607;
  wire       [7:0]    _zz_dataOut_payload_0_8608;
  wire       [7:0]    _zz_dataOut_payload_0_8609;
  wire                _zz_dataOut_payload_0_8610;
  wire       [7:0]    _zz_dataOut_payload_0_8611;
  wire       [7:0]    _zz_dataOut_payload_0_8612;
  wire                _zz_dataOut_payload_0_8613;
  wire       [7:0]    _zz_dataOut_payload_0_8614;
  wire       [7:0]    _zz_dataOut_payload_0_8615;
  wire                _zz_dataOut_payload_0_8616;
  wire       [7:0]    _zz_dataOut_payload_0_8617;
  wire       [7:0]    _zz_dataOut_payload_0_8618;
  wire                _zz_dataOut_payload_0_8619;
  wire       [7:0]    _zz_dataOut_payload_0_8620;
  wire       [7:0]    _zz_dataOut_payload_0_8621;
  wire                _zz_dataOut_payload_0_8622;
  wire       [7:0]    _zz_dataOut_payload_0_8623;
  wire       [7:0]    _zz_dataOut_payload_0_8624;
  wire                _zz_dataOut_payload_0_8625;
  wire       [7:0]    _zz_dataOut_payload_0_8626;
  wire       [7:0]    _zz_dataOut_payload_0_8627;
  wire                _zz_dataOut_payload_0_8628;
  wire       [7:0]    _zz_dataOut_payload_0_8629;
  wire       [7:0]    _zz_dataOut_payload_0_8630;
  wire                _zz_dataOut_payload_0_8631;
  wire       [7:0]    _zz_dataOut_payload_0_8632;
  wire       [7:0]    _zz_dataOut_payload_0_8633;
  wire                _zz_dataOut_payload_0_8634;
  wire                _zz_dataOut_payload_0_8635;
  reg        [7:0]    _zz_dataOut_payload_0_8636;
  reg        [7:0]    _zz_dataOut_payload_0_8637;
  reg        [7:0]    _zz_dataOut_payload_0_8638;
  reg        [7:0]    _zz_dataOut_payload_0_8639;
  wire                _zz_dataOut_payload_0_8640;
  wire       [7:0]    _zz_dataOut_payload_0_8641;
  wire       [7:0]    _zz_dataOut_payload_0_8642;
  wire                _zz_dataOut_payload_0_8643;
  wire       [7:0]    _zz_dataOut_payload_0_8644;
  wire       [7:0]    _zz_dataOut_payload_0_8645;
  wire                _zz_dataOut_payload_0_8646;
  wire                _zz_dataOut_payload_0_8647;
  reg        [7:0]    _zz_dataOut_payload_0_8648;
  reg        [7:0]    _zz_dataOut_payload_0_8649;
  reg        [7:0]    _zz_dataOut_payload_0_8650;
  reg        [7:0]    _zz_dataOut_payload_0_8651;
  reg        [7:0]    _zz_dataOut_payload_0_8652;
  reg        [7:0]    _zz_dataOut_payload_0_8653;
  reg        [7:0]    _zz_dataOut_payload_0_8654;
  reg        [7:0]    _zz_dataOut_payload_0_8655;
  reg        [7:0]    _zz_dataOut_payload_0_8656;
  reg        [7:0]    _zz_dataOut_payload_0_8657;
  reg        [7:0]    _zz_dataOut_payload_0_8658;
  reg        [7:0]    _zz_dataOut_payload_0_8659;
  wire                _zz_dataOut_payload_0_8660;
  wire       [7:0]    _zz_dataOut_payload_0_8661;
  wire       [7:0]    _zz_dataOut_payload_0_8662;
  wire                _zz_dataOut_payload_0_8663;
  wire       [7:0]    _zz_dataOut_payload_0_8664;
  wire       [7:0]    _zz_dataOut_payload_0_8665;
  wire                _zz_dataOut_payload_0_8666;
  wire       [7:0]    _zz_dataOut_payload_0_8667;
  wire       [7:0]    _zz_dataOut_payload_0_8668;
  wire                _zz_dataOut_payload_0_8669;
  wire       [7:0]    _zz_dataOut_payload_0_8670;
  wire       [7:0]    _zz_dataOut_payload_0_8671;
  wire                _zz_dataOut_payload_0_8672;
  wire       [7:0]    _zz_dataOut_payload_0_8673;
  wire       [7:0]    _zz_dataOut_payload_0_8674;
  wire                _zz_dataOut_payload_0_8675;
  wire       [7:0]    _zz_dataOut_payload_0_8676;
  wire       [7:0]    _zz_dataOut_payload_0_8677;
  wire                _zz_dataOut_payload_0_8678;
  wire                _zz_dataOut_payload_0_8679;
  reg        [7:0]    _zz_dataOut_payload_0_8680;
  reg        [7:0]    _zz_dataOut_payload_0_8681;
  reg        [7:0]    _zz_dataOut_payload_0_8682;
  reg        [7:0]    _zz_dataOut_payload_0_8683;
  wire                _zz_dataOut_payload_0_8684;
  wire       [7:0]    _zz_dataOut_payload_0_8685;
  wire       [7:0]    _zz_dataOut_payload_0_8686;
  wire                _zz_dataOut_payload_0_8687;
  wire       [7:0]    _zz_dataOut_payload_0_8688;
  wire       [7:0]    _zz_dataOut_payload_0_8689;
  wire                _zz_dataOut_payload_0_8690;
  wire                _zz_dataOut_payload_0_8691;
  reg        [7:0]    _zz_dataOut_payload_0_8692;
  reg        [7:0]    _zz_dataOut_payload_0_8693;
  reg        [7:0]    _zz_dataOut_payload_0_8694;
  reg        [7:0]    _zz_dataOut_payload_0_8695;
  reg        [7:0]    _zz_dataOut_payload_0_8696;
  reg        [7:0]    _zz_dataOut_payload_0_8697;
  reg        [7:0]    _zz_dataOut_payload_0_8698;
  reg        [7:0]    _zz_dataOut_payload_0_8699;
  reg        [7:0]    _zz_dataOut_payload_0_8700;
  reg        [7:0]    _zz_dataOut_payload_0_8701;
  reg        [7:0]    _zz_dataOut_payload_0_8702;
  reg        [7:0]    _zz_dataOut_payload_0_8703;
  reg        [7:0]    _zz_dataOut_payload_0_8704;
  reg        [7:0]    _zz_dataOut_payload_0_8705;
  reg        [7:0]    _zz_dataOut_payload_0_8706;
  reg        [7:0]    _zz_dataOut_payload_0_8707;
  reg        [7:0]    _zz_dataOut_payload_0_8708;
  reg        [7:0]    _zz_dataOut_payload_0_8709;
  reg        [7:0]    _zz_dataOut_payload_0_8710;
  reg        [7:0]    _zz_dataOut_payload_0_8711;
  reg        [7:0]    _zz_dataOut_payload_0_8712;
  reg        [7:0]    _zz_dataOut_payload_0_8713;
  reg        [7:0]    _zz_dataOut_payload_0_8714;
  reg        [7:0]    _zz_dataOut_payload_0_8715;
  reg        [7:0]    _zz_dataOut_payload_0_8716;
  reg        [7:0]    _zz_dataOut_payload_0_8717;
  reg        [7:0]    _zz_dataOut_payload_0_8718;
  reg        [7:0]    _zz_dataOut_payload_0_8719;
  reg        [7:0]    _zz_dataOut_payload_0_8720;
  reg        [7:0]    _zz_dataOut_payload_0_8721;
  reg        [7:0]    _zz_dataOut_payload_0_8722;
  reg        [7:0]    _zz_dataOut_payload_0_8723;
  reg        [7:0]    _zz_dataOut_payload_0_8724;
  reg        [7:0]    _zz_dataOut_payload_0_8725;
  reg        [7:0]    _zz_dataOut_payload_0_8726;
  reg        [7:0]    _zz_dataOut_payload_0_8727;
  reg        [7:0]    _zz_dataOut_payload_0_8728;
  reg        [7:0]    _zz_dataOut_payload_0_8729;
  reg        [7:0]    _zz_dataOut_payload_0_8730;
  reg        [7:0]    _zz_dataOut_payload_0_8731;
  reg        [7:0]    _zz_dataOut_payload_0_8732;
  reg        [7:0]    _zz_dataOut_payload_0_8733;
  reg        [7:0]    _zz_dataOut_payload_0_8734;
  reg        [7:0]    _zz_dataOut_payload_0_8735;
  reg        [7:0]    _zz_dataOut_payload_0_8736;
  reg        [7:0]    _zz_dataOut_payload_0_8737;
  reg        [7:0]    _zz_dataOut_payload_0_8738;
  reg        [7:0]    _zz_dataOut_payload_0_8739;
  reg        [7:0]    _zz_dataOut_payload_0_8740;
  reg        [7:0]    _zz_dataOut_payload_0_8741;
  reg        [7:0]    _zz_dataOut_payload_0_8742;
  reg        [7:0]    _zz_dataOut_payload_0_8743;
  reg        [7:0]    _zz_dataOut_payload_0_8744;
  reg        [7:0]    _zz_dataOut_payload_0_8745;
  reg        [7:0]    _zz_dataOut_payload_0_8746;
  reg        [7:0]    _zz_dataOut_payload_0_8747;
  reg        [7:0]    _zz_dataOut_payload_0_8748;
  reg        [7:0]    _zz_dataOut_payload_0_8749;
  reg        [7:0]    _zz_dataOut_payload_0_8750;
  reg        [7:0]    _zz_dataOut_payload_0_8751;
  wire                _zz_dataOut_payload_0_8752;
  wire       [7:0]    _zz_dataOut_payload_0_8753;
  wire       [7:0]    _zz_dataOut_payload_0_8754;
  wire                _zz_dataOut_payload_0_8755;
  wire       [7:0]    _zz_dataOut_payload_0_8756;
  wire       [7:0]    _zz_dataOut_payload_0_8757;
  wire                _zz_dataOut_payload_0_8758;
  wire       [7:0]    _zz_dataOut_payload_0_8759;
  wire       [7:0]    _zz_dataOut_payload_0_8760;
  wire                _zz_dataOut_payload_0_8761;
  wire       [7:0]    _zz_dataOut_payload_0_8762;
  wire       [7:0]    _zz_dataOut_payload_0_8763;
  wire                _zz_dataOut_payload_0_8764;
  wire       [7:0]    _zz_dataOut_payload_0_8765;
  wire       [7:0]    _zz_dataOut_payload_0_8766;
  wire                _zz_dataOut_payload_0_8767;
  wire       [7:0]    _zz_dataOut_payload_0_8768;
  wire       [7:0]    _zz_dataOut_payload_0_8769;
  wire                _zz_dataOut_payload_0_8770;
  wire       [7:0]    _zz_dataOut_payload_0_8771;
  wire       [7:0]    _zz_dataOut_payload_0_8772;
  wire                _zz_dataOut_payload_0_8773;
  wire       [7:0]    _zz_dataOut_payload_0_8774;
  wire       [7:0]    _zz_dataOut_payload_0_8775;
  wire                _zz_dataOut_payload_0_8776;
  wire       [7:0]    _zz_dataOut_payload_0_8777;
  wire       [7:0]    _zz_dataOut_payload_0_8778;
  wire                _zz_dataOut_payload_0_8779;
  wire       [7:0]    _zz_dataOut_payload_0_8780;
  wire       [7:0]    _zz_dataOut_payload_0_8781;
  wire                _zz_dataOut_payload_0_8782;
  wire       [7:0]    _zz_dataOut_payload_0_8783;
  wire       [7:0]    _zz_dataOut_payload_0_8784;
  wire                _zz_dataOut_payload_0_8785;
  wire       [7:0]    _zz_dataOut_payload_0_8786;
  wire       [7:0]    _zz_dataOut_payload_0_8787;
  wire                _zz_dataOut_payload_0_8788;
  wire       [7:0]    _zz_dataOut_payload_0_8789;
  wire       [7:0]    _zz_dataOut_payload_0_8790;
  wire                _zz_dataOut_payload_0_8791;
  wire       [7:0]    _zz_dataOut_payload_0_8792;
  wire       [7:0]    _zz_dataOut_payload_0_8793;
  wire                _zz_dataOut_payload_0_8794;
  wire       [7:0]    _zz_dataOut_payload_0_8795;
  wire       [7:0]    _zz_dataOut_payload_0_8796;
  wire                _zz_dataOut_payload_0_8797;
  wire       [7:0]    _zz_dataOut_payload_0_8798;
  wire       [7:0]    _zz_dataOut_payload_0_8799;
  wire                _zz_dataOut_payload_0_8800;
  wire       [7:0]    _zz_dataOut_payload_0_8801;
  wire       [7:0]    _zz_dataOut_payload_0_8802;
  wire                _zz_dataOut_payload_0_8803;
  wire       [7:0]    _zz_dataOut_payload_0_8804;
  wire       [7:0]    _zz_dataOut_payload_0_8805;
  wire                _zz_dataOut_payload_0_8806;
  wire       [7:0]    _zz_dataOut_payload_0_8807;
  wire       [7:0]    _zz_dataOut_payload_0_8808;
  wire                _zz_dataOut_payload_0_8809;
  wire       [7:0]    _zz_dataOut_payload_0_8810;
  wire       [7:0]    _zz_dataOut_payload_0_8811;
  wire                _zz_dataOut_payload_0_8812;
  wire       [7:0]    _zz_dataOut_payload_0_8813;
  wire       [7:0]    _zz_dataOut_payload_0_8814;
  wire                _zz_dataOut_payload_0_8815;
  wire       [7:0]    _zz_dataOut_payload_0_8816;
  wire       [7:0]    _zz_dataOut_payload_0_8817;
  wire                _zz_dataOut_payload_0_8818;
  wire       [7:0]    _zz_dataOut_payload_0_8819;
  wire       [7:0]    _zz_dataOut_payload_0_8820;
  wire                _zz_dataOut_payload_0_8821;
  wire       [7:0]    _zz_dataOut_payload_0_8822;
  wire       [7:0]    _zz_dataOut_payload_0_8823;
  wire                _zz_dataOut_payload_0_8824;
  wire       [7:0]    _zz_dataOut_payload_0_8825;
  wire       [7:0]    _zz_dataOut_payload_0_8826;
  wire                _zz_dataOut_payload_0_8827;
  wire       [7:0]    _zz_dataOut_payload_0_8828;
  wire       [7:0]    _zz_dataOut_payload_0_8829;
  wire                _zz_dataOut_payload_0_8830;
  wire       [7:0]    _zz_dataOut_payload_0_8831;
  wire       [7:0]    _zz_dataOut_payload_0_8832;
  wire                _zz_dataOut_payload_0_8833;
  wire       [7:0]    _zz_dataOut_payload_0_8834;
  wire       [7:0]    _zz_dataOut_payload_0_8835;
  wire                _zz_dataOut_payload_0_8836;
  wire       [7:0]    _zz_dataOut_payload_0_8837;
  wire       [7:0]    _zz_dataOut_payload_0_8838;
  wire                _zz_dataOut_payload_0_8839;
  wire       [7:0]    _zz_dataOut_payload_0_8840;
  wire       [7:0]    _zz_dataOut_payload_0_8841;
  wire                _zz_dataOut_payload_0_8842;
  wire                _zz_dataOut_payload_0_8843;
  reg        [7:0]    _zz_dataOut_payload_0_8844;
  reg        [7:0]    _zz_dataOut_payload_0_8845;
  reg        [7:0]    _zz_dataOut_payload_0_8846;
  reg        [7:0]    _zz_dataOut_payload_0_8847;
  wire                _zz_dataOut_payload_0_8848;
  wire       [7:0]    _zz_dataOut_payload_0_8849;
  wire       [7:0]    _zz_dataOut_payload_0_8850;
  wire                _zz_dataOut_payload_0_8851;
  wire       [7:0]    _zz_dataOut_payload_0_8852;
  wire       [7:0]    _zz_dataOut_payload_0_8853;
  wire                _zz_dataOut_payload_0_8854;
  wire                _zz_dataOut_payload_0_8855;
  reg        [7:0]    _zz_dataOut_payload_0_8856;
  reg        [7:0]    _zz_dataOut_payload_0_8857;
  reg        [7:0]    _zz_dataOut_payload_0_8858;
  reg        [7:0]    _zz_dataOut_payload_0_8859;
  reg        [7:0]    _zz_dataOut_payload_0_8860;
  reg        [7:0]    _zz_dataOut_payload_0_8861;
  reg        [7:0]    _zz_dataOut_payload_0_8862;
  reg        [7:0]    _zz_dataOut_payload_0_8863;
  reg        [7:0]    _zz_dataOut_payload_0_8864;
  reg        [7:0]    _zz_dataOut_payload_0_8865;
  reg        [7:0]    _zz_dataOut_payload_0_8866;
  reg        [7:0]    _zz_dataOut_payload_0_8867;
  wire                _zz_dataOut_payload_0_8868;
  wire       [7:0]    _zz_dataOut_payload_0_8869;
  wire       [7:0]    _zz_dataOut_payload_0_8870;
  wire                _zz_dataOut_payload_0_8871;
  wire       [7:0]    _zz_dataOut_payload_0_8872;
  wire       [7:0]    _zz_dataOut_payload_0_8873;
  wire                _zz_dataOut_payload_0_8874;
  wire       [7:0]    _zz_dataOut_payload_0_8875;
  wire       [7:0]    _zz_dataOut_payload_0_8876;
  wire                _zz_dataOut_payload_0_8877;
  wire       [7:0]    _zz_dataOut_payload_0_8878;
  wire       [7:0]    _zz_dataOut_payload_0_8879;
  wire                _zz_dataOut_payload_0_8880;
  wire       [7:0]    _zz_dataOut_payload_0_8881;
  wire       [7:0]    _zz_dataOut_payload_0_8882;
  wire                _zz_dataOut_payload_0_8883;
  wire       [7:0]    _zz_dataOut_payload_0_8884;
  wire       [7:0]    _zz_dataOut_payload_0_8885;
  wire                _zz_dataOut_payload_0_8886;
  wire                _zz_dataOut_payload_0_8887;
  reg        [7:0]    _zz_dataOut_payload_0_8888;
  reg        [7:0]    _zz_dataOut_payload_0_8889;
  reg        [7:0]    _zz_dataOut_payload_0_8890;
  reg        [7:0]    _zz_dataOut_payload_0_8891;
  wire                _zz_dataOut_payload_0_8892;
  wire       [7:0]    _zz_dataOut_payload_0_8893;
  wire       [7:0]    _zz_dataOut_payload_0_8894;
  wire                _zz_dataOut_payload_0_8895;
  wire       [7:0]    _zz_dataOut_payload_0_8896;
  wire       [7:0]    _zz_dataOut_payload_0_8897;
  wire                _zz_dataOut_payload_0_8898;
  wire                _zz_dataOut_payload_0_8899;
  reg        [7:0]    _zz_dataOut_payload_0_8900;
  reg        [7:0]    _zz_dataOut_payload_0_8901;
  reg        [7:0]    _zz_dataOut_payload_0_8902;
  reg        [7:0]    _zz_dataOut_payload_0_8903;
  reg        [7:0]    _zz_dataOut_payload_0_8904;
  reg        [7:0]    _zz_dataOut_payload_0_8905;
  reg        [7:0]    _zz_dataOut_payload_0_8906;
  reg        [7:0]    _zz_dataOut_payload_0_8907;
  reg        [7:0]    _zz_dataOut_payload_0_8908;
  reg        [7:0]    _zz_dataOut_payload_0_8909;
  reg        [7:0]    _zz_dataOut_payload_0_8910;
  reg        [7:0]    _zz_dataOut_payload_0_8911;
  reg        [7:0]    _zz_dataOut_payload_0_8912;
  reg        [7:0]    _zz_dataOut_payload_0_8913;
  reg        [7:0]    _zz_dataOut_payload_0_8914;
  reg        [7:0]    _zz_dataOut_payload_0_8915;
  reg        [7:0]    _zz_dataOut_payload_0_8916;
  reg        [7:0]    _zz_dataOut_payload_0_8917;
  reg        [7:0]    _zz_dataOut_payload_0_8918;
  reg        [7:0]    _zz_dataOut_payload_0_8919;
  reg        [7:0]    _zz_dataOut_payload_0_8920;
  reg        [7:0]    _zz_dataOut_payload_0_8921;
  reg        [7:0]    _zz_dataOut_payload_0_8922;
  reg        [7:0]    _zz_dataOut_payload_0_8923;
  reg        [7:0]    _zz_dataOut_payload_0_8924;
  reg        [7:0]    _zz_dataOut_payload_0_8925;
  reg        [7:0]    _zz_dataOut_payload_0_8926;
  reg        [7:0]    _zz_dataOut_payload_0_8927;
  wire                _zz_dataOut_payload_0_8928;
  wire       [7:0]    _zz_dataOut_payload_0_8929;
  wire       [7:0]    _zz_dataOut_payload_0_8930;
  wire                _zz_dataOut_payload_0_8931;
  wire       [7:0]    _zz_dataOut_payload_0_8932;
  wire       [7:0]    _zz_dataOut_payload_0_8933;
  wire                _zz_dataOut_payload_0_8934;
  wire       [7:0]    _zz_dataOut_payload_0_8935;
  wire       [7:0]    _zz_dataOut_payload_0_8936;
  wire                _zz_dataOut_payload_0_8937;
  wire       [7:0]    _zz_dataOut_payload_0_8938;
  wire       [7:0]    _zz_dataOut_payload_0_8939;
  wire                _zz_dataOut_payload_0_8940;
  wire       [7:0]    _zz_dataOut_payload_0_8941;
  wire       [7:0]    _zz_dataOut_payload_0_8942;
  wire                _zz_dataOut_payload_0_8943;
  wire       [7:0]    _zz_dataOut_payload_0_8944;
  wire       [7:0]    _zz_dataOut_payload_0_8945;
  wire                _zz_dataOut_payload_0_8946;
  wire       [7:0]    _zz_dataOut_payload_0_8947;
  wire       [7:0]    _zz_dataOut_payload_0_8948;
  wire                _zz_dataOut_payload_0_8949;
  wire       [7:0]    _zz_dataOut_payload_0_8950;
  wire       [7:0]    _zz_dataOut_payload_0_8951;
  wire                _zz_dataOut_payload_0_8952;
  wire       [7:0]    _zz_dataOut_payload_0_8953;
  wire       [7:0]    _zz_dataOut_payload_0_8954;
  wire                _zz_dataOut_payload_0_8955;
  wire       [7:0]    _zz_dataOut_payload_0_8956;
  wire       [7:0]    _zz_dataOut_payload_0_8957;
  wire                _zz_dataOut_payload_0_8958;
  wire       [7:0]    _zz_dataOut_payload_0_8959;
  wire       [7:0]    _zz_dataOut_payload_0_8960;
  wire                _zz_dataOut_payload_0_8961;
  wire       [7:0]    _zz_dataOut_payload_0_8962;
  wire       [7:0]    _zz_dataOut_payload_0_8963;
  wire                _zz_dataOut_payload_0_8964;
  wire       [7:0]    _zz_dataOut_payload_0_8965;
  wire       [7:0]    _zz_dataOut_payload_0_8966;
  wire                _zz_dataOut_payload_0_8967;
  wire       [7:0]    _zz_dataOut_payload_0_8968;
  wire       [7:0]    _zz_dataOut_payload_0_8969;
  wire                _zz_dataOut_payload_0_8970;
  wire                _zz_dataOut_payload_0_8971;
  reg        [7:0]    _zz_dataOut_payload_0_8972;
  reg        [7:0]    _zz_dataOut_payload_0_8973;
  reg        [7:0]    _zz_dataOut_payload_0_8974;
  reg        [7:0]    _zz_dataOut_payload_0_8975;
  wire                _zz_dataOut_payload_0_8976;
  wire       [7:0]    _zz_dataOut_payload_0_8977;
  wire       [7:0]    _zz_dataOut_payload_0_8978;
  wire                _zz_dataOut_payload_0_8979;
  wire       [7:0]    _zz_dataOut_payload_0_8980;
  wire       [7:0]    _zz_dataOut_payload_0_8981;
  wire                _zz_dataOut_payload_0_8982;
  wire                _zz_dataOut_payload_0_8983;
  reg        [7:0]    _zz_dataOut_payload_0_8984;
  reg        [7:0]    _zz_dataOut_payload_0_8985;
  reg        [7:0]    _zz_dataOut_payload_0_8986;
  reg        [7:0]    _zz_dataOut_payload_0_8987;
  reg        [7:0]    _zz_dataOut_payload_0_8988;
  reg        [7:0]    _zz_dataOut_payload_0_8989;
  reg        [7:0]    _zz_dataOut_payload_0_8990;
  reg        [7:0]    _zz_dataOut_payload_0_8991;
  reg        [7:0]    _zz_dataOut_payload_0_8992;
  reg        [7:0]    _zz_dataOut_payload_0_8993;
  reg        [7:0]    _zz_dataOut_payload_0_8994;
  reg        [7:0]    _zz_dataOut_payload_0_8995;
  wire                _zz_dataOut_payload_0_8996;
  wire       [7:0]    _zz_dataOut_payload_0_8997;
  wire       [7:0]    _zz_dataOut_payload_0_8998;
  wire                _zz_dataOut_payload_0_8999;
  wire       [7:0]    _zz_dataOut_payload_0_9000;
  wire       [7:0]    _zz_dataOut_payload_0_9001;
  wire                _zz_dataOut_payload_0_9002;
  wire       [7:0]    _zz_dataOut_payload_0_9003;
  wire       [7:0]    _zz_dataOut_payload_0_9004;
  wire                _zz_dataOut_payload_0_9005;
  wire       [7:0]    _zz_dataOut_payload_0_9006;
  wire       [7:0]    _zz_dataOut_payload_0_9007;
  wire                _zz_dataOut_payload_0_9008;
  wire       [7:0]    _zz_dataOut_payload_0_9009;
  wire       [7:0]    _zz_dataOut_payload_0_9010;
  wire                _zz_dataOut_payload_0_9011;
  wire       [7:0]    _zz_dataOut_payload_0_9012;
  wire       [7:0]    _zz_dataOut_payload_0_9013;
  wire                _zz_dataOut_payload_0_9014;
  wire                _zz_dataOut_payload_0_9015;
  reg        [7:0]    _zz_dataOut_payload_0_9016;
  reg        [7:0]    _zz_dataOut_payload_0_9017;
  reg        [7:0]    _zz_dataOut_payload_0_9018;
  reg        [7:0]    _zz_dataOut_payload_0_9019;
  wire                _zz_dataOut_payload_0_9020;
  wire       [7:0]    _zz_dataOut_payload_0_9021;
  wire       [7:0]    _zz_dataOut_payload_0_9022;
  wire                _zz_dataOut_payload_0_9023;
  wire       [7:0]    _zz_dataOut_payload_0_9024;
  wire       [7:0]    _zz_dataOut_payload_0_9025;
  wire                _zz_dataOut_payload_0_9026;
  wire                _zz_dataOut_payload_0_9027;
  reg        [7:0]    _zz_dataOut_payload_0_9028;
  reg        [7:0]    _zz_dataOut_payload_0_9029;
  reg        [7:0]    _zz_dataOut_payload_0_9030;
  reg        [7:0]    _zz_dataOut_payload_0_9031;
  reg        [7:0]    _zz_dataOut_payload_0_9032;
  reg        [7:0]    _zz_dataOut_payload_0_9033;
  reg        [7:0]    _zz_dataOut_payload_0_9034;
  reg        [7:0]    _zz_dataOut_payload_0_9035;
  reg        [7:0]    _zz_dataOut_payload_0_9036;
  reg        [7:0]    _zz_dataOut_payload_0_9037;
  reg        [7:0]    _zz_dataOut_payload_0_9038;
  reg        [7:0]    _zz_dataOut_payload_0_9039;
  reg        [7:0]    _zz_dataOut_payload_0_9040;
  reg        [7:0]    _zz_dataOut_payload_0_9041;
  reg        [7:0]    _zz_dataOut_payload_0_9042;
  reg        [7:0]    _zz_dataOut_payload_0_9043;
  reg        [7:0]    _zz_dataOut_payload_0_9044;
  reg        [7:0]    _zz_dataOut_payload_0_9045;
  reg        [7:0]    _zz_dataOut_payload_0_9046;
  reg        [7:0]    _zz_dataOut_payload_0_9047;
  reg        [7:0]    _zz_dataOut_payload_0_9048;
  reg        [7:0]    _zz_dataOut_payload_0_9049;
  reg        [7:0]    _zz_dataOut_payload_0_9050;
  reg        [7:0]    _zz_dataOut_payload_0_9051;
  reg        [7:0]    _zz_dataOut_payload_0_9052;
  reg        [7:0]    _zz_dataOut_payload_0_9053;
  reg        [7:0]    _zz_dataOut_payload_0_9054;
  reg        [7:0]    _zz_dataOut_payload_0_9055;
  reg        [7:0]    _zz_dataOut_payload_0_9056;
  reg        [7:0]    _zz_dataOut_payload_0_9057;
  reg        [7:0]    _zz_dataOut_payload_0_9058;
  reg        [7:0]    _zz_dataOut_payload_0_9059;
  reg        [7:0]    _zz_dataOut_payload_0_9060;
  reg        [7:0]    _zz_dataOut_payload_0_9061;
  reg        [7:0]    _zz_dataOut_payload_0_9062;
  reg        [7:0]    _zz_dataOut_payload_0_9063;
  reg        [7:0]    _zz_dataOut_payload_0_9064;
  reg        [7:0]    _zz_dataOut_payload_0_9065;
  reg        [7:0]    _zz_dataOut_payload_0_9066;
  reg        [7:0]    _zz_dataOut_payload_0_9067;
  reg        [7:0]    _zz_dataOut_payload_0_9068;
  reg        [7:0]    _zz_dataOut_payload_0_9069;
  reg        [7:0]    _zz_dataOut_payload_0_9070;
  reg        [7:0]    _zz_dataOut_payload_0_9071;
  reg        [7:0]    _zz_dataOut_payload_0_9072;
  reg        [7:0]    _zz_dataOut_payload_0_9073;
  reg        [7:0]    _zz_dataOut_payload_0_9074;
  reg        [7:0]    _zz_dataOut_payload_0_9075;
  reg        [7:0]    _zz_dataOut_payload_0_9076;
  reg        [7:0]    _zz_dataOut_payload_0_9077;
  reg        [7:0]    _zz_dataOut_payload_0_9078;
  reg        [7:0]    _zz_dataOut_payload_0_9079;
  reg        [7:0]    _zz_dataOut_payload_0_9080;
  reg        [7:0]    _zz_dataOut_payload_0_9081;
  reg        [7:0]    _zz_dataOut_payload_0_9082;
  reg        [7:0]    _zz_dataOut_payload_0_9083;
  reg        [7:0]    _zz_dataOut_payload_0_9084;
  reg        [7:0]    _zz_dataOut_payload_0_9085;
  reg        [7:0]    _zz_dataOut_payload_0_9086;
  reg        [7:0]    _zz_dataOut_payload_0_9087;
  reg        [7:0]    _zz_dataOut_payload_0_9088;
  reg        [7:0]    _zz_dataOut_payload_0_9089;
  reg        [7:0]    _zz_dataOut_payload_0_9090;
  reg        [7:0]    _zz_dataOut_payload_0_9091;
  reg        [7:0]    _zz_dataOut_payload_0_9092;
  reg        [7:0]    _zz_dataOut_payload_0_9093;
  reg        [7:0]    _zz_dataOut_payload_0_9094;
  reg        [7:0]    _zz_dataOut_payload_0_9095;
  reg        [7:0]    _zz_dataOut_payload_0_9096;
  reg        [7:0]    _zz_dataOut_payload_0_9097;
  reg        [7:0]    _zz_dataOut_payload_0_9098;
  reg        [7:0]    _zz_dataOut_payload_0_9099;
  reg        [7:0]    _zz_dataOut_payload_0_9100;
  reg        [7:0]    _zz_dataOut_payload_0_9101;
  reg        [7:0]    _zz_dataOut_payload_0_9102;
  reg        [7:0]    _zz_dataOut_payload_0_9103;
  reg        [7:0]    _zz_dataOut_payload_0_9104;
  reg        [7:0]    _zz_dataOut_payload_0_9105;
  reg        [7:0]    _zz_dataOut_payload_0_9106;
  reg        [7:0]    _zz_dataOut_payload_0_9107;
  reg        [7:0]    _zz_dataOut_payload_0_9108;
  reg        [7:0]    _zz_dataOut_payload_0_9109;
  reg        [7:0]    _zz_dataOut_payload_0_9110;
  reg        [7:0]    _zz_dataOut_payload_0_9111;
  reg        [7:0]    _zz_dataOut_payload_0_9112;
  reg        [7:0]    _zz_dataOut_payload_0_9113;
  reg        [7:0]    _zz_dataOut_payload_0_9114;
  reg        [7:0]    _zz_dataOut_payload_0_9115;
  reg        [7:0]    _zz_dataOut_payload_0_9116;
  reg        [7:0]    _zz_dataOut_payload_0_9117;
  reg        [7:0]    _zz_dataOut_payload_0_9118;
  reg        [7:0]    _zz_dataOut_payload_0_9119;
  reg        [7:0]    _zz_dataOut_payload_0_9120;
  reg        [7:0]    _zz_dataOut_payload_0_9121;
  reg        [7:0]    _zz_dataOut_payload_0_9122;
  reg        [7:0]    _zz_dataOut_payload_0_9123;
  reg        [7:0]    _zz_dataOut_payload_0_9124;
  reg        [7:0]    _zz_dataOut_payload_0_9125;
  reg        [7:0]    _zz_dataOut_payload_0_9126;
  reg        [7:0]    _zz_dataOut_payload_0_9127;
  reg        [7:0]    _zz_dataOut_payload_0_9128;
  reg        [7:0]    _zz_dataOut_payload_0_9129;
  reg        [7:0]    _zz_dataOut_payload_0_9130;
  reg        [7:0]    _zz_dataOut_payload_0_9131;
  reg        [7:0]    _zz_dataOut_payload_0_9132;
  reg        [7:0]    _zz_dataOut_payload_0_9133;
  reg        [7:0]    _zz_dataOut_payload_0_9134;
  reg        [7:0]    _zz_dataOut_payload_0_9135;
  reg        [7:0]    _zz_dataOut_payload_0_9136;
  reg        [7:0]    _zz_dataOut_payload_0_9137;
  reg        [7:0]    _zz_dataOut_payload_0_9138;
  reg        [7:0]    _zz_dataOut_payload_0_9139;
  reg        [7:0]    _zz_dataOut_payload_0_9140;
  reg        [7:0]    _zz_dataOut_payload_0_9141;
  reg        [7:0]    _zz_dataOut_payload_0_9142;
  reg        [7:0]    _zz_dataOut_payload_0_9143;
  reg        [7:0]    _zz_dataOut_payload_0_9144;
  reg        [7:0]    _zz_dataOut_payload_0_9145;
  reg        [7:0]    _zz_dataOut_payload_0_9146;
  reg        [7:0]    _zz_dataOut_payload_0_9147;
  reg        [7:0]    _zz_dataOut_payload_0_9148;
  reg        [7:0]    _zz_dataOut_payload_0_9149;
  reg        [7:0]    _zz_dataOut_payload_0_9150;
  reg        [7:0]    _zz_dataOut_payload_0_9151;
  wire                _zz_dataOut_payload_0_9152;
  wire       [7:0]    _zz_dataOut_payload_0_9153;
  wire       [7:0]    _zz_dataOut_payload_0_9154;
  wire                _zz_dataOut_payload_0_9155;
  wire       [7:0]    _zz_dataOut_payload_0_9156;
  wire       [7:0]    _zz_dataOut_payload_0_9157;
  wire                _zz_dataOut_payload_0_9158;
  wire       [7:0]    _zz_dataOut_payload_0_9159;
  wire       [7:0]    _zz_dataOut_payload_0_9160;
  wire                _zz_dataOut_payload_0_9161;
  wire       [7:0]    _zz_dataOut_payload_0_9162;
  wire       [7:0]    _zz_dataOut_payload_0_9163;
  wire                _zz_dataOut_payload_0_9164;
  wire       [7:0]    _zz_dataOut_payload_0_9165;
  wire       [7:0]    _zz_dataOut_payload_0_9166;
  wire                _zz_dataOut_payload_0_9167;
  wire       [7:0]    _zz_dataOut_payload_0_9168;
  wire       [7:0]    _zz_dataOut_payload_0_9169;
  wire                _zz_dataOut_payload_0_9170;
  wire       [7:0]    _zz_dataOut_payload_0_9171;
  wire       [7:0]    _zz_dataOut_payload_0_9172;
  wire                _zz_dataOut_payload_0_9173;
  wire       [7:0]    _zz_dataOut_payload_0_9174;
  wire       [7:0]    _zz_dataOut_payload_0_9175;
  wire                _zz_dataOut_payload_0_9176;
  wire       [7:0]    _zz_dataOut_payload_0_9177;
  wire       [7:0]    _zz_dataOut_payload_0_9178;
  wire                _zz_dataOut_payload_0_9179;
  wire       [7:0]    _zz_dataOut_payload_0_9180;
  wire       [7:0]    _zz_dataOut_payload_0_9181;
  wire                _zz_dataOut_payload_0_9182;
  wire       [7:0]    _zz_dataOut_payload_0_9183;
  wire       [7:0]    _zz_dataOut_payload_0_9184;
  wire                _zz_dataOut_payload_0_9185;
  wire       [7:0]    _zz_dataOut_payload_0_9186;
  wire       [7:0]    _zz_dataOut_payload_0_9187;
  wire                _zz_dataOut_payload_0_9188;
  wire       [7:0]    _zz_dataOut_payload_0_9189;
  wire       [7:0]    _zz_dataOut_payload_0_9190;
  wire                _zz_dataOut_payload_0_9191;
  wire       [7:0]    _zz_dataOut_payload_0_9192;
  wire       [7:0]    _zz_dataOut_payload_0_9193;
  wire                _zz_dataOut_payload_0_9194;
  wire       [7:0]    _zz_dataOut_payload_0_9195;
  wire       [7:0]    _zz_dataOut_payload_0_9196;
  wire                _zz_dataOut_payload_0_9197;
  wire       [7:0]    _zz_dataOut_payload_0_9198;
  wire       [7:0]    _zz_dataOut_payload_0_9199;
  wire                _zz_dataOut_payload_0_9200;
  wire       [7:0]    _zz_dataOut_payload_0_9201;
  wire       [7:0]    _zz_dataOut_payload_0_9202;
  wire                _zz_dataOut_payload_0_9203;
  wire       [7:0]    _zz_dataOut_payload_0_9204;
  wire       [7:0]    _zz_dataOut_payload_0_9205;
  wire                _zz_dataOut_payload_0_9206;
  wire       [7:0]    _zz_dataOut_payload_0_9207;
  wire       [7:0]    _zz_dataOut_payload_0_9208;
  wire                _zz_dataOut_payload_0_9209;
  wire       [7:0]    _zz_dataOut_payload_0_9210;
  wire       [7:0]    _zz_dataOut_payload_0_9211;
  wire                _zz_dataOut_payload_0_9212;
  wire       [7:0]    _zz_dataOut_payload_0_9213;
  wire       [7:0]    _zz_dataOut_payload_0_9214;
  wire                _zz_dataOut_payload_0_9215;
  wire       [7:0]    _zz_dataOut_payload_0_9216;
  wire       [7:0]    _zz_dataOut_payload_0_9217;
  wire                _zz_dataOut_payload_0_9218;
  wire       [7:0]    _zz_dataOut_payload_0_9219;
  wire       [7:0]    _zz_dataOut_payload_0_9220;
  wire                _zz_dataOut_payload_0_9221;
  wire       [7:0]    _zz_dataOut_payload_0_9222;
  wire       [7:0]    _zz_dataOut_payload_0_9223;
  wire                _zz_dataOut_payload_0_9224;
  wire       [7:0]    _zz_dataOut_payload_0_9225;
  wire       [7:0]    _zz_dataOut_payload_0_9226;
  wire                _zz_dataOut_payload_0_9227;
  wire       [7:0]    _zz_dataOut_payload_0_9228;
  wire       [7:0]    _zz_dataOut_payload_0_9229;
  wire                _zz_dataOut_payload_0_9230;
  wire       [7:0]    _zz_dataOut_payload_0_9231;
  wire       [7:0]    _zz_dataOut_payload_0_9232;
  wire                _zz_dataOut_payload_0_9233;
  wire       [7:0]    _zz_dataOut_payload_0_9234;
  wire       [7:0]    _zz_dataOut_payload_0_9235;
  wire                _zz_dataOut_payload_0_9236;
  wire       [7:0]    _zz_dataOut_payload_0_9237;
  wire       [7:0]    _zz_dataOut_payload_0_9238;
  wire                _zz_dataOut_payload_0_9239;
  wire       [7:0]    _zz_dataOut_payload_0_9240;
  wire       [7:0]    _zz_dataOut_payload_0_9241;
  wire                _zz_dataOut_payload_0_9242;
  wire       [7:0]    _zz_dataOut_payload_0_9243;
  wire       [7:0]    _zz_dataOut_payload_0_9244;
  wire                _zz_dataOut_payload_0_9245;
  wire       [7:0]    _zz_dataOut_payload_0_9246;
  wire       [7:0]    _zz_dataOut_payload_0_9247;
  wire                _zz_dataOut_payload_0_9248;
  wire       [7:0]    _zz_dataOut_payload_0_9249;
  wire       [7:0]    _zz_dataOut_payload_0_9250;
  wire                _zz_dataOut_payload_0_9251;
  wire       [7:0]    _zz_dataOut_payload_0_9252;
  wire       [7:0]    _zz_dataOut_payload_0_9253;
  wire                _zz_dataOut_payload_0_9254;
  wire       [7:0]    _zz_dataOut_payload_0_9255;
  wire       [7:0]    _zz_dataOut_payload_0_9256;
  wire                _zz_dataOut_payload_0_9257;
  wire       [7:0]    _zz_dataOut_payload_0_9258;
  wire       [7:0]    _zz_dataOut_payload_0_9259;
  wire                _zz_dataOut_payload_0_9260;
  wire       [7:0]    _zz_dataOut_payload_0_9261;
  wire       [7:0]    _zz_dataOut_payload_0_9262;
  wire                _zz_dataOut_payload_0_9263;
  wire       [7:0]    _zz_dataOut_payload_0_9264;
  wire       [7:0]    _zz_dataOut_payload_0_9265;
  wire                _zz_dataOut_payload_0_9266;
  wire       [7:0]    _zz_dataOut_payload_0_9267;
  wire       [7:0]    _zz_dataOut_payload_0_9268;
  wire                _zz_dataOut_payload_0_9269;
  wire       [7:0]    _zz_dataOut_payload_0_9270;
  wire       [7:0]    _zz_dataOut_payload_0_9271;
  wire                _zz_dataOut_payload_0_9272;
  wire       [7:0]    _zz_dataOut_payload_0_9273;
  wire       [7:0]    _zz_dataOut_payload_0_9274;
  wire                _zz_dataOut_payload_0_9275;
  wire       [7:0]    _zz_dataOut_payload_0_9276;
  wire       [7:0]    _zz_dataOut_payload_0_9277;
  wire                _zz_dataOut_payload_0_9278;
  wire       [7:0]    _zz_dataOut_payload_0_9279;
  wire       [7:0]    _zz_dataOut_payload_0_9280;
  wire                _zz_dataOut_payload_0_9281;
  wire       [7:0]    _zz_dataOut_payload_0_9282;
  wire       [7:0]    _zz_dataOut_payload_0_9283;
  wire                _zz_dataOut_payload_0_9284;
  wire       [7:0]    _zz_dataOut_payload_0_9285;
  wire       [7:0]    _zz_dataOut_payload_0_9286;
  wire                _zz_dataOut_payload_0_9287;
  wire       [7:0]    _zz_dataOut_payload_0_9288;
  wire       [7:0]    _zz_dataOut_payload_0_9289;
  wire                _zz_dataOut_payload_0_9290;
  wire       [7:0]    _zz_dataOut_payload_0_9291;
  wire       [7:0]    _zz_dataOut_payload_0_9292;
  wire                _zz_dataOut_payload_0_9293;
  wire       [7:0]    _zz_dataOut_payload_0_9294;
  wire       [7:0]    _zz_dataOut_payload_0_9295;
  wire                _zz_dataOut_payload_0_9296;
  wire       [7:0]    _zz_dataOut_payload_0_9297;
  wire       [7:0]    _zz_dataOut_payload_0_9298;
  wire                _zz_dataOut_payload_0_9299;
  wire       [7:0]    _zz_dataOut_payload_0_9300;
  wire       [7:0]    _zz_dataOut_payload_0_9301;
  wire                _zz_dataOut_payload_0_9302;
  wire       [7:0]    _zz_dataOut_payload_0_9303;
  wire       [7:0]    _zz_dataOut_payload_0_9304;
  wire                _zz_dataOut_payload_0_9305;
  wire       [7:0]    _zz_dataOut_payload_0_9306;
  wire       [7:0]    _zz_dataOut_payload_0_9307;
  wire                _zz_dataOut_payload_0_9308;
  wire       [7:0]    _zz_dataOut_payload_0_9309;
  wire       [7:0]    _zz_dataOut_payload_0_9310;
  wire                _zz_dataOut_payload_0_9311;
  wire       [7:0]    _zz_dataOut_payload_0_9312;
  wire       [7:0]    _zz_dataOut_payload_0_9313;
  wire                _zz_dataOut_payload_0_9314;
  wire       [7:0]    _zz_dataOut_payload_0_9315;
  wire       [7:0]    _zz_dataOut_payload_0_9316;
  wire                _zz_dataOut_payload_0_9317;
  wire       [7:0]    _zz_dataOut_payload_0_9318;
  wire       [7:0]    _zz_dataOut_payload_0_9319;
  wire                _zz_dataOut_payload_0_9320;
  wire       [7:0]    _zz_dataOut_payload_0_9321;
  wire       [7:0]    _zz_dataOut_payload_0_9322;
  wire                _zz_dataOut_payload_0_9323;
  wire       [7:0]    _zz_dataOut_payload_0_9324;
  wire       [7:0]    _zz_dataOut_payload_0_9325;
  wire                _zz_dataOut_payload_0_9326;
  wire       [7:0]    _zz_dataOut_payload_0_9327;
  wire       [7:0]    _zz_dataOut_payload_0_9328;
  wire                _zz_dataOut_payload_0_9329;
  wire       [7:0]    _zz_dataOut_payload_0_9330;
  wire       [7:0]    _zz_dataOut_payload_0_9331;
  wire                _zz_dataOut_payload_0_9332;
  wire       [7:0]    _zz_dataOut_payload_0_9333;
  wire       [7:0]    _zz_dataOut_payload_0_9334;
  wire                _zz_dataOut_payload_0_9335;
  wire       [7:0]    _zz_dataOut_payload_0_9336;
  wire       [7:0]    _zz_dataOut_payload_0_9337;
  wire                _zz_dataOut_payload_0_9338;
  wire                _zz_dataOut_payload_0_9339;
  reg        [7:0]    _zz_dataOut_payload_0_9340;
  reg        [7:0]    _zz_dataOut_payload_0_9341;
  reg        [7:0]    _zz_dataOut_payload_0_9342;
  reg        [7:0]    _zz_dataOut_payload_0_9343;
  wire                _zz_dataOut_payload_0_9344;
  wire       [7:0]    _zz_dataOut_payload_0_9345;
  wire       [7:0]    _zz_dataOut_payload_0_9346;
  wire                _zz_dataOut_payload_0_9347;
  wire       [7:0]    _zz_dataOut_payload_0_9348;
  wire       [7:0]    _zz_dataOut_payload_0_9349;
  wire                _zz_dataOut_payload_0_9350;
  wire                _zz_dataOut_payload_0_9351;
  reg        [7:0]    _zz_dataOut_payload_0_9352;
  reg        [7:0]    _zz_dataOut_payload_0_9353;
  reg        [7:0]    _zz_dataOut_payload_0_9354;
  reg        [7:0]    _zz_dataOut_payload_0_9355;
  reg        [7:0]    _zz_dataOut_payload_0_9356;
  reg        [7:0]    _zz_dataOut_payload_0_9357;
  reg        [7:0]    _zz_dataOut_payload_0_9358;
  reg        [7:0]    _zz_dataOut_payload_0_9359;
  reg        [7:0]    _zz_dataOut_payload_0_9360;
  reg        [7:0]    _zz_dataOut_payload_0_9361;
  reg        [7:0]    _zz_dataOut_payload_0_9362;
  reg        [7:0]    _zz_dataOut_payload_0_9363;
  wire                _zz_dataOut_payload_0_9364;
  wire       [7:0]    _zz_dataOut_payload_0_9365;
  wire       [7:0]    _zz_dataOut_payload_0_9366;
  wire                _zz_dataOut_payload_0_9367;
  wire       [7:0]    _zz_dataOut_payload_0_9368;
  wire       [7:0]    _zz_dataOut_payload_0_9369;
  wire                _zz_dataOut_payload_0_9370;
  wire       [7:0]    _zz_dataOut_payload_0_9371;
  wire       [7:0]    _zz_dataOut_payload_0_9372;
  wire                _zz_dataOut_payload_0_9373;
  wire       [7:0]    _zz_dataOut_payload_0_9374;
  wire       [7:0]    _zz_dataOut_payload_0_9375;
  wire                _zz_dataOut_payload_0_9376;
  wire       [7:0]    _zz_dataOut_payload_0_9377;
  wire       [7:0]    _zz_dataOut_payload_0_9378;
  wire                _zz_dataOut_payload_0_9379;
  wire       [7:0]    _zz_dataOut_payload_0_9380;
  wire       [7:0]    _zz_dataOut_payload_0_9381;
  wire                _zz_dataOut_payload_0_9382;
  wire                _zz_dataOut_payload_0_9383;
  reg        [7:0]    _zz_dataOut_payload_0_9384;
  reg        [7:0]    _zz_dataOut_payload_0_9385;
  reg        [7:0]    _zz_dataOut_payload_0_9386;
  reg        [7:0]    _zz_dataOut_payload_0_9387;
  wire                _zz_dataOut_payload_0_9388;
  wire       [7:0]    _zz_dataOut_payload_0_9389;
  wire       [7:0]    _zz_dataOut_payload_0_9390;
  wire                _zz_dataOut_payload_0_9391;
  wire       [7:0]    _zz_dataOut_payload_0_9392;
  wire       [7:0]    _zz_dataOut_payload_0_9393;
  wire                _zz_dataOut_payload_0_9394;
  wire                _zz_dataOut_payload_0_9395;
  reg        [7:0]    _zz_dataOut_payload_0_9396;
  reg        [7:0]    _zz_dataOut_payload_0_9397;
  reg        [7:0]    _zz_dataOut_payload_0_9398;
  reg        [7:0]    _zz_dataOut_payload_0_9399;
  reg        [7:0]    _zz_dataOut_payload_0_9400;
  reg        [7:0]    _zz_dataOut_payload_0_9401;
  reg        [7:0]    _zz_dataOut_payload_0_9402;
  reg        [7:0]    _zz_dataOut_payload_0_9403;
  reg        [7:0]    _zz_dataOut_payload_0_9404;
  reg        [7:0]    _zz_dataOut_payload_0_9405;
  reg        [7:0]    _zz_dataOut_payload_0_9406;
  reg        [7:0]    _zz_dataOut_payload_0_9407;
  reg        [7:0]    _zz_dataOut_payload_0_9408;
  reg        [7:0]    _zz_dataOut_payload_0_9409;
  reg        [7:0]    _zz_dataOut_payload_0_9410;
  reg        [7:0]    _zz_dataOut_payload_0_9411;
  reg        [7:0]    _zz_dataOut_payload_0_9412;
  reg        [7:0]    _zz_dataOut_payload_0_9413;
  reg        [7:0]    _zz_dataOut_payload_0_9414;
  reg        [7:0]    _zz_dataOut_payload_0_9415;
  reg        [7:0]    _zz_dataOut_payload_0_9416;
  reg        [7:0]    _zz_dataOut_payload_0_9417;
  reg        [7:0]    _zz_dataOut_payload_0_9418;
  reg        [7:0]    _zz_dataOut_payload_0_9419;
  reg        [7:0]    _zz_dataOut_payload_0_9420;
  reg        [7:0]    _zz_dataOut_payload_0_9421;
  reg        [7:0]    _zz_dataOut_payload_0_9422;
  reg        [7:0]    _zz_dataOut_payload_0_9423;
  wire                _zz_dataOut_payload_0_9424;
  wire       [7:0]    _zz_dataOut_payload_0_9425;
  wire       [7:0]    _zz_dataOut_payload_0_9426;
  wire                _zz_dataOut_payload_0_9427;
  wire       [7:0]    _zz_dataOut_payload_0_9428;
  wire       [7:0]    _zz_dataOut_payload_0_9429;
  wire                _zz_dataOut_payload_0_9430;
  wire       [7:0]    _zz_dataOut_payload_0_9431;
  wire       [7:0]    _zz_dataOut_payload_0_9432;
  wire                _zz_dataOut_payload_0_9433;
  wire       [7:0]    _zz_dataOut_payload_0_9434;
  wire       [7:0]    _zz_dataOut_payload_0_9435;
  wire                _zz_dataOut_payload_0_9436;
  wire       [7:0]    _zz_dataOut_payload_0_9437;
  wire       [7:0]    _zz_dataOut_payload_0_9438;
  wire                _zz_dataOut_payload_0_9439;
  wire       [7:0]    _zz_dataOut_payload_0_9440;
  wire       [7:0]    _zz_dataOut_payload_0_9441;
  wire                _zz_dataOut_payload_0_9442;
  wire       [7:0]    _zz_dataOut_payload_0_9443;
  wire       [7:0]    _zz_dataOut_payload_0_9444;
  wire                _zz_dataOut_payload_0_9445;
  wire       [7:0]    _zz_dataOut_payload_0_9446;
  wire       [7:0]    _zz_dataOut_payload_0_9447;
  wire                _zz_dataOut_payload_0_9448;
  wire       [7:0]    _zz_dataOut_payload_0_9449;
  wire       [7:0]    _zz_dataOut_payload_0_9450;
  wire                _zz_dataOut_payload_0_9451;
  wire       [7:0]    _zz_dataOut_payload_0_9452;
  wire       [7:0]    _zz_dataOut_payload_0_9453;
  wire                _zz_dataOut_payload_0_9454;
  wire       [7:0]    _zz_dataOut_payload_0_9455;
  wire       [7:0]    _zz_dataOut_payload_0_9456;
  wire                _zz_dataOut_payload_0_9457;
  wire       [7:0]    _zz_dataOut_payload_0_9458;
  wire       [7:0]    _zz_dataOut_payload_0_9459;
  wire                _zz_dataOut_payload_0_9460;
  wire       [7:0]    _zz_dataOut_payload_0_9461;
  wire       [7:0]    _zz_dataOut_payload_0_9462;
  wire                _zz_dataOut_payload_0_9463;
  wire       [7:0]    _zz_dataOut_payload_0_9464;
  wire       [7:0]    _zz_dataOut_payload_0_9465;
  wire                _zz_dataOut_payload_0_9466;
  wire                _zz_dataOut_payload_0_9467;
  reg        [7:0]    _zz_dataOut_payload_0_9468;
  reg        [7:0]    _zz_dataOut_payload_0_9469;
  reg        [7:0]    _zz_dataOut_payload_0_9470;
  reg        [7:0]    _zz_dataOut_payload_0_9471;
  wire                _zz_dataOut_payload_0_9472;
  wire       [7:0]    _zz_dataOut_payload_0_9473;
  wire       [7:0]    _zz_dataOut_payload_0_9474;
  wire                _zz_dataOut_payload_0_9475;
  wire       [7:0]    _zz_dataOut_payload_0_9476;
  wire       [7:0]    _zz_dataOut_payload_0_9477;
  wire                _zz_dataOut_payload_0_9478;
  wire                _zz_dataOut_payload_0_9479;
  reg        [7:0]    _zz_dataOut_payload_0_9480;
  reg        [7:0]    _zz_dataOut_payload_0_9481;
  reg        [7:0]    _zz_dataOut_payload_0_9482;
  reg        [7:0]    _zz_dataOut_payload_0_9483;
  reg        [7:0]    _zz_dataOut_payload_0_9484;
  reg        [7:0]    _zz_dataOut_payload_0_9485;
  reg        [7:0]    _zz_dataOut_payload_0_9486;
  reg        [7:0]    _zz_dataOut_payload_0_9487;
  reg        [7:0]    _zz_dataOut_payload_0_9488;
  reg        [7:0]    _zz_dataOut_payload_0_9489;
  reg        [7:0]    _zz_dataOut_payload_0_9490;
  reg        [7:0]    _zz_dataOut_payload_0_9491;
  wire                _zz_dataOut_payload_0_9492;
  wire       [7:0]    _zz_dataOut_payload_0_9493;
  wire       [7:0]    _zz_dataOut_payload_0_9494;
  wire                _zz_dataOut_payload_0_9495;
  wire       [7:0]    _zz_dataOut_payload_0_9496;
  wire       [7:0]    _zz_dataOut_payload_0_9497;
  wire                _zz_dataOut_payload_0_9498;
  wire       [7:0]    _zz_dataOut_payload_0_9499;
  wire       [7:0]    _zz_dataOut_payload_0_9500;
  wire                _zz_dataOut_payload_0_9501;
  wire       [7:0]    _zz_dataOut_payload_0_9502;
  wire       [7:0]    _zz_dataOut_payload_0_9503;
  wire                _zz_dataOut_payload_0_9504;
  wire       [7:0]    _zz_dataOut_payload_0_9505;
  wire       [7:0]    _zz_dataOut_payload_0_9506;
  wire                _zz_dataOut_payload_0_9507;
  wire       [7:0]    _zz_dataOut_payload_0_9508;
  wire       [7:0]    _zz_dataOut_payload_0_9509;
  wire                _zz_dataOut_payload_0_9510;
  wire                _zz_dataOut_payload_0_9511;
  reg        [7:0]    _zz_dataOut_payload_0_9512;
  reg        [7:0]    _zz_dataOut_payload_0_9513;
  reg        [7:0]    _zz_dataOut_payload_0_9514;
  reg        [7:0]    _zz_dataOut_payload_0_9515;
  wire                _zz_dataOut_payload_0_9516;
  wire       [7:0]    _zz_dataOut_payload_0_9517;
  wire       [7:0]    _zz_dataOut_payload_0_9518;
  wire                _zz_dataOut_payload_0_9519;
  wire       [7:0]    _zz_dataOut_payload_0_9520;
  wire       [7:0]    _zz_dataOut_payload_0_9521;
  wire                _zz_dataOut_payload_0_9522;
  wire                _zz_dataOut_payload_0_9523;
  reg        [7:0]    _zz_dataOut_payload_0_9524;
  reg        [7:0]    _zz_dataOut_payload_0_9525;
  reg        [7:0]    _zz_dataOut_payload_0_9526;
  reg        [7:0]    _zz_dataOut_payload_0_9527;
  reg        [7:0]    _zz_dataOut_payload_0_9528;
  reg        [7:0]    _zz_dataOut_payload_0_9529;
  reg        [7:0]    _zz_dataOut_payload_0_9530;
  reg        [7:0]    _zz_dataOut_payload_0_9531;
  reg        [7:0]    _zz_dataOut_payload_0_9532;
  reg        [7:0]    _zz_dataOut_payload_0_9533;
  reg        [7:0]    _zz_dataOut_payload_0_9534;
  reg        [7:0]    _zz_dataOut_payload_0_9535;
  reg        [7:0]    _zz_dataOut_payload_0_9536;
  reg        [7:0]    _zz_dataOut_payload_0_9537;
  reg        [7:0]    _zz_dataOut_payload_0_9538;
  reg        [7:0]    _zz_dataOut_payload_0_9539;
  reg        [7:0]    _zz_dataOut_payload_0_9540;
  reg        [7:0]    _zz_dataOut_payload_0_9541;
  reg        [7:0]    _zz_dataOut_payload_0_9542;
  reg        [7:0]    _zz_dataOut_payload_0_9543;
  reg        [7:0]    _zz_dataOut_payload_0_9544;
  reg        [7:0]    _zz_dataOut_payload_0_9545;
  reg        [7:0]    _zz_dataOut_payload_0_9546;
  reg        [7:0]    _zz_dataOut_payload_0_9547;
  reg        [7:0]    _zz_dataOut_payload_0_9548;
  reg        [7:0]    _zz_dataOut_payload_0_9549;
  reg        [7:0]    _zz_dataOut_payload_0_9550;
  reg        [7:0]    _zz_dataOut_payload_0_9551;
  reg        [7:0]    _zz_dataOut_payload_0_9552;
  reg        [7:0]    _zz_dataOut_payload_0_9553;
  reg        [7:0]    _zz_dataOut_payload_0_9554;
  reg        [7:0]    _zz_dataOut_payload_0_9555;
  reg        [7:0]    _zz_dataOut_payload_0_9556;
  reg        [7:0]    _zz_dataOut_payload_0_9557;
  reg        [7:0]    _zz_dataOut_payload_0_9558;
  reg        [7:0]    _zz_dataOut_payload_0_9559;
  reg        [7:0]    _zz_dataOut_payload_0_9560;
  reg        [7:0]    _zz_dataOut_payload_0_9561;
  reg        [7:0]    _zz_dataOut_payload_0_9562;
  reg        [7:0]    _zz_dataOut_payload_0_9563;
  reg        [7:0]    _zz_dataOut_payload_0_9564;
  reg        [7:0]    _zz_dataOut_payload_0_9565;
  reg        [7:0]    _zz_dataOut_payload_0_9566;
  reg        [7:0]    _zz_dataOut_payload_0_9567;
  reg        [7:0]    _zz_dataOut_payload_0_9568;
  reg        [7:0]    _zz_dataOut_payload_0_9569;
  reg        [7:0]    _zz_dataOut_payload_0_9570;
  reg        [7:0]    _zz_dataOut_payload_0_9571;
  reg        [7:0]    _zz_dataOut_payload_0_9572;
  reg        [7:0]    _zz_dataOut_payload_0_9573;
  reg        [7:0]    _zz_dataOut_payload_0_9574;
  reg        [7:0]    _zz_dataOut_payload_0_9575;
  reg        [7:0]    _zz_dataOut_payload_0_9576;
  reg        [7:0]    _zz_dataOut_payload_0_9577;
  reg        [7:0]    _zz_dataOut_payload_0_9578;
  reg        [7:0]    _zz_dataOut_payload_0_9579;
  reg        [7:0]    _zz_dataOut_payload_0_9580;
  reg        [7:0]    _zz_dataOut_payload_0_9581;
  reg        [7:0]    _zz_dataOut_payload_0_9582;
  reg        [7:0]    _zz_dataOut_payload_0_9583;
  wire                _zz_dataOut_payload_0_9584;
  wire       [7:0]    _zz_dataOut_payload_0_9585;
  wire       [7:0]    _zz_dataOut_payload_0_9586;
  wire                _zz_dataOut_payload_0_9587;
  wire       [7:0]    _zz_dataOut_payload_0_9588;
  wire       [7:0]    _zz_dataOut_payload_0_9589;
  wire                _zz_dataOut_payload_0_9590;
  wire       [7:0]    _zz_dataOut_payload_0_9591;
  wire       [7:0]    _zz_dataOut_payload_0_9592;
  wire                _zz_dataOut_payload_0_9593;
  wire       [7:0]    _zz_dataOut_payload_0_9594;
  wire       [7:0]    _zz_dataOut_payload_0_9595;
  wire                _zz_dataOut_payload_0_9596;
  wire       [7:0]    _zz_dataOut_payload_0_9597;
  wire       [7:0]    _zz_dataOut_payload_0_9598;
  wire                _zz_dataOut_payload_0_9599;
  wire       [7:0]    _zz_dataOut_payload_0_9600;
  wire       [7:0]    _zz_dataOut_payload_0_9601;
  wire                _zz_dataOut_payload_0_9602;
  wire       [7:0]    _zz_dataOut_payload_0_9603;
  wire       [7:0]    _zz_dataOut_payload_0_9604;
  wire                _zz_dataOut_payload_0_9605;
  wire       [7:0]    _zz_dataOut_payload_0_9606;
  wire       [7:0]    _zz_dataOut_payload_0_9607;
  wire                _zz_dataOut_payload_0_9608;
  wire       [7:0]    _zz_dataOut_payload_0_9609;
  wire       [7:0]    _zz_dataOut_payload_0_9610;
  wire                _zz_dataOut_payload_0_9611;
  wire       [7:0]    _zz_dataOut_payload_0_9612;
  wire       [7:0]    _zz_dataOut_payload_0_9613;
  wire                _zz_dataOut_payload_0_9614;
  wire       [7:0]    _zz_dataOut_payload_0_9615;
  wire       [7:0]    _zz_dataOut_payload_0_9616;
  wire                _zz_dataOut_payload_0_9617;
  wire       [7:0]    _zz_dataOut_payload_0_9618;
  wire       [7:0]    _zz_dataOut_payload_0_9619;
  wire                _zz_dataOut_payload_0_9620;
  wire       [7:0]    _zz_dataOut_payload_0_9621;
  wire       [7:0]    _zz_dataOut_payload_0_9622;
  wire                _zz_dataOut_payload_0_9623;
  wire       [7:0]    _zz_dataOut_payload_0_9624;
  wire       [7:0]    _zz_dataOut_payload_0_9625;
  wire                _zz_dataOut_payload_0_9626;
  wire       [7:0]    _zz_dataOut_payload_0_9627;
  wire       [7:0]    _zz_dataOut_payload_0_9628;
  wire                _zz_dataOut_payload_0_9629;
  wire       [7:0]    _zz_dataOut_payload_0_9630;
  wire       [7:0]    _zz_dataOut_payload_0_9631;
  wire                _zz_dataOut_payload_0_9632;
  wire       [7:0]    _zz_dataOut_payload_0_9633;
  wire       [7:0]    _zz_dataOut_payload_0_9634;
  wire                _zz_dataOut_payload_0_9635;
  wire       [7:0]    _zz_dataOut_payload_0_9636;
  wire       [7:0]    _zz_dataOut_payload_0_9637;
  wire                _zz_dataOut_payload_0_9638;
  wire       [7:0]    _zz_dataOut_payload_0_9639;
  wire       [7:0]    _zz_dataOut_payload_0_9640;
  wire                _zz_dataOut_payload_0_9641;
  wire       [7:0]    _zz_dataOut_payload_0_9642;
  wire       [7:0]    _zz_dataOut_payload_0_9643;
  wire                _zz_dataOut_payload_0_9644;
  wire       [7:0]    _zz_dataOut_payload_0_9645;
  wire       [7:0]    _zz_dataOut_payload_0_9646;
  wire                _zz_dataOut_payload_0_9647;
  wire       [7:0]    _zz_dataOut_payload_0_9648;
  wire       [7:0]    _zz_dataOut_payload_0_9649;
  wire                _zz_dataOut_payload_0_9650;
  wire       [7:0]    _zz_dataOut_payload_0_9651;
  wire       [7:0]    _zz_dataOut_payload_0_9652;
  wire                _zz_dataOut_payload_0_9653;
  wire       [7:0]    _zz_dataOut_payload_0_9654;
  wire       [7:0]    _zz_dataOut_payload_0_9655;
  wire                _zz_dataOut_payload_0_9656;
  wire       [7:0]    _zz_dataOut_payload_0_9657;
  wire       [7:0]    _zz_dataOut_payload_0_9658;
  wire                _zz_dataOut_payload_0_9659;
  wire       [7:0]    _zz_dataOut_payload_0_9660;
  wire       [7:0]    _zz_dataOut_payload_0_9661;
  wire                _zz_dataOut_payload_0_9662;
  wire       [7:0]    _zz_dataOut_payload_0_9663;
  wire       [7:0]    _zz_dataOut_payload_0_9664;
  wire                _zz_dataOut_payload_0_9665;
  wire       [7:0]    _zz_dataOut_payload_0_9666;
  wire       [7:0]    _zz_dataOut_payload_0_9667;
  wire                _zz_dataOut_payload_0_9668;
  wire       [7:0]    _zz_dataOut_payload_0_9669;
  wire       [7:0]    _zz_dataOut_payload_0_9670;
  wire                _zz_dataOut_payload_0_9671;
  wire       [7:0]    _zz_dataOut_payload_0_9672;
  wire       [7:0]    _zz_dataOut_payload_0_9673;
  wire                _zz_dataOut_payload_0_9674;
  wire                _zz_dataOut_payload_0_9675;
  reg        [7:0]    _zz_dataOut_payload_0_9676;
  reg        [7:0]    _zz_dataOut_payload_0_9677;
  reg        [7:0]    _zz_dataOut_payload_0_9678;
  reg        [7:0]    _zz_dataOut_payload_0_9679;
  wire                _zz_dataOut_payload_0_9680;
  wire       [7:0]    _zz_dataOut_payload_0_9681;
  wire       [7:0]    _zz_dataOut_payload_0_9682;
  wire                _zz_dataOut_payload_0_9683;
  wire       [7:0]    _zz_dataOut_payload_0_9684;
  wire       [7:0]    _zz_dataOut_payload_0_9685;
  wire                _zz_dataOut_payload_0_9686;
  wire                _zz_dataOut_payload_0_9687;
  reg        [7:0]    _zz_dataOut_payload_0_9688;
  reg        [7:0]    _zz_dataOut_payload_0_9689;
  reg        [7:0]    _zz_dataOut_payload_0_9690;
  reg        [7:0]    _zz_dataOut_payload_0_9691;
  reg        [7:0]    _zz_dataOut_payload_0_9692;
  reg        [7:0]    _zz_dataOut_payload_0_9693;
  reg        [7:0]    _zz_dataOut_payload_0_9694;
  reg        [7:0]    _zz_dataOut_payload_0_9695;
  reg        [7:0]    _zz_dataOut_payload_0_9696;
  reg        [7:0]    _zz_dataOut_payload_0_9697;
  reg        [7:0]    _zz_dataOut_payload_0_9698;
  reg        [7:0]    _zz_dataOut_payload_0_9699;
  wire                _zz_dataOut_payload_0_9700;
  wire       [7:0]    _zz_dataOut_payload_0_9701;
  wire       [7:0]    _zz_dataOut_payload_0_9702;
  wire                _zz_dataOut_payload_0_9703;
  wire       [7:0]    _zz_dataOut_payload_0_9704;
  wire       [7:0]    _zz_dataOut_payload_0_9705;
  wire                _zz_dataOut_payload_0_9706;
  wire       [7:0]    _zz_dataOut_payload_0_9707;
  wire       [7:0]    _zz_dataOut_payload_0_9708;
  wire                _zz_dataOut_payload_0_9709;
  wire       [7:0]    _zz_dataOut_payload_0_9710;
  wire       [7:0]    _zz_dataOut_payload_0_9711;
  wire                _zz_dataOut_payload_0_9712;
  wire       [7:0]    _zz_dataOut_payload_0_9713;
  wire       [7:0]    _zz_dataOut_payload_0_9714;
  wire                _zz_dataOut_payload_0_9715;
  wire       [7:0]    _zz_dataOut_payload_0_9716;
  wire       [7:0]    _zz_dataOut_payload_0_9717;
  wire                _zz_dataOut_payload_0_9718;
  wire                _zz_dataOut_payload_0_9719;
  reg        [7:0]    _zz_dataOut_payload_0_9720;
  reg        [7:0]    _zz_dataOut_payload_0_9721;
  reg        [7:0]    _zz_dataOut_payload_0_9722;
  reg        [7:0]    _zz_dataOut_payload_0_9723;
  wire                _zz_dataOut_payload_0_9724;
  wire       [7:0]    _zz_dataOut_payload_0_9725;
  wire       [7:0]    _zz_dataOut_payload_0_9726;
  wire                _zz_dataOut_payload_0_9727;
  wire       [7:0]    _zz_dataOut_payload_0_9728;
  wire       [7:0]    _zz_dataOut_payload_0_9729;
  wire                _zz_dataOut_payload_0_9730;
  wire                _zz_dataOut_payload_0_9731;
  reg        [7:0]    _zz_dataOut_payload_0_9732;
  reg        [7:0]    _zz_dataOut_payload_0_9733;
  reg        [7:0]    _zz_dataOut_payload_0_9734;
  reg        [7:0]    _zz_dataOut_payload_0_9735;
  reg        [7:0]    _zz_dataOut_payload_0_9736;
  reg        [7:0]    _zz_dataOut_payload_0_9737;
  reg        [7:0]    _zz_dataOut_payload_0_9738;
  reg        [7:0]    _zz_dataOut_payload_0_9739;
  reg        [7:0]    _zz_dataOut_payload_0_9740;
  reg        [7:0]    _zz_dataOut_payload_0_9741;
  reg        [7:0]    _zz_dataOut_payload_0_9742;
  reg        [7:0]    _zz_dataOut_payload_0_9743;
  reg        [7:0]    _zz_dataOut_payload_0_9744;
  reg        [7:0]    _zz_dataOut_payload_0_9745;
  reg        [7:0]    _zz_dataOut_payload_0_9746;
  reg        [7:0]    _zz_dataOut_payload_0_9747;
  reg        [7:0]    _zz_dataOut_payload_0_9748;
  reg        [7:0]    _zz_dataOut_payload_0_9749;
  reg        [7:0]    _zz_dataOut_payload_0_9750;
  reg        [7:0]    _zz_dataOut_payload_0_9751;
  reg        [7:0]    _zz_dataOut_payload_0_9752;
  reg        [7:0]    _zz_dataOut_payload_0_9753;
  reg        [7:0]    _zz_dataOut_payload_0_9754;
  reg        [7:0]    _zz_dataOut_payload_0_9755;
  reg        [7:0]    _zz_dataOut_payload_0_9756;
  reg        [7:0]    _zz_dataOut_payload_0_9757;
  reg        [7:0]    _zz_dataOut_payload_0_9758;
  reg        [7:0]    _zz_dataOut_payload_0_9759;
  wire                _zz_dataOut_payload_0_9760;
  wire       [7:0]    _zz_dataOut_payload_0_9761;
  wire       [7:0]    _zz_dataOut_payload_0_9762;
  wire                _zz_dataOut_payload_0_9763;
  wire       [7:0]    _zz_dataOut_payload_0_9764;
  wire       [7:0]    _zz_dataOut_payload_0_9765;
  wire                _zz_dataOut_payload_0_9766;
  wire       [7:0]    _zz_dataOut_payload_0_9767;
  wire       [7:0]    _zz_dataOut_payload_0_9768;
  wire                _zz_dataOut_payload_0_9769;
  wire       [7:0]    _zz_dataOut_payload_0_9770;
  wire       [7:0]    _zz_dataOut_payload_0_9771;
  wire                _zz_dataOut_payload_0_9772;
  wire       [7:0]    _zz_dataOut_payload_0_9773;
  wire       [7:0]    _zz_dataOut_payload_0_9774;
  wire                _zz_dataOut_payload_0_9775;
  wire       [7:0]    _zz_dataOut_payload_0_9776;
  wire       [7:0]    _zz_dataOut_payload_0_9777;
  wire                _zz_dataOut_payload_0_9778;
  wire       [7:0]    _zz_dataOut_payload_0_9779;
  wire       [7:0]    _zz_dataOut_payload_0_9780;
  wire                _zz_dataOut_payload_0_9781;
  wire       [7:0]    _zz_dataOut_payload_0_9782;
  wire       [7:0]    _zz_dataOut_payload_0_9783;
  wire                _zz_dataOut_payload_0_9784;
  wire       [7:0]    _zz_dataOut_payload_0_9785;
  wire       [7:0]    _zz_dataOut_payload_0_9786;
  wire                _zz_dataOut_payload_0_9787;
  wire       [7:0]    _zz_dataOut_payload_0_9788;
  wire       [7:0]    _zz_dataOut_payload_0_9789;
  wire                _zz_dataOut_payload_0_9790;
  wire       [7:0]    _zz_dataOut_payload_0_9791;
  wire       [7:0]    _zz_dataOut_payload_0_9792;
  wire                _zz_dataOut_payload_0_9793;
  wire       [7:0]    _zz_dataOut_payload_0_9794;
  wire       [7:0]    _zz_dataOut_payload_0_9795;
  wire                _zz_dataOut_payload_0_9796;
  wire       [7:0]    _zz_dataOut_payload_0_9797;
  wire       [7:0]    _zz_dataOut_payload_0_9798;
  wire                _zz_dataOut_payload_0_9799;
  wire       [7:0]    _zz_dataOut_payload_0_9800;
  wire       [7:0]    _zz_dataOut_payload_0_9801;
  wire                _zz_dataOut_payload_0_9802;
  wire                _zz_dataOut_payload_0_9803;
  reg        [7:0]    _zz_dataOut_payload_0_9804;
  reg        [7:0]    _zz_dataOut_payload_0_9805;
  reg        [7:0]    _zz_dataOut_payload_0_9806;
  reg        [7:0]    _zz_dataOut_payload_0_9807;
  wire                _zz_dataOut_payload_0_9808;
  wire       [7:0]    _zz_dataOut_payload_0_9809;
  wire       [7:0]    _zz_dataOut_payload_0_9810;
  wire                _zz_dataOut_payload_0_9811;
  wire       [7:0]    _zz_dataOut_payload_0_9812;
  wire       [7:0]    _zz_dataOut_payload_0_9813;
  wire                _zz_dataOut_payload_0_9814;
  wire                _zz_dataOut_payload_0_9815;
  reg        [7:0]    _zz_dataOut_payload_0_9816;
  reg        [7:0]    _zz_dataOut_payload_0_9817;
  reg        [7:0]    _zz_dataOut_payload_0_9818;
  reg        [7:0]    _zz_dataOut_payload_0_9819;
  reg        [7:0]    _zz_dataOut_payload_0_9820;
  reg        [7:0]    _zz_dataOut_payload_0_9821;
  reg        [7:0]    _zz_dataOut_payload_0_9822;
  reg        [7:0]    _zz_dataOut_payload_0_9823;
  reg        [7:0]    _zz_dataOut_payload_0_9824;
  reg        [7:0]    _zz_dataOut_payload_0_9825;
  reg        [7:0]    _zz_dataOut_payload_0_9826;
  reg        [7:0]    _zz_dataOut_payload_0_9827;
  wire                _zz_dataOut_payload_0_9828;
  wire       [7:0]    _zz_dataOut_payload_0_9829;
  wire       [7:0]    _zz_dataOut_payload_0_9830;
  wire                _zz_dataOut_payload_0_9831;
  wire       [7:0]    _zz_dataOut_payload_0_9832;
  wire       [7:0]    _zz_dataOut_payload_0_9833;
  wire                _zz_dataOut_payload_0_9834;
  wire       [7:0]    _zz_dataOut_payload_0_9835;
  wire       [7:0]    _zz_dataOut_payload_0_9836;
  wire                _zz_dataOut_payload_0_9837;
  wire       [7:0]    _zz_dataOut_payload_0_9838;
  wire       [7:0]    _zz_dataOut_payload_0_9839;
  wire                _zz_dataOut_payload_0_9840;
  wire       [7:0]    _zz_dataOut_payload_0_9841;
  wire       [7:0]    _zz_dataOut_payload_0_9842;
  wire                _zz_dataOut_payload_0_9843;
  wire       [7:0]    _zz_dataOut_payload_0_9844;
  wire       [7:0]    _zz_dataOut_payload_0_9845;
  wire                _zz_dataOut_payload_0_9846;
  wire                _zz_dataOut_payload_0_9847;
  reg        [7:0]    _zz_dataOut_payload_0_9848;
  reg        [7:0]    _zz_dataOut_payload_0_9849;
  reg        [7:0]    _zz_dataOut_payload_0_9850;
  reg        [7:0]    _zz_dataOut_payload_0_9851;
  wire                _zz_dataOut_payload_0_9852;
  wire       [7:0]    _zz_dataOut_payload_0_9853;
  wire       [7:0]    _zz_dataOut_payload_0_9854;
  wire                _zz_dataOut_payload_0_9855;
  wire       [7:0]    _zz_dataOut_payload_0_9856;
  wire       [7:0]    _zz_dataOut_payload_0_9857;
  wire                _zz_dataOut_payload_0_9858;
  wire                _zz_dataOut_payload_0_9859;
  reg        [7:0]    _zz_dataOut_payload_0_9860;
  reg        [7:0]    _zz_dataOut_payload_0_9861;
  reg        [7:0]    _zz_dataOut_payload_0_9862;
  reg        [7:0]    _zz_dataOut_payload_0_9863;
  reg        [7:0]    _zz_dataOut_payload_0_9864;
  reg        [7:0]    _zz_dataOut_payload_0_9865;
  reg        [7:0]    _zz_dataOut_payload_0_9866;
  reg        [7:0]    _zz_dataOut_payload_0_9867;
  reg        [7:0]    _zz_dataOut_payload_0_9868;
  reg        [7:0]    _zz_dataOut_payload_0_9869;
  reg        [7:0]    _zz_dataOut_payload_0_9870;
  reg        [7:0]    _zz_dataOut_payload_0_9871;
  reg        [7:0]    _zz_dataOut_payload_0_9872;
  reg        [7:0]    _zz_dataOut_payload_0_9873;
  reg        [7:0]    _zz_dataOut_payload_0_9874;
  reg        [7:0]    _zz_dataOut_payload_0_9875;
  reg        [7:0]    _zz_dataOut_payload_0_9876;
  reg        [7:0]    _zz_dataOut_payload_0_9877;
  reg        [7:0]    _zz_dataOut_payload_0_9878;
  reg        [7:0]    _zz_dataOut_payload_0_9879;
  reg        [7:0]    _zz_dataOut_payload_0_9880;
  reg        [7:0]    _zz_dataOut_payload_0_9881;
  reg        [7:0]    _zz_dataOut_payload_0_9882;
  reg        [7:0]    _zz_dataOut_payload_0_9883;
  reg        [7:0]    _zz_dataOut_payload_0_9884;
  reg        [7:0]    _zz_dataOut_payload_0_9885;
  reg        [7:0]    _zz_dataOut_payload_0_9886;
  reg        [7:0]    _zz_dataOut_payload_0_9887;
  reg        [7:0]    _zz_dataOut_payload_0_9888;
  reg        [7:0]    _zz_dataOut_payload_0_9889;
  reg        [7:0]    _zz_dataOut_payload_0_9890;
  reg        [7:0]    _zz_dataOut_payload_0_9891;
  reg        [7:0]    _zz_dataOut_payload_0_9892;
  reg        [7:0]    _zz_dataOut_payload_0_9893;
  reg        [7:0]    _zz_dataOut_payload_0_9894;
  reg        [7:0]    _zz_dataOut_payload_0_9895;
  reg        [7:0]    _zz_dataOut_payload_0_9896;
  reg        [7:0]    _zz_dataOut_payload_0_9897;
  reg        [7:0]    _zz_dataOut_payload_0_9898;
  reg        [7:0]    _zz_dataOut_payload_0_9899;
  reg        [7:0]    _zz_dataOut_payload_0_9900;
  reg        [7:0]    _zz_dataOut_payload_0_9901;
  reg        [7:0]    _zz_dataOut_payload_0_9902;
  reg        [7:0]    _zz_dataOut_payload_0_9903;
  reg        [7:0]    _zz_dataOut_payload_0_9904;
  reg        [7:0]    _zz_dataOut_payload_0_9905;
  reg        [7:0]    _zz_dataOut_payload_0_9906;
  reg        [7:0]    _zz_dataOut_payload_0_9907;
  reg        [7:0]    _zz_dataOut_payload_0_9908;
  reg        [7:0]    _zz_dataOut_payload_0_9909;
  reg        [7:0]    _zz_dataOut_payload_0_9910;
  reg        [7:0]    _zz_dataOut_payload_0_9911;
  reg        [7:0]    _zz_dataOut_payload_0_9912;
  reg        [7:0]    _zz_dataOut_payload_0_9913;
  reg        [7:0]    _zz_dataOut_payload_0_9914;
  reg        [7:0]    _zz_dataOut_payload_0_9915;
  reg        [7:0]    _zz_dataOut_payload_0_9916;
  reg        [7:0]    _zz_dataOut_payload_0_9917;
  reg        [7:0]    _zz_dataOut_payload_0_9918;
  reg        [7:0]    _zz_dataOut_payload_0_9919;
  reg        [7:0]    _zz_dataOut_payload_0_9920;
  reg        [7:0]    _zz_dataOut_payload_0_9921;
  reg        [7:0]    _zz_dataOut_payload_0_9922;
  reg        [7:0]    _zz_dataOut_payload_0_9923;
  reg        [7:0]    _zz_dataOut_payload_0_9924;
  reg        [7:0]    _zz_dataOut_payload_0_9925;
  reg        [7:0]    _zz_dataOut_payload_0_9926;
  reg        [7:0]    _zz_dataOut_payload_0_9927;
  reg        [7:0]    _zz_dataOut_payload_0_9928;
  reg        [7:0]    _zz_dataOut_payload_0_9929;
  reg        [7:0]    _zz_dataOut_payload_0_9930;
  reg        [7:0]    _zz_dataOut_payload_0_9931;
  reg        [7:0]    _zz_dataOut_payload_0_9932;
  reg        [7:0]    _zz_dataOut_payload_0_9933;
  reg        [7:0]    _zz_dataOut_payload_0_9934;
  reg        [7:0]    _zz_dataOut_payload_0_9935;
  reg        [7:0]    _zz_dataOut_payload_0_9936;
  reg        [7:0]    _zz_dataOut_payload_0_9937;
  reg        [7:0]    _zz_dataOut_payload_0_9938;
  reg        [7:0]    _zz_dataOut_payload_0_9939;
  reg        [7:0]    _zz_dataOut_payload_0_9940;
  reg        [7:0]    _zz_dataOut_payload_0_9941;
  reg        [7:0]    _zz_dataOut_payload_0_9942;
  reg        [7:0]    _zz_dataOut_payload_0_9943;
  reg        [7:0]    _zz_dataOut_payload_0_9944;
  reg        [7:0]    _zz_dataOut_payload_0_9945;
  reg        [7:0]    _zz_dataOut_payload_0_9946;
  reg        [7:0]    _zz_dataOut_payload_0_9947;
  reg        [7:0]    _zz_dataOut_payload_0_9948;
  reg        [7:0]    _zz_dataOut_payload_0_9949;
  reg        [7:0]    _zz_dataOut_payload_0_9950;
  reg        [7:0]    _zz_dataOut_payload_0_9951;
  reg        [7:0]    _zz_dataOut_payload_0_9952;
  reg        [7:0]    _zz_dataOut_payload_0_9953;
  reg        [7:0]    _zz_dataOut_payload_0_9954;
  reg        [7:0]    _zz_dataOut_payload_0_9955;
  reg        [7:0]    _zz_dataOut_payload_0_9956;
  reg        [7:0]    _zz_dataOut_payload_0_9957;
  reg        [7:0]    _zz_dataOut_payload_0_9958;
  reg        [7:0]    _zz_dataOut_payload_0_9959;
  reg        [7:0]    _zz_dataOut_payload_0_9960;
  reg        [7:0]    _zz_dataOut_payload_0_9961;
  reg        [7:0]    _zz_dataOut_payload_0_9962;
  reg        [7:0]    _zz_dataOut_payload_0_9963;
  reg        [7:0]    _zz_dataOut_payload_0_9964;
  reg        [7:0]    _zz_dataOut_payload_0_9965;
  reg        [7:0]    _zz_dataOut_payload_0_9966;
  reg        [7:0]    _zz_dataOut_payload_0_9967;
  reg        [7:0]    _zz_dataOut_payload_0_9968;
  reg        [7:0]    _zz_dataOut_payload_0_9969;
  reg        [7:0]    _zz_dataOut_payload_0_9970;
  reg        [7:0]    _zz_dataOut_payload_0_9971;
  reg        [7:0]    _zz_dataOut_payload_0_9972;
  reg        [7:0]    _zz_dataOut_payload_0_9973;
  reg        [7:0]    _zz_dataOut_payload_0_9974;
  reg        [7:0]    _zz_dataOut_payload_0_9975;
  reg        [7:0]    _zz_dataOut_payload_0_9976;
  reg        [7:0]    _zz_dataOut_payload_0_9977;
  reg        [7:0]    _zz_dataOut_payload_0_9978;
  reg        [7:0]    _zz_dataOut_payload_0_9979;
  reg        [7:0]    _zz_dataOut_payload_0_9980;
  reg        [7:0]    _zz_dataOut_payload_0_9981;
  reg        [7:0]    _zz_dataOut_payload_0_9982;
  reg        [7:0]    _zz_dataOut_payload_0_9983;
  wire                _zz_dataOut_payload_0_9984;
  wire       [7:0]    _zz_dataOut_payload_0_9985;
  wire       [7:0]    _zz_dataOut_payload_0_9986;
  wire                _zz_dataOut_payload_0_9987;
  wire       [7:0]    _zz_dataOut_payload_0_9988;
  wire       [7:0]    _zz_dataOut_payload_0_9989;
  wire                _zz_dataOut_payload_0_9990;
  wire       [7:0]    _zz_dataOut_payload_0_9991;
  wire       [7:0]    _zz_dataOut_payload_0_9992;
  wire                _zz_dataOut_payload_0_9993;
  wire       [7:0]    _zz_dataOut_payload_0_9994;
  wire       [7:0]    _zz_dataOut_payload_0_9995;
  wire                _zz_dataOut_payload_0_9996;
  wire       [7:0]    _zz_dataOut_payload_0_9997;
  wire       [7:0]    _zz_dataOut_payload_0_9998;
  wire                _zz_dataOut_payload_0_9999;
  wire       [7:0]    _zz_dataOut_payload_0_10000;
  wire       [7:0]    _zz_dataOut_payload_0_10001;
  wire                _zz_dataOut_payload_0_10002;
  wire       [7:0]    _zz_dataOut_payload_0_10003;
  wire       [7:0]    _zz_dataOut_payload_0_10004;
  wire                _zz_dataOut_payload_0_10005;
  wire       [7:0]    _zz_dataOut_payload_0_10006;
  wire       [7:0]    _zz_dataOut_payload_0_10007;
  wire                _zz_dataOut_payload_0_10008;
  wire       [7:0]    _zz_dataOut_payload_0_10009;
  wire       [7:0]    _zz_dataOut_payload_0_10010;
  wire                _zz_dataOut_payload_0_10011;
  wire       [7:0]    _zz_dataOut_payload_0_10012;
  wire       [7:0]    _zz_dataOut_payload_0_10013;
  wire                _zz_dataOut_payload_0_10014;
  wire       [7:0]    _zz_dataOut_payload_0_10015;
  wire       [7:0]    _zz_dataOut_payload_0_10016;
  wire                _zz_dataOut_payload_0_10017;
  wire       [7:0]    _zz_dataOut_payload_0_10018;
  wire       [7:0]    _zz_dataOut_payload_0_10019;
  wire                _zz_dataOut_payload_0_10020;
  wire       [7:0]    _zz_dataOut_payload_0_10021;
  wire       [7:0]    _zz_dataOut_payload_0_10022;
  wire                _zz_dataOut_payload_0_10023;
  wire       [7:0]    _zz_dataOut_payload_0_10024;
  wire       [7:0]    _zz_dataOut_payload_0_10025;
  wire                _zz_dataOut_payload_0_10026;
  wire       [7:0]    _zz_dataOut_payload_0_10027;
  wire       [7:0]    _zz_dataOut_payload_0_10028;
  wire                _zz_dataOut_payload_0_10029;
  wire       [7:0]    _zz_dataOut_payload_0_10030;
  wire       [7:0]    _zz_dataOut_payload_0_10031;
  wire                _zz_dataOut_payload_0_10032;
  wire       [7:0]    _zz_dataOut_payload_0_10033;
  wire       [7:0]    _zz_dataOut_payload_0_10034;
  wire                _zz_dataOut_payload_0_10035;
  wire       [7:0]    _zz_dataOut_payload_0_10036;
  wire       [7:0]    _zz_dataOut_payload_0_10037;
  wire                _zz_dataOut_payload_0_10038;
  wire       [7:0]    _zz_dataOut_payload_0_10039;
  wire       [7:0]    _zz_dataOut_payload_0_10040;
  wire                _zz_dataOut_payload_0_10041;
  wire       [7:0]    _zz_dataOut_payload_0_10042;
  wire       [7:0]    _zz_dataOut_payload_0_10043;
  wire                _zz_dataOut_payload_0_10044;
  wire       [7:0]    _zz_dataOut_payload_0_10045;
  wire       [7:0]    _zz_dataOut_payload_0_10046;
  wire                _zz_dataOut_payload_0_10047;
  wire       [7:0]    _zz_dataOut_payload_0_10048;
  wire       [7:0]    _zz_dataOut_payload_0_10049;
  wire                _zz_dataOut_payload_0_10050;
  wire       [7:0]    _zz_dataOut_payload_0_10051;
  wire       [7:0]    _zz_dataOut_payload_0_10052;
  wire                _zz_dataOut_payload_0_10053;
  wire       [7:0]    _zz_dataOut_payload_0_10054;
  wire       [7:0]    _zz_dataOut_payload_0_10055;
  wire                _zz_dataOut_payload_0_10056;
  wire       [7:0]    _zz_dataOut_payload_0_10057;
  wire       [7:0]    _zz_dataOut_payload_0_10058;
  wire                _zz_dataOut_payload_0_10059;
  wire       [7:0]    _zz_dataOut_payload_0_10060;
  wire       [7:0]    _zz_dataOut_payload_0_10061;
  wire                _zz_dataOut_payload_0_10062;
  wire       [7:0]    _zz_dataOut_payload_0_10063;
  wire       [7:0]    _zz_dataOut_payload_0_10064;
  wire                _zz_dataOut_payload_0_10065;
  wire       [7:0]    _zz_dataOut_payload_0_10066;
  wire       [7:0]    _zz_dataOut_payload_0_10067;
  wire                _zz_dataOut_payload_0_10068;
  wire       [7:0]    _zz_dataOut_payload_0_10069;
  wire       [7:0]    _zz_dataOut_payload_0_10070;
  wire                _zz_dataOut_payload_0_10071;
  wire       [7:0]    _zz_dataOut_payload_0_10072;
  wire       [7:0]    _zz_dataOut_payload_0_10073;
  wire                _zz_dataOut_payload_0_10074;
  wire       [7:0]    _zz_dataOut_payload_0_10075;
  wire       [7:0]    _zz_dataOut_payload_0_10076;
  wire                _zz_dataOut_payload_0_10077;
  wire       [7:0]    _zz_dataOut_payload_0_10078;
  wire       [7:0]    _zz_dataOut_payload_0_10079;
  wire                _zz_dataOut_payload_0_10080;
  wire       [7:0]    _zz_dataOut_payload_0_10081;
  wire       [7:0]    _zz_dataOut_payload_0_10082;
  wire                _zz_dataOut_payload_0_10083;
  wire       [7:0]    _zz_dataOut_payload_0_10084;
  wire       [7:0]    _zz_dataOut_payload_0_10085;
  wire                _zz_dataOut_payload_0_10086;
  wire       [7:0]    _zz_dataOut_payload_0_10087;
  wire       [7:0]    _zz_dataOut_payload_0_10088;
  wire                _zz_dataOut_payload_0_10089;
  wire       [7:0]    _zz_dataOut_payload_0_10090;
  wire       [7:0]    _zz_dataOut_payload_0_10091;
  wire                _zz_dataOut_payload_0_10092;
  wire       [7:0]    _zz_dataOut_payload_0_10093;
  wire       [7:0]    _zz_dataOut_payload_0_10094;
  wire                _zz_dataOut_payload_0_10095;
  wire       [7:0]    _zz_dataOut_payload_0_10096;
  wire       [7:0]    _zz_dataOut_payload_0_10097;
  wire                _zz_dataOut_payload_0_10098;
  wire       [7:0]    _zz_dataOut_payload_0_10099;
  wire       [7:0]    _zz_dataOut_payload_0_10100;
  wire                _zz_dataOut_payload_0_10101;
  wire       [7:0]    _zz_dataOut_payload_0_10102;
  wire       [7:0]    _zz_dataOut_payload_0_10103;
  wire                _zz_dataOut_payload_0_10104;
  wire       [7:0]    _zz_dataOut_payload_0_10105;
  wire       [7:0]    _zz_dataOut_payload_0_10106;
  wire                _zz_dataOut_payload_0_10107;
  wire       [7:0]    _zz_dataOut_payload_0_10108;
  wire       [7:0]    _zz_dataOut_payload_0_10109;
  wire                _zz_dataOut_payload_0_10110;
  wire       [7:0]    _zz_dataOut_payload_0_10111;
  wire       [7:0]    _zz_dataOut_payload_0_10112;
  wire                _zz_dataOut_payload_0_10113;
  wire       [7:0]    _zz_dataOut_payload_0_10114;
  wire       [7:0]    _zz_dataOut_payload_0_10115;
  wire                _zz_dataOut_payload_0_10116;
  wire       [7:0]    _zz_dataOut_payload_0_10117;
  wire       [7:0]    _zz_dataOut_payload_0_10118;
  wire                _zz_dataOut_payload_0_10119;
  wire       [7:0]    _zz_dataOut_payload_0_10120;
  wire       [7:0]    _zz_dataOut_payload_0_10121;
  wire                _zz_dataOut_payload_0_10122;
  wire       [7:0]    _zz_dataOut_payload_0_10123;
  wire       [7:0]    _zz_dataOut_payload_0_10124;
  wire                _zz_dataOut_payload_0_10125;
  wire       [7:0]    _zz_dataOut_payload_0_10126;
  wire       [7:0]    _zz_dataOut_payload_0_10127;
  wire                _zz_dataOut_payload_0_10128;
  wire       [7:0]    _zz_dataOut_payload_0_10129;
  wire       [7:0]    _zz_dataOut_payload_0_10130;
  wire                _zz_dataOut_payload_0_10131;
  wire       [7:0]    _zz_dataOut_payload_0_10132;
  wire       [7:0]    _zz_dataOut_payload_0_10133;
  wire                _zz_dataOut_payload_0_10134;
  wire       [7:0]    _zz_dataOut_payload_0_10135;
  wire       [7:0]    _zz_dataOut_payload_0_10136;
  wire                _zz_dataOut_payload_0_10137;
  wire       [7:0]    _zz_dataOut_payload_0_10138;
  wire       [7:0]    _zz_dataOut_payload_0_10139;
  wire                _zz_dataOut_payload_0_10140;
  wire       [7:0]    _zz_dataOut_payload_0_10141;
  wire       [7:0]    _zz_dataOut_payload_0_10142;
  wire                _zz_dataOut_payload_0_10143;
  wire       [7:0]    _zz_dataOut_payload_0_10144;
  wire       [7:0]    _zz_dataOut_payload_0_10145;
  wire                _zz_dataOut_payload_0_10146;
  wire       [7:0]    _zz_dataOut_payload_0_10147;
  wire       [7:0]    _zz_dataOut_payload_0_10148;
  wire                _zz_dataOut_payload_0_10149;
  wire       [7:0]    _zz_dataOut_payload_0_10150;
  wire       [7:0]    _zz_dataOut_payload_0_10151;
  wire                _zz_dataOut_payload_0_10152;
  wire       [7:0]    _zz_dataOut_payload_0_10153;
  wire       [7:0]    _zz_dataOut_payload_0_10154;
  wire                _zz_dataOut_payload_0_10155;
  wire       [7:0]    _zz_dataOut_payload_0_10156;
  wire       [7:0]    _zz_dataOut_payload_0_10157;
  wire                _zz_dataOut_payload_0_10158;
  wire       [7:0]    _zz_dataOut_payload_0_10159;
  wire       [7:0]    _zz_dataOut_payload_0_10160;
  wire                _zz_dataOut_payload_0_10161;
  wire       [7:0]    _zz_dataOut_payload_0_10162;
  wire       [7:0]    _zz_dataOut_payload_0_10163;
  wire                _zz_dataOut_payload_0_10164;
  wire       [7:0]    _zz_dataOut_payload_0_10165;
  wire       [7:0]    _zz_dataOut_payload_0_10166;
  wire                _zz_dataOut_payload_0_10167;
  wire       [7:0]    _zz_dataOut_payload_0_10168;
  wire       [7:0]    _zz_dataOut_payload_0_10169;
  wire                _zz_dataOut_payload_0_10170;
  wire                _zz_dataOut_payload_0_10171;
  reg        [7:0]    _zz_dataOut_payload_0_10172;
  reg        [7:0]    _zz_dataOut_payload_0_10173;
  reg        [7:0]    _zz_dataOut_payload_0_10174;
  reg        [7:0]    _zz_dataOut_payload_0_10175;
  wire                _zz_dataOut_payload_0_10176;
  wire       [7:0]    _zz_dataOut_payload_0_10177;
  wire       [7:0]    _zz_dataOut_payload_0_10178;
  wire                _zz_dataOut_payload_0_10179;
  wire       [7:0]    _zz_dataOut_payload_0_10180;
  wire       [7:0]    _zz_dataOut_payload_0_10181;
  wire                _zz_dataOut_payload_0_10182;
  wire                _zz_dataOut_payload_0_10183;
  reg        [7:0]    _zz_dataOut_payload_0_10184;
  reg        [7:0]    _zz_dataOut_payload_0_10185;
  reg        [7:0]    _zz_dataOut_payload_0_10186;
  reg        [7:0]    _zz_dataOut_payload_0_10187;
  reg        [7:0]    _zz_dataOut_payload_0_10188;
  reg        [7:0]    _zz_dataOut_payload_0_10189;
  reg        [7:0]    _zz_dataOut_payload_0_10190;
  reg        [7:0]    _zz_dataOut_payload_0_10191;
  reg        [7:0]    _zz_dataOut_payload_0_10192;
  reg        [7:0]    _zz_dataOut_payload_0_10193;
  reg        [7:0]    _zz_dataOut_payload_0_10194;
  reg        [7:0]    _zz_dataOut_payload_0_10195;
  wire                _zz_dataOut_payload_0_10196;
  wire       [7:0]    _zz_dataOut_payload_0_10197;
  wire       [7:0]    _zz_dataOut_payload_0_10198;
  wire                _zz_dataOut_payload_0_10199;
  wire       [7:0]    _zz_dataOut_payload_0_10200;
  wire       [7:0]    _zz_dataOut_payload_0_10201;
  wire                _zz_dataOut_payload_0_10202;
  wire       [7:0]    _zz_dataOut_payload_0_10203;
  wire       [7:0]    _zz_dataOut_payload_0_10204;
  wire                _zz_dataOut_payload_0_10205;
  wire       [7:0]    _zz_dataOut_payload_0_10206;
  wire       [7:0]    _zz_dataOut_payload_0_10207;
  wire                _zz_dataOut_payload_0_10208;
  wire       [7:0]    _zz_dataOut_payload_0_10209;
  wire       [7:0]    _zz_dataOut_payload_0_10210;
  wire                _zz_dataOut_payload_0_10211;
  wire       [7:0]    _zz_dataOut_payload_0_10212;
  wire       [7:0]    _zz_dataOut_payload_0_10213;
  wire                _zz_dataOut_payload_0_10214;
  wire                _zz_dataOut_payload_0_10215;
  reg        [7:0]    _zz_dataOut_payload_0_10216;
  reg        [7:0]    _zz_dataOut_payload_0_10217;
  reg        [7:0]    _zz_dataOut_payload_0_10218;
  reg        [7:0]    _zz_dataOut_payload_0_10219;
  wire                _zz_dataOut_payload_0_10220;
  wire       [7:0]    _zz_dataOut_payload_0_10221;
  wire       [7:0]    _zz_dataOut_payload_0_10222;
  wire                _zz_dataOut_payload_0_10223;
  wire       [7:0]    _zz_dataOut_payload_0_10224;
  wire       [7:0]    _zz_dataOut_payload_0_10225;
  wire                _zz_dataOut_payload_0_10226;
  wire                _zz_dataOut_payload_0_10227;
  reg        [7:0]    _zz_dataOut_payload_0_10228;
  reg        [7:0]    _zz_dataOut_payload_0_10229;
  reg        [7:0]    _zz_dataOut_payload_0_10230;
  reg        [7:0]    _zz_dataOut_payload_0_10231;
  reg        [7:0]    _zz_dataOut_payload_0_10232;
  reg        [7:0]    _zz_dataOut_payload_0_10233;
  reg        [7:0]    _zz_dataOut_payload_0_10234;
  reg        [7:0]    _zz_dataOut_payload_0_10235;
  reg        [7:0]    _zz_dataOut_payload_0_10236;
  reg        [7:0]    _zz_dataOut_payload_0_10237;
  reg        [7:0]    _zz_dataOut_payload_0_10238;
  reg        [7:0]    _zz_dataOut_payload_0_10239;
  reg        [7:0]    _zz_dataOut_payload_0_10240;
  reg        [7:0]    _zz_dataOut_payload_0_10241;
  reg        [7:0]    _zz_dataOut_payload_0_10242;
  reg        [7:0]    _zz_dataOut_payload_0_10243;
  reg        [7:0]    _zz_dataOut_payload_0_10244;
  reg        [7:0]    _zz_dataOut_payload_0_10245;
  reg        [7:0]    _zz_dataOut_payload_0_10246;
  reg        [7:0]    _zz_dataOut_payload_0_10247;
  reg        [7:0]    _zz_dataOut_payload_0_10248;
  reg        [7:0]    _zz_dataOut_payload_0_10249;
  reg        [7:0]    _zz_dataOut_payload_0_10250;
  reg        [7:0]    _zz_dataOut_payload_0_10251;
  reg        [7:0]    _zz_dataOut_payload_0_10252;
  reg        [7:0]    _zz_dataOut_payload_0_10253;
  reg        [7:0]    _zz_dataOut_payload_0_10254;
  reg        [7:0]    _zz_dataOut_payload_0_10255;
  wire                _zz_dataOut_payload_0_10256;
  wire       [7:0]    _zz_dataOut_payload_0_10257;
  wire       [7:0]    _zz_dataOut_payload_0_10258;
  wire                _zz_dataOut_payload_0_10259;
  wire       [7:0]    _zz_dataOut_payload_0_10260;
  wire       [7:0]    _zz_dataOut_payload_0_10261;
  wire                _zz_dataOut_payload_0_10262;
  wire       [7:0]    _zz_dataOut_payload_0_10263;
  wire       [7:0]    _zz_dataOut_payload_0_10264;
  wire                _zz_dataOut_payload_0_10265;
  wire       [7:0]    _zz_dataOut_payload_0_10266;
  wire       [7:0]    _zz_dataOut_payload_0_10267;
  wire                _zz_dataOut_payload_0_10268;
  wire       [7:0]    _zz_dataOut_payload_0_10269;
  wire       [7:0]    _zz_dataOut_payload_0_10270;
  wire                _zz_dataOut_payload_0_10271;
  wire       [7:0]    _zz_dataOut_payload_0_10272;
  wire       [7:0]    _zz_dataOut_payload_0_10273;
  wire                _zz_dataOut_payload_0_10274;
  wire       [7:0]    _zz_dataOut_payload_0_10275;
  wire       [7:0]    _zz_dataOut_payload_0_10276;
  wire                _zz_dataOut_payload_0_10277;
  wire       [7:0]    _zz_dataOut_payload_0_10278;
  wire       [7:0]    _zz_dataOut_payload_0_10279;
  wire                _zz_dataOut_payload_0_10280;
  wire       [7:0]    _zz_dataOut_payload_0_10281;
  wire       [7:0]    _zz_dataOut_payload_0_10282;
  wire                _zz_dataOut_payload_0_10283;
  wire       [7:0]    _zz_dataOut_payload_0_10284;
  wire       [7:0]    _zz_dataOut_payload_0_10285;
  wire                _zz_dataOut_payload_0_10286;
  wire       [7:0]    _zz_dataOut_payload_0_10287;
  wire       [7:0]    _zz_dataOut_payload_0_10288;
  wire                _zz_dataOut_payload_0_10289;
  wire       [7:0]    _zz_dataOut_payload_0_10290;
  wire       [7:0]    _zz_dataOut_payload_0_10291;
  wire                _zz_dataOut_payload_0_10292;
  wire       [7:0]    _zz_dataOut_payload_0_10293;
  wire       [7:0]    _zz_dataOut_payload_0_10294;
  wire                _zz_dataOut_payload_0_10295;
  wire       [7:0]    _zz_dataOut_payload_0_10296;
  wire       [7:0]    _zz_dataOut_payload_0_10297;
  wire                _zz_dataOut_payload_0_10298;
  wire                _zz_dataOut_payload_0_10299;
  reg        [7:0]    _zz_dataOut_payload_0_10300;
  reg        [7:0]    _zz_dataOut_payload_0_10301;
  reg        [7:0]    _zz_dataOut_payload_0_10302;
  reg        [7:0]    _zz_dataOut_payload_0_10303;
  wire                _zz_dataOut_payload_0_10304;
  wire       [7:0]    _zz_dataOut_payload_0_10305;
  wire       [7:0]    _zz_dataOut_payload_0_10306;
  wire                _zz_dataOut_payload_0_10307;
  wire       [7:0]    _zz_dataOut_payload_0_10308;
  wire       [7:0]    _zz_dataOut_payload_0_10309;
  wire                _zz_dataOut_payload_0_10310;
  wire                _zz_dataOut_payload_0_10311;
  reg        [7:0]    _zz_dataOut_payload_0_10312;
  reg        [7:0]    _zz_dataOut_payload_0_10313;
  reg        [7:0]    _zz_dataOut_payload_0_10314;
  reg        [7:0]    _zz_dataOut_payload_0_10315;
  reg        [7:0]    _zz_dataOut_payload_0_10316;
  reg        [7:0]    _zz_dataOut_payload_0_10317;
  reg        [7:0]    _zz_dataOut_payload_0_10318;
  reg        [7:0]    _zz_dataOut_payload_0_10319;
  reg        [7:0]    _zz_dataOut_payload_0_10320;
  reg        [7:0]    _zz_dataOut_payload_0_10321;
  reg        [7:0]    _zz_dataOut_payload_0_10322;
  reg        [7:0]    _zz_dataOut_payload_0_10323;
  wire                _zz_dataOut_payload_0_10324;
  wire       [7:0]    _zz_dataOut_payload_0_10325;
  wire       [7:0]    _zz_dataOut_payload_0_10326;
  wire                _zz_dataOut_payload_0_10327;
  wire       [7:0]    _zz_dataOut_payload_0_10328;
  wire       [7:0]    _zz_dataOut_payload_0_10329;
  wire                _zz_dataOut_payload_0_10330;
  wire       [7:0]    _zz_dataOut_payload_0_10331;
  wire       [7:0]    _zz_dataOut_payload_0_10332;
  wire                _zz_dataOut_payload_0_10333;
  wire       [7:0]    _zz_dataOut_payload_0_10334;
  wire       [7:0]    _zz_dataOut_payload_0_10335;
  wire                _zz_dataOut_payload_0_10336;
  wire       [7:0]    _zz_dataOut_payload_0_10337;
  wire       [7:0]    _zz_dataOut_payload_0_10338;
  wire                _zz_dataOut_payload_0_10339;
  wire       [7:0]    _zz_dataOut_payload_0_10340;
  wire       [7:0]    _zz_dataOut_payload_0_10341;
  wire                _zz_dataOut_payload_0_10342;
  wire                _zz_dataOut_payload_0_10343;
  reg        [7:0]    _zz_dataOut_payload_0_10344;
  reg        [7:0]    _zz_dataOut_payload_0_10345;
  reg        [7:0]    _zz_dataOut_payload_0_10346;
  reg        [7:0]    _zz_dataOut_payload_0_10347;
  wire                _zz_dataOut_payload_0_10348;
  wire       [7:0]    _zz_dataOut_payload_0_10349;
  wire       [7:0]    _zz_dataOut_payload_0_10350;
  wire                _zz_dataOut_payload_0_10351;
  wire       [7:0]    _zz_dataOut_payload_0_10352;
  wire       [7:0]    _zz_dataOut_payload_0_10353;
  wire                _zz_dataOut_payload_0_10354;
  wire                _zz_dataOut_payload_0_10355;
  reg        [7:0]    _zz_dataOut_payload_0_10356;
  reg        [7:0]    _zz_dataOut_payload_0_10357;
  reg        [7:0]    _zz_dataOut_payload_0_10358;
  reg        [7:0]    _zz_dataOut_payload_0_10359;
  reg        [7:0]    _zz_dataOut_payload_0_10360;
  reg        [7:0]    _zz_dataOut_payload_0_10361;
  reg        [7:0]    _zz_dataOut_payload_0_10362;
  reg        [7:0]    _zz_dataOut_payload_0_10363;
  reg        [7:0]    _zz_dataOut_payload_0_10364;
  reg        [7:0]    _zz_dataOut_payload_0_10365;
  reg        [7:0]    _zz_dataOut_payload_0_10366;
  reg        [7:0]    _zz_dataOut_payload_0_10367;
  reg        [7:0]    _zz_dataOut_payload_0_10368;
  reg        [7:0]    _zz_dataOut_payload_0_10369;
  reg        [7:0]    _zz_dataOut_payload_0_10370;
  reg        [7:0]    _zz_dataOut_payload_0_10371;
  reg        [7:0]    _zz_dataOut_payload_0_10372;
  reg        [7:0]    _zz_dataOut_payload_0_10373;
  reg        [7:0]    _zz_dataOut_payload_0_10374;
  reg        [7:0]    _zz_dataOut_payload_0_10375;
  reg        [7:0]    _zz_dataOut_payload_0_10376;
  reg        [7:0]    _zz_dataOut_payload_0_10377;
  reg        [7:0]    _zz_dataOut_payload_0_10378;
  reg        [7:0]    _zz_dataOut_payload_0_10379;
  reg        [7:0]    _zz_dataOut_payload_0_10380;
  reg        [7:0]    _zz_dataOut_payload_0_10381;
  reg        [7:0]    _zz_dataOut_payload_0_10382;
  reg        [7:0]    _zz_dataOut_payload_0_10383;
  reg        [7:0]    _zz_dataOut_payload_0_10384;
  reg        [7:0]    _zz_dataOut_payload_0_10385;
  reg        [7:0]    _zz_dataOut_payload_0_10386;
  reg        [7:0]    _zz_dataOut_payload_0_10387;
  reg        [7:0]    _zz_dataOut_payload_0_10388;
  reg        [7:0]    _zz_dataOut_payload_0_10389;
  reg        [7:0]    _zz_dataOut_payload_0_10390;
  reg        [7:0]    _zz_dataOut_payload_0_10391;
  reg        [7:0]    _zz_dataOut_payload_0_10392;
  reg        [7:0]    _zz_dataOut_payload_0_10393;
  reg        [7:0]    _zz_dataOut_payload_0_10394;
  reg        [7:0]    _zz_dataOut_payload_0_10395;
  reg        [7:0]    _zz_dataOut_payload_0_10396;
  reg        [7:0]    _zz_dataOut_payload_0_10397;
  reg        [7:0]    _zz_dataOut_payload_0_10398;
  reg        [7:0]    _zz_dataOut_payload_0_10399;
  reg        [7:0]    _zz_dataOut_payload_0_10400;
  reg        [7:0]    _zz_dataOut_payload_0_10401;
  reg        [7:0]    _zz_dataOut_payload_0_10402;
  reg        [7:0]    _zz_dataOut_payload_0_10403;
  reg        [7:0]    _zz_dataOut_payload_0_10404;
  reg        [7:0]    _zz_dataOut_payload_0_10405;
  reg        [7:0]    _zz_dataOut_payload_0_10406;
  reg        [7:0]    _zz_dataOut_payload_0_10407;
  reg        [7:0]    _zz_dataOut_payload_0_10408;
  reg        [7:0]    _zz_dataOut_payload_0_10409;
  reg        [7:0]    _zz_dataOut_payload_0_10410;
  reg        [7:0]    _zz_dataOut_payload_0_10411;
  reg        [7:0]    _zz_dataOut_payload_0_10412;
  reg        [7:0]    _zz_dataOut_payload_0_10413;
  reg        [7:0]    _zz_dataOut_payload_0_10414;
  reg        [7:0]    _zz_dataOut_payload_0_10415;
  wire                _zz_dataOut_payload_0_10416;
  wire       [7:0]    _zz_dataOut_payload_0_10417;
  wire       [7:0]    _zz_dataOut_payload_0_10418;
  wire                _zz_dataOut_payload_0_10419;
  wire       [7:0]    _zz_dataOut_payload_0_10420;
  wire       [7:0]    _zz_dataOut_payload_0_10421;
  wire                _zz_dataOut_payload_0_10422;
  wire       [7:0]    _zz_dataOut_payload_0_10423;
  wire       [7:0]    _zz_dataOut_payload_0_10424;
  wire                _zz_dataOut_payload_0_10425;
  wire       [7:0]    _zz_dataOut_payload_0_10426;
  wire       [7:0]    _zz_dataOut_payload_0_10427;
  wire                _zz_dataOut_payload_0_10428;
  wire       [7:0]    _zz_dataOut_payload_0_10429;
  wire       [7:0]    _zz_dataOut_payload_0_10430;
  wire                _zz_dataOut_payload_0_10431;
  wire       [7:0]    _zz_dataOut_payload_0_10432;
  wire       [7:0]    _zz_dataOut_payload_0_10433;
  wire                _zz_dataOut_payload_0_10434;
  wire       [7:0]    _zz_dataOut_payload_0_10435;
  wire       [7:0]    _zz_dataOut_payload_0_10436;
  wire                _zz_dataOut_payload_0_10437;
  wire       [7:0]    _zz_dataOut_payload_0_10438;
  wire       [7:0]    _zz_dataOut_payload_0_10439;
  wire                _zz_dataOut_payload_0_10440;
  wire       [7:0]    _zz_dataOut_payload_0_10441;
  wire       [7:0]    _zz_dataOut_payload_0_10442;
  wire                _zz_dataOut_payload_0_10443;
  wire       [7:0]    _zz_dataOut_payload_0_10444;
  wire       [7:0]    _zz_dataOut_payload_0_10445;
  wire                _zz_dataOut_payload_0_10446;
  wire       [7:0]    _zz_dataOut_payload_0_10447;
  wire       [7:0]    _zz_dataOut_payload_0_10448;
  wire                _zz_dataOut_payload_0_10449;
  wire       [7:0]    _zz_dataOut_payload_0_10450;
  wire       [7:0]    _zz_dataOut_payload_0_10451;
  wire                _zz_dataOut_payload_0_10452;
  wire       [7:0]    _zz_dataOut_payload_0_10453;
  wire       [7:0]    _zz_dataOut_payload_0_10454;
  wire                _zz_dataOut_payload_0_10455;
  wire       [7:0]    _zz_dataOut_payload_0_10456;
  wire       [7:0]    _zz_dataOut_payload_0_10457;
  wire                _zz_dataOut_payload_0_10458;
  wire       [7:0]    _zz_dataOut_payload_0_10459;
  wire       [7:0]    _zz_dataOut_payload_0_10460;
  wire                _zz_dataOut_payload_0_10461;
  wire       [7:0]    _zz_dataOut_payload_0_10462;
  wire       [7:0]    _zz_dataOut_payload_0_10463;
  wire                _zz_dataOut_payload_0_10464;
  wire       [7:0]    _zz_dataOut_payload_0_10465;
  wire       [7:0]    _zz_dataOut_payload_0_10466;
  wire                _zz_dataOut_payload_0_10467;
  wire       [7:0]    _zz_dataOut_payload_0_10468;
  wire       [7:0]    _zz_dataOut_payload_0_10469;
  wire                _zz_dataOut_payload_0_10470;
  wire       [7:0]    _zz_dataOut_payload_0_10471;
  wire       [7:0]    _zz_dataOut_payload_0_10472;
  wire                _zz_dataOut_payload_0_10473;
  wire       [7:0]    _zz_dataOut_payload_0_10474;
  wire       [7:0]    _zz_dataOut_payload_0_10475;
  wire                _zz_dataOut_payload_0_10476;
  wire       [7:0]    _zz_dataOut_payload_0_10477;
  wire       [7:0]    _zz_dataOut_payload_0_10478;
  wire                _zz_dataOut_payload_0_10479;
  wire       [7:0]    _zz_dataOut_payload_0_10480;
  wire       [7:0]    _zz_dataOut_payload_0_10481;
  wire                _zz_dataOut_payload_0_10482;
  wire       [7:0]    _zz_dataOut_payload_0_10483;
  wire       [7:0]    _zz_dataOut_payload_0_10484;
  wire                _zz_dataOut_payload_0_10485;
  wire       [7:0]    _zz_dataOut_payload_0_10486;
  wire       [7:0]    _zz_dataOut_payload_0_10487;
  wire                _zz_dataOut_payload_0_10488;
  wire       [7:0]    _zz_dataOut_payload_0_10489;
  wire       [7:0]    _zz_dataOut_payload_0_10490;
  wire                _zz_dataOut_payload_0_10491;
  wire       [7:0]    _zz_dataOut_payload_0_10492;
  wire       [7:0]    _zz_dataOut_payload_0_10493;
  wire                _zz_dataOut_payload_0_10494;
  wire       [7:0]    _zz_dataOut_payload_0_10495;
  wire       [7:0]    _zz_dataOut_payload_0_10496;
  wire                _zz_dataOut_payload_0_10497;
  wire       [7:0]    _zz_dataOut_payload_0_10498;
  wire       [7:0]    _zz_dataOut_payload_0_10499;
  wire                _zz_dataOut_payload_0_10500;
  wire       [7:0]    _zz_dataOut_payload_0_10501;
  wire       [7:0]    _zz_dataOut_payload_0_10502;
  wire                _zz_dataOut_payload_0_10503;
  wire       [7:0]    _zz_dataOut_payload_0_10504;
  wire       [7:0]    _zz_dataOut_payload_0_10505;
  wire                _zz_dataOut_payload_0_10506;
  wire                _zz_dataOut_payload_0_10507;
  reg        [7:0]    _zz_dataOut_payload_0_10508;
  reg        [7:0]    _zz_dataOut_payload_0_10509;
  reg        [7:0]    _zz_dataOut_payload_0_10510;
  reg        [7:0]    _zz_dataOut_payload_0_10511;
  wire                _zz_dataOut_payload_0_10512;
  wire       [7:0]    _zz_dataOut_payload_0_10513;
  wire       [7:0]    _zz_dataOut_payload_0_10514;
  wire                _zz_dataOut_payload_0_10515;
  wire       [7:0]    _zz_dataOut_payload_0_10516;
  wire       [7:0]    _zz_dataOut_payload_0_10517;
  wire                _zz_dataOut_payload_0_10518;
  wire                _zz_dataOut_payload_0_10519;
  reg        [7:0]    _zz_dataOut_payload_0_10520;
  reg        [7:0]    _zz_dataOut_payload_0_10521;
  reg        [7:0]    _zz_dataOut_payload_0_10522;
  reg        [7:0]    _zz_dataOut_payload_0_10523;
  reg        [7:0]    _zz_dataOut_payload_0_10524;
  reg        [7:0]    _zz_dataOut_payload_0_10525;
  reg        [7:0]    _zz_dataOut_payload_0_10526;
  reg        [7:0]    _zz_dataOut_payload_0_10527;
  reg        [7:0]    _zz_dataOut_payload_0_10528;
  reg        [7:0]    _zz_dataOut_payload_0_10529;
  reg        [7:0]    _zz_dataOut_payload_0_10530;
  reg        [7:0]    _zz_dataOut_payload_0_10531;
  wire                _zz_dataOut_payload_0_10532;
  wire       [7:0]    _zz_dataOut_payload_0_10533;
  wire       [7:0]    _zz_dataOut_payload_0_10534;
  wire                _zz_dataOut_payload_0_10535;
  wire       [7:0]    _zz_dataOut_payload_0_10536;
  wire       [7:0]    _zz_dataOut_payload_0_10537;
  wire                _zz_dataOut_payload_0_10538;
  wire       [7:0]    _zz_dataOut_payload_0_10539;
  wire       [7:0]    _zz_dataOut_payload_0_10540;
  wire                _zz_dataOut_payload_0_10541;
  wire       [7:0]    _zz_dataOut_payload_0_10542;
  wire       [7:0]    _zz_dataOut_payload_0_10543;
  wire                _zz_dataOut_payload_0_10544;
  wire       [7:0]    _zz_dataOut_payload_0_10545;
  wire       [7:0]    _zz_dataOut_payload_0_10546;
  wire                _zz_dataOut_payload_0_10547;
  wire       [7:0]    _zz_dataOut_payload_0_10548;
  wire       [7:0]    _zz_dataOut_payload_0_10549;
  wire                _zz_dataOut_payload_0_10550;
  wire                _zz_dataOut_payload_0_10551;
  reg        [7:0]    _zz_dataOut_payload_0_10552;
  reg        [7:0]    _zz_dataOut_payload_0_10553;
  reg        [7:0]    _zz_dataOut_payload_0_10554;
  reg        [7:0]    _zz_dataOut_payload_0_10555;
  wire                _zz_dataOut_payload_0_10556;
  wire       [7:0]    _zz_dataOut_payload_0_10557;
  wire       [7:0]    _zz_dataOut_payload_0_10558;
  wire                _zz_dataOut_payload_0_10559;
  wire       [7:0]    _zz_dataOut_payload_0_10560;
  wire       [7:0]    _zz_dataOut_payload_0_10561;
  wire                _zz_dataOut_payload_0_10562;
  wire                _zz_dataOut_payload_0_10563;
  reg        [7:0]    _zz_dataOut_payload_0_10564;
  reg        [7:0]    _zz_dataOut_payload_0_10565;
  reg        [7:0]    _zz_dataOut_payload_0_10566;
  reg        [7:0]    _zz_dataOut_payload_0_10567;
  reg        [7:0]    _zz_dataOut_payload_0_10568;
  reg        [7:0]    _zz_dataOut_payload_0_10569;
  reg        [7:0]    _zz_dataOut_payload_0_10570;
  reg        [7:0]    _zz_dataOut_payload_0_10571;
  reg        [7:0]    _zz_dataOut_payload_0_10572;
  reg        [7:0]    _zz_dataOut_payload_0_10573;
  reg        [7:0]    _zz_dataOut_payload_0_10574;
  reg        [7:0]    _zz_dataOut_payload_0_10575;
  reg        [7:0]    _zz_dataOut_payload_0_10576;
  reg        [7:0]    _zz_dataOut_payload_0_10577;
  reg        [7:0]    _zz_dataOut_payload_0_10578;
  reg        [7:0]    _zz_dataOut_payload_0_10579;
  reg        [7:0]    _zz_dataOut_payload_0_10580;
  reg        [7:0]    _zz_dataOut_payload_0_10581;
  reg        [7:0]    _zz_dataOut_payload_0_10582;
  reg        [7:0]    _zz_dataOut_payload_0_10583;
  reg        [7:0]    _zz_dataOut_payload_0_10584;
  reg        [7:0]    _zz_dataOut_payload_0_10585;
  reg        [7:0]    _zz_dataOut_payload_0_10586;
  reg        [7:0]    _zz_dataOut_payload_0_10587;
  reg        [7:0]    _zz_dataOut_payload_0_10588;
  reg        [7:0]    _zz_dataOut_payload_0_10589;
  reg        [7:0]    _zz_dataOut_payload_0_10590;
  reg        [7:0]    _zz_dataOut_payload_0_10591;
  wire                _zz_dataOut_payload_0_10592;
  wire       [7:0]    _zz_dataOut_payload_0_10593;
  wire       [7:0]    _zz_dataOut_payload_0_10594;
  wire                _zz_dataOut_payload_0_10595;
  wire       [7:0]    _zz_dataOut_payload_0_10596;
  wire       [7:0]    _zz_dataOut_payload_0_10597;
  wire                _zz_dataOut_payload_0_10598;
  wire       [7:0]    _zz_dataOut_payload_0_10599;
  wire       [7:0]    _zz_dataOut_payload_0_10600;
  wire                _zz_dataOut_payload_0_10601;
  wire       [7:0]    _zz_dataOut_payload_0_10602;
  wire       [7:0]    _zz_dataOut_payload_0_10603;
  wire                _zz_dataOut_payload_0_10604;
  wire       [7:0]    _zz_dataOut_payload_0_10605;
  wire       [7:0]    _zz_dataOut_payload_0_10606;
  wire                _zz_dataOut_payload_0_10607;
  wire       [7:0]    _zz_dataOut_payload_0_10608;
  wire       [7:0]    _zz_dataOut_payload_0_10609;
  wire                _zz_dataOut_payload_0_10610;
  wire       [7:0]    _zz_dataOut_payload_0_10611;
  wire       [7:0]    _zz_dataOut_payload_0_10612;
  wire                _zz_dataOut_payload_0_10613;
  wire       [7:0]    _zz_dataOut_payload_0_10614;
  wire       [7:0]    _zz_dataOut_payload_0_10615;
  wire                _zz_dataOut_payload_0_10616;
  wire       [7:0]    _zz_dataOut_payload_0_10617;
  wire       [7:0]    _zz_dataOut_payload_0_10618;
  wire                _zz_dataOut_payload_0_10619;
  wire       [7:0]    _zz_dataOut_payload_0_10620;
  wire       [7:0]    _zz_dataOut_payload_0_10621;
  wire                _zz_dataOut_payload_0_10622;
  wire       [7:0]    _zz_dataOut_payload_0_10623;
  wire       [7:0]    _zz_dataOut_payload_0_10624;
  wire                _zz_dataOut_payload_0_10625;
  wire       [7:0]    _zz_dataOut_payload_0_10626;
  wire       [7:0]    _zz_dataOut_payload_0_10627;
  wire                _zz_dataOut_payload_0_10628;
  wire       [7:0]    _zz_dataOut_payload_0_10629;
  wire       [7:0]    _zz_dataOut_payload_0_10630;
  wire                _zz_dataOut_payload_0_10631;
  wire       [7:0]    _zz_dataOut_payload_0_10632;
  wire       [7:0]    _zz_dataOut_payload_0_10633;
  wire                _zz_dataOut_payload_0_10634;
  wire                _zz_dataOut_payload_0_10635;
  reg        [7:0]    _zz_dataOut_payload_0_10636;
  reg        [7:0]    _zz_dataOut_payload_0_10637;
  reg        [7:0]    _zz_dataOut_payload_0_10638;
  reg        [7:0]    _zz_dataOut_payload_0_10639;
  wire                _zz_dataOut_payload_0_10640;
  wire       [7:0]    _zz_dataOut_payload_0_10641;
  wire       [7:0]    _zz_dataOut_payload_0_10642;
  wire                _zz_dataOut_payload_0_10643;
  wire       [7:0]    _zz_dataOut_payload_0_10644;
  wire       [7:0]    _zz_dataOut_payload_0_10645;
  wire                _zz_dataOut_payload_0_10646;
  wire                _zz_dataOut_payload_0_10647;
  reg        [7:0]    _zz_dataOut_payload_0_10648;
  reg        [7:0]    _zz_dataOut_payload_0_10649;
  reg        [7:0]    _zz_dataOut_payload_0_10650;
  reg        [7:0]    _zz_dataOut_payload_0_10651;
  reg        [7:0]    _zz_dataOut_payload_0_10652;
  reg        [7:0]    _zz_dataOut_payload_0_10653;
  reg        [7:0]    _zz_dataOut_payload_0_10654;
  reg        [7:0]    _zz_dataOut_payload_0_10655;
  reg        [7:0]    _zz_dataOut_payload_0_10656;
  reg        [7:0]    _zz_dataOut_payload_0_10657;
  reg        [7:0]    _zz_dataOut_payload_0_10658;
  reg        [7:0]    _zz_dataOut_payload_0_10659;
  wire                _zz_dataOut_payload_0_10660;
  wire       [7:0]    _zz_dataOut_payload_0_10661;
  wire       [7:0]    _zz_dataOut_payload_0_10662;
  wire                _zz_dataOut_payload_0_10663;
  wire       [7:0]    _zz_dataOut_payload_0_10664;
  wire       [7:0]    _zz_dataOut_payload_0_10665;
  wire                _zz_dataOut_payload_0_10666;
  wire       [7:0]    _zz_dataOut_payload_0_10667;
  wire       [7:0]    _zz_dataOut_payload_0_10668;
  wire                _zz_dataOut_payload_0_10669;
  wire       [7:0]    _zz_dataOut_payload_0_10670;
  wire       [7:0]    _zz_dataOut_payload_0_10671;
  wire                _zz_dataOut_payload_0_10672;
  wire       [7:0]    _zz_dataOut_payload_0_10673;
  wire       [7:0]    _zz_dataOut_payload_0_10674;
  wire                _zz_dataOut_payload_0_10675;
  wire       [7:0]    _zz_dataOut_payload_0_10676;
  wire       [7:0]    _zz_dataOut_payload_0_10677;
  wire                _zz_dataOut_payload_0_10678;
  wire                _zz_dataOut_payload_0_10679;
  reg        [7:0]    _zz_dataOut_payload_0_10680;
  reg        [7:0]    _zz_dataOut_payload_0_10681;
  reg        [7:0]    _zz_dataOut_payload_0_10682;
  reg        [7:0]    _zz_dataOut_payload_0_10683;
  wire                _zz_dataOut_payload_0_10684;
  wire       [7:0]    _zz_dataOut_payload_0_10685;
  wire       [7:0]    _zz_dataOut_payload_0_10686;
  wire                _zz_dataOut_payload_0_10687;
  wire       [7:0]    _zz_dataOut_payload_0_10688;
  wire       [7:0]    _zz_dataOut_payload_0_10689;
  wire                _zz_dataOut_payload_0_10690;
  wire                _zz_dataOut_payload_0_10691;
  reg        [7:0]    _zz_dataOut_payload_0_10692;
  reg        [7:0]    _zz_dataOut_payload_0_10693;
  reg        [7:0]    _zz_dataOut_payload_0_10694;
  reg        [7:0]    _zz_dataOut_payload_0_10695;
  reg        [7:0]    _zz_dataOut_payload_0_10696;
  reg        [7:0]    _zz_dataOut_payload_0_10697;
  reg        [7:0]    _zz_dataOut_payload_0_10698;
  reg        [7:0]    _zz_dataOut_payload_0_10699;
  reg        [7:0]    _zz_dataOut_payload_0_10700;
  reg        [7:0]    _zz_dataOut_payload_0_10701;
  reg        [7:0]    _zz_dataOut_payload_0_10702;
  reg        [7:0]    _zz_dataOut_payload_0_10703;
  reg        [7:0]    _zz_dataOut_payload_0_10704;
  reg        [7:0]    _zz_dataOut_payload_0_10705;
  reg        [7:0]    _zz_dataOut_payload_0_10706;
  reg        [7:0]    _zz_dataOut_payload_0_10707;
  reg        [7:0]    _zz_dataOut_payload_0_10708;
  reg        [7:0]    _zz_dataOut_payload_0_10709;
  reg        [7:0]    _zz_dataOut_payload_0_10710;
  reg        [7:0]    _zz_dataOut_payload_0_10711;
  reg        [7:0]    _zz_dataOut_payload_0_10712;
  reg        [7:0]    _zz_dataOut_payload_0_10713;
  reg        [7:0]    _zz_dataOut_payload_0_10714;
  reg        [7:0]    _zz_dataOut_payload_0_10715;
  reg        [7:0]    _zz_dataOut_payload_0_10716;
  reg        [7:0]    _zz_dataOut_payload_0_10717;
  reg        [7:0]    _zz_dataOut_payload_0_10718;
  reg        [7:0]    _zz_dataOut_payload_0_10719;
  reg        [7:0]    _zz_dataOut_payload_0_10720;
  reg        [7:0]    _zz_dataOut_payload_0_10721;
  reg        [7:0]    _zz_dataOut_payload_0_10722;
  reg        [7:0]    _zz_dataOut_payload_0_10723;
  reg        [7:0]    _zz_dataOut_payload_0_10724;
  reg        [7:0]    _zz_dataOut_payload_0_10725;
  reg        [7:0]    _zz_dataOut_payload_0_10726;
  reg        [7:0]    _zz_dataOut_payload_0_10727;
  reg        [7:0]    _zz_dataOut_payload_0_10728;
  reg        [7:0]    _zz_dataOut_payload_0_10729;
  reg        [7:0]    _zz_dataOut_payload_0_10730;
  reg        [7:0]    _zz_dataOut_payload_0_10731;
  reg        [7:0]    _zz_dataOut_payload_0_10732;
  reg        [7:0]    _zz_dataOut_payload_0_10733;
  reg        [7:0]    _zz_dataOut_payload_0_10734;
  reg        [7:0]    _zz_dataOut_payload_0_10735;
  reg        [7:0]    _zz_dataOut_payload_0_10736;
  reg        [7:0]    _zz_dataOut_payload_0_10737;
  reg        [7:0]    _zz_dataOut_payload_0_10738;
  reg        [7:0]    _zz_dataOut_payload_0_10739;
  reg        [7:0]    _zz_dataOut_payload_0_10740;
  reg        [7:0]    _zz_dataOut_payload_0_10741;
  reg        [7:0]    _zz_dataOut_payload_0_10742;
  reg        [7:0]    _zz_dataOut_payload_0_10743;
  reg        [7:0]    _zz_dataOut_payload_0_10744;
  reg        [7:0]    _zz_dataOut_payload_0_10745;
  reg        [7:0]    _zz_dataOut_payload_0_10746;
  reg        [7:0]    _zz_dataOut_payload_0_10747;
  reg        [7:0]    _zz_dataOut_payload_0_10748;
  reg        [7:0]    _zz_dataOut_payload_0_10749;
  reg        [7:0]    _zz_dataOut_payload_0_10750;
  reg        [7:0]    _zz_dataOut_payload_0_10751;
  reg        [7:0]    _zz_dataOut_payload_0_10752;
  reg        [7:0]    _zz_dataOut_payload_0_10753;
  reg        [7:0]    _zz_dataOut_payload_0_10754;
  reg        [7:0]    _zz_dataOut_payload_0_10755;
  reg        [7:0]    _zz_dataOut_payload_0_10756;
  reg        [7:0]    _zz_dataOut_payload_0_10757;
  reg        [7:0]    _zz_dataOut_payload_0_10758;
  reg        [7:0]    _zz_dataOut_payload_0_10759;
  reg        [7:0]    _zz_dataOut_payload_0_10760;
  reg        [7:0]    _zz_dataOut_payload_0_10761;
  reg        [7:0]    _zz_dataOut_payload_0_10762;
  reg        [7:0]    _zz_dataOut_payload_0_10763;
  reg        [7:0]    _zz_dataOut_payload_0_10764;
  reg        [7:0]    _zz_dataOut_payload_0_10765;
  reg        [7:0]    _zz_dataOut_payload_0_10766;
  reg        [7:0]    _zz_dataOut_payload_0_10767;
  reg        [7:0]    _zz_dataOut_payload_0_10768;
  reg        [7:0]    _zz_dataOut_payload_0_10769;
  reg        [7:0]    _zz_dataOut_payload_0_10770;
  reg        [7:0]    _zz_dataOut_payload_0_10771;
  reg        [7:0]    _zz_dataOut_payload_0_10772;
  reg        [7:0]    _zz_dataOut_payload_0_10773;
  reg        [7:0]    _zz_dataOut_payload_0_10774;
  reg        [7:0]    _zz_dataOut_payload_0_10775;
  reg        [7:0]    _zz_dataOut_payload_0_10776;
  reg        [7:0]    _zz_dataOut_payload_0_10777;
  reg        [7:0]    _zz_dataOut_payload_0_10778;
  reg        [7:0]    _zz_dataOut_payload_0_10779;
  reg        [7:0]    _zz_dataOut_payload_0_10780;
  reg        [7:0]    _zz_dataOut_payload_0_10781;
  reg        [7:0]    _zz_dataOut_payload_0_10782;
  reg        [7:0]    _zz_dataOut_payload_0_10783;
  reg        [7:0]    _zz_dataOut_payload_0_10784;
  reg        [7:0]    _zz_dataOut_payload_0_10785;
  reg        [7:0]    _zz_dataOut_payload_0_10786;
  reg        [7:0]    _zz_dataOut_payload_0_10787;
  reg        [7:0]    _zz_dataOut_payload_0_10788;
  reg        [7:0]    _zz_dataOut_payload_0_10789;
  reg        [7:0]    _zz_dataOut_payload_0_10790;
  reg        [7:0]    _zz_dataOut_payload_0_10791;
  reg        [7:0]    _zz_dataOut_payload_0_10792;
  reg        [7:0]    _zz_dataOut_payload_0_10793;
  reg        [7:0]    _zz_dataOut_payload_0_10794;
  reg        [7:0]    _zz_dataOut_payload_0_10795;
  reg        [7:0]    _zz_dataOut_payload_0_10796;
  reg        [7:0]    _zz_dataOut_payload_0_10797;
  reg        [7:0]    _zz_dataOut_payload_0_10798;
  reg        [7:0]    _zz_dataOut_payload_0_10799;
  reg        [7:0]    _zz_dataOut_payload_0_10800;
  reg        [7:0]    _zz_dataOut_payload_0_10801;
  reg        [7:0]    _zz_dataOut_payload_0_10802;
  reg        [7:0]    _zz_dataOut_payload_0_10803;
  reg        [7:0]    _zz_dataOut_payload_0_10804;
  reg        [7:0]    _zz_dataOut_payload_0_10805;
  reg        [7:0]    _zz_dataOut_payload_0_10806;
  reg        [7:0]    _zz_dataOut_payload_0_10807;
  reg        [7:0]    _zz_dataOut_payload_0_10808;
  reg        [7:0]    _zz_dataOut_payload_0_10809;
  reg        [7:0]    _zz_dataOut_payload_0_10810;
  reg        [7:0]    _zz_dataOut_payload_0_10811;
  reg        [7:0]    _zz_dataOut_payload_0_10812;
  reg        [7:0]    _zz_dataOut_payload_0_10813;
  reg        [7:0]    _zz_dataOut_payload_0_10814;
  reg        [7:0]    _zz_dataOut_payload_0_10815;
  wire                _zz_dataOut_payload_0_10816;
  wire       [7:0]    _zz_dataOut_payload_0_10817;
  wire       [7:0]    _zz_dataOut_payload_0_10818;
  wire                _zz_dataOut_payload_0_10819;
  wire       [7:0]    _zz_dataOut_payload_0_10820;
  wire       [7:0]    _zz_dataOut_payload_0_10821;
  wire                _zz_dataOut_payload_0_10822;
  wire       [7:0]    _zz_dataOut_payload_0_10823;
  wire       [7:0]    _zz_dataOut_payload_0_10824;
  wire                _zz_dataOut_payload_0_10825;
  wire       [7:0]    _zz_dataOut_payload_0_10826;
  wire       [7:0]    _zz_dataOut_payload_0_10827;
  wire                _zz_dataOut_payload_0_10828;
  wire       [7:0]    _zz_dataOut_payload_0_10829;
  wire       [7:0]    _zz_dataOut_payload_0_10830;
  wire                _zz_dataOut_payload_0_10831;
  wire       [7:0]    _zz_dataOut_payload_0_10832;
  wire       [7:0]    _zz_dataOut_payload_0_10833;
  wire                _zz_dataOut_payload_0_10834;
  wire       [7:0]    _zz_dataOut_payload_0_10835;
  wire       [7:0]    _zz_dataOut_payload_0_10836;
  wire                _zz_dataOut_payload_0_10837;
  wire       [7:0]    _zz_dataOut_payload_0_10838;
  wire       [7:0]    _zz_dataOut_payload_0_10839;
  wire                _zz_dataOut_payload_0_10840;
  wire       [7:0]    _zz_dataOut_payload_0_10841;
  wire       [7:0]    _zz_dataOut_payload_0_10842;
  wire                _zz_dataOut_payload_0_10843;
  wire       [7:0]    _zz_dataOut_payload_0_10844;
  wire       [7:0]    _zz_dataOut_payload_0_10845;
  wire                _zz_dataOut_payload_0_10846;
  wire       [7:0]    _zz_dataOut_payload_0_10847;
  wire       [7:0]    _zz_dataOut_payload_0_10848;
  wire                _zz_dataOut_payload_0_10849;
  wire       [7:0]    _zz_dataOut_payload_0_10850;
  wire       [7:0]    _zz_dataOut_payload_0_10851;
  wire                _zz_dataOut_payload_0_10852;
  wire       [7:0]    _zz_dataOut_payload_0_10853;
  wire       [7:0]    _zz_dataOut_payload_0_10854;
  wire                _zz_dataOut_payload_0_10855;
  wire       [7:0]    _zz_dataOut_payload_0_10856;
  wire       [7:0]    _zz_dataOut_payload_0_10857;
  wire                _zz_dataOut_payload_0_10858;
  wire       [7:0]    _zz_dataOut_payload_0_10859;
  wire       [7:0]    _zz_dataOut_payload_0_10860;
  wire                _zz_dataOut_payload_0_10861;
  wire       [7:0]    _zz_dataOut_payload_0_10862;
  wire       [7:0]    _zz_dataOut_payload_0_10863;
  wire                _zz_dataOut_payload_0_10864;
  wire       [7:0]    _zz_dataOut_payload_0_10865;
  wire       [7:0]    _zz_dataOut_payload_0_10866;
  wire                _zz_dataOut_payload_0_10867;
  wire       [7:0]    _zz_dataOut_payload_0_10868;
  wire       [7:0]    _zz_dataOut_payload_0_10869;
  wire                _zz_dataOut_payload_0_10870;
  wire       [7:0]    _zz_dataOut_payload_0_10871;
  wire       [7:0]    _zz_dataOut_payload_0_10872;
  wire                _zz_dataOut_payload_0_10873;
  wire       [7:0]    _zz_dataOut_payload_0_10874;
  wire       [7:0]    _zz_dataOut_payload_0_10875;
  wire                _zz_dataOut_payload_0_10876;
  wire       [7:0]    _zz_dataOut_payload_0_10877;
  wire       [7:0]    _zz_dataOut_payload_0_10878;
  wire                _zz_dataOut_payload_0_10879;
  wire       [7:0]    _zz_dataOut_payload_0_10880;
  wire       [7:0]    _zz_dataOut_payload_0_10881;
  wire                _zz_dataOut_payload_0_10882;
  wire       [7:0]    _zz_dataOut_payload_0_10883;
  wire       [7:0]    _zz_dataOut_payload_0_10884;
  wire                _zz_dataOut_payload_0_10885;
  wire       [7:0]    _zz_dataOut_payload_0_10886;
  wire       [7:0]    _zz_dataOut_payload_0_10887;
  wire                _zz_dataOut_payload_0_10888;
  wire       [7:0]    _zz_dataOut_payload_0_10889;
  wire       [7:0]    _zz_dataOut_payload_0_10890;
  wire                _zz_dataOut_payload_0_10891;
  wire       [7:0]    _zz_dataOut_payload_0_10892;
  wire       [7:0]    _zz_dataOut_payload_0_10893;
  wire                _zz_dataOut_payload_0_10894;
  wire       [7:0]    _zz_dataOut_payload_0_10895;
  wire       [7:0]    _zz_dataOut_payload_0_10896;
  wire                _zz_dataOut_payload_0_10897;
  wire       [7:0]    _zz_dataOut_payload_0_10898;
  wire       [7:0]    _zz_dataOut_payload_0_10899;
  wire                _zz_dataOut_payload_0_10900;
  wire       [7:0]    _zz_dataOut_payload_0_10901;
  wire       [7:0]    _zz_dataOut_payload_0_10902;
  wire                _zz_dataOut_payload_0_10903;
  wire       [7:0]    _zz_dataOut_payload_0_10904;
  wire       [7:0]    _zz_dataOut_payload_0_10905;
  wire                _zz_dataOut_payload_0_10906;
  wire       [7:0]    _zz_dataOut_payload_0_10907;
  wire       [7:0]    _zz_dataOut_payload_0_10908;
  wire                _zz_dataOut_payload_0_10909;
  wire       [7:0]    _zz_dataOut_payload_0_10910;
  wire       [7:0]    _zz_dataOut_payload_0_10911;
  wire                _zz_dataOut_payload_0_10912;
  wire       [7:0]    _zz_dataOut_payload_0_10913;
  wire       [7:0]    _zz_dataOut_payload_0_10914;
  wire                _zz_dataOut_payload_0_10915;
  wire       [7:0]    _zz_dataOut_payload_0_10916;
  wire       [7:0]    _zz_dataOut_payload_0_10917;
  wire                _zz_dataOut_payload_0_10918;
  wire       [7:0]    _zz_dataOut_payload_0_10919;
  wire       [7:0]    _zz_dataOut_payload_0_10920;
  wire                _zz_dataOut_payload_0_10921;
  wire       [7:0]    _zz_dataOut_payload_0_10922;
  wire       [7:0]    _zz_dataOut_payload_0_10923;
  wire                _zz_dataOut_payload_0_10924;
  wire       [7:0]    _zz_dataOut_payload_0_10925;
  wire       [7:0]    _zz_dataOut_payload_0_10926;
  wire                _zz_dataOut_payload_0_10927;
  wire       [7:0]    _zz_dataOut_payload_0_10928;
  wire       [7:0]    _zz_dataOut_payload_0_10929;
  wire                _zz_dataOut_payload_0_10930;
  wire       [7:0]    _zz_dataOut_payload_0_10931;
  wire       [7:0]    _zz_dataOut_payload_0_10932;
  wire                _zz_dataOut_payload_0_10933;
  wire       [7:0]    _zz_dataOut_payload_0_10934;
  wire       [7:0]    _zz_dataOut_payload_0_10935;
  wire                _zz_dataOut_payload_0_10936;
  wire       [7:0]    _zz_dataOut_payload_0_10937;
  wire       [7:0]    _zz_dataOut_payload_0_10938;
  wire                _zz_dataOut_payload_0_10939;
  wire       [7:0]    _zz_dataOut_payload_0_10940;
  wire       [7:0]    _zz_dataOut_payload_0_10941;
  wire                _zz_dataOut_payload_0_10942;
  wire       [7:0]    _zz_dataOut_payload_0_10943;
  wire       [7:0]    _zz_dataOut_payload_0_10944;
  wire                _zz_dataOut_payload_0_10945;
  wire       [7:0]    _zz_dataOut_payload_0_10946;
  wire       [7:0]    _zz_dataOut_payload_0_10947;
  wire                _zz_dataOut_payload_0_10948;
  wire       [7:0]    _zz_dataOut_payload_0_10949;
  wire       [7:0]    _zz_dataOut_payload_0_10950;
  wire                _zz_dataOut_payload_0_10951;
  wire       [7:0]    _zz_dataOut_payload_0_10952;
  wire       [7:0]    _zz_dataOut_payload_0_10953;
  wire                _zz_dataOut_payload_0_10954;
  wire       [7:0]    _zz_dataOut_payload_0_10955;
  wire       [7:0]    _zz_dataOut_payload_0_10956;
  wire                _zz_dataOut_payload_0_10957;
  wire       [7:0]    _zz_dataOut_payload_0_10958;
  wire       [7:0]    _zz_dataOut_payload_0_10959;
  wire                _zz_dataOut_payload_0_10960;
  wire       [7:0]    _zz_dataOut_payload_0_10961;
  wire       [7:0]    _zz_dataOut_payload_0_10962;
  wire                _zz_dataOut_payload_0_10963;
  wire       [7:0]    _zz_dataOut_payload_0_10964;
  wire       [7:0]    _zz_dataOut_payload_0_10965;
  wire                _zz_dataOut_payload_0_10966;
  wire       [7:0]    _zz_dataOut_payload_0_10967;
  wire       [7:0]    _zz_dataOut_payload_0_10968;
  wire                _zz_dataOut_payload_0_10969;
  wire       [7:0]    _zz_dataOut_payload_0_10970;
  wire       [7:0]    _zz_dataOut_payload_0_10971;
  wire                _zz_dataOut_payload_0_10972;
  wire       [7:0]    _zz_dataOut_payload_0_10973;
  wire       [7:0]    _zz_dataOut_payload_0_10974;
  wire                _zz_dataOut_payload_0_10975;
  wire       [7:0]    _zz_dataOut_payload_0_10976;
  wire       [7:0]    _zz_dataOut_payload_0_10977;
  wire                _zz_dataOut_payload_0_10978;
  wire       [7:0]    _zz_dataOut_payload_0_10979;
  wire       [7:0]    _zz_dataOut_payload_0_10980;
  wire                _zz_dataOut_payload_0_10981;
  wire       [7:0]    _zz_dataOut_payload_0_10982;
  wire       [7:0]    _zz_dataOut_payload_0_10983;
  wire                _zz_dataOut_payload_0_10984;
  wire       [7:0]    _zz_dataOut_payload_0_10985;
  wire       [7:0]    _zz_dataOut_payload_0_10986;
  wire                _zz_dataOut_payload_0_10987;
  wire       [7:0]    _zz_dataOut_payload_0_10988;
  wire       [7:0]    _zz_dataOut_payload_0_10989;
  wire                _zz_dataOut_payload_0_10990;
  wire       [7:0]    _zz_dataOut_payload_0_10991;
  wire       [7:0]    _zz_dataOut_payload_0_10992;
  wire                _zz_dataOut_payload_0_10993;
  wire       [7:0]    _zz_dataOut_payload_0_10994;
  wire       [7:0]    _zz_dataOut_payload_0_10995;
  wire                _zz_dataOut_payload_0_10996;
  wire       [7:0]    _zz_dataOut_payload_0_10997;
  wire       [7:0]    _zz_dataOut_payload_0_10998;
  wire                _zz_dataOut_payload_0_10999;
  wire       [7:0]    _zz_dataOut_payload_0_11000;
  wire       [7:0]    _zz_dataOut_payload_0_11001;
  wire                _zz_dataOut_payload_0_11002;
  wire                _zz_dataOut_payload_0_11003;
  reg        [7:0]    _zz_dataOut_payload_0_11004;
  reg        [7:0]    _zz_dataOut_payload_0_11005;
  reg        [7:0]    _zz_dataOut_payload_0_11006;
  reg        [7:0]    _zz_dataOut_payload_0_11007;
  wire                _zz_dataOut_payload_0_11008;
  wire       [7:0]    _zz_dataOut_payload_0_11009;
  wire       [7:0]    _zz_dataOut_payload_0_11010;
  wire                _zz_dataOut_payload_0_11011;
  wire       [7:0]    _zz_dataOut_payload_0_11012;
  wire       [7:0]    _zz_dataOut_payload_0_11013;
  wire                _zz_dataOut_payload_0_11014;
  wire                _zz_dataOut_payload_0_11015;
  reg        [7:0]    _zz_dataOut_payload_0_11016;
  reg        [7:0]    _zz_dataOut_payload_0_11017;
  reg        [7:0]    _zz_dataOut_payload_0_11018;
  reg        [7:0]    _zz_dataOut_payload_0_11019;
  reg        [7:0]    _zz_dataOut_payload_0_11020;
  reg        [7:0]    _zz_dataOut_payload_0_11021;
  reg        [7:0]    _zz_dataOut_payload_0_11022;
  reg        [7:0]    _zz_dataOut_payload_0_11023;
  reg        [7:0]    _zz_dataOut_payload_0_11024;
  reg        [7:0]    _zz_dataOut_payload_0_11025;
  reg        [7:0]    _zz_dataOut_payload_0_11026;
  reg        [7:0]    _zz_dataOut_payload_0_11027;
  wire                _zz_dataOut_payload_0_11028;
  wire       [7:0]    _zz_dataOut_payload_0_11029;
  wire       [7:0]    _zz_dataOut_payload_0_11030;
  wire                _zz_dataOut_payload_0_11031;
  wire       [7:0]    _zz_dataOut_payload_0_11032;
  wire       [7:0]    _zz_dataOut_payload_0_11033;
  wire                _zz_dataOut_payload_0_11034;
  wire       [7:0]    _zz_dataOut_payload_0_11035;
  wire       [7:0]    _zz_dataOut_payload_0_11036;
  wire                _zz_dataOut_payload_0_11037;
  wire       [7:0]    _zz_dataOut_payload_0_11038;
  wire       [7:0]    _zz_dataOut_payload_0_11039;
  wire                _zz_dataOut_payload_0_11040;
  wire       [7:0]    _zz_dataOut_payload_0_11041;
  wire       [7:0]    _zz_dataOut_payload_0_11042;
  wire                _zz_dataOut_payload_0_11043;
  wire       [7:0]    _zz_dataOut_payload_0_11044;
  wire       [7:0]    _zz_dataOut_payload_0_11045;
  wire                _zz_dataOut_payload_0_11046;
  wire                _zz_dataOut_payload_0_11047;
  reg        [7:0]    _zz_dataOut_payload_0_11048;
  reg        [7:0]    _zz_dataOut_payload_0_11049;
  reg        [7:0]    _zz_dataOut_payload_0_11050;
  reg        [7:0]    _zz_dataOut_payload_0_11051;
  wire                _zz_dataOut_payload_0_11052;
  wire       [7:0]    _zz_dataOut_payload_0_11053;
  wire       [7:0]    _zz_dataOut_payload_0_11054;
  wire                _zz_dataOut_payload_0_11055;
  wire       [7:0]    _zz_dataOut_payload_0_11056;
  wire       [7:0]    _zz_dataOut_payload_0_11057;
  wire                _zz_dataOut_payload_0_11058;
  wire                _zz_dataOut_payload_0_11059;
  reg        [7:0]    _zz_dataOut_payload_0_11060;
  reg        [7:0]    _zz_dataOut_payload_0_11061;
  reg        [7:0]    _zz_dataOut_payload_0_11062;
  reg        [7:0]    _zz_dataOut_payload_0_11063;
  reg        [7:0]    _zz_dataOut_payload_0_11064;
  reg        [7:0]    _zz_dataOut_payload_0_11065;
  reg        [7:0]    _zz_dataOut_payload_0_11066;
  reg        [7:0]    _zz_dataOut_payload_0_11067;
  reg        [7:0]    _zz_dataOut_payload_0_11068;
  reg        [7:0]    _zz_dataOut_payload_0_11069;
  reg        [7:0]    _zz_dataOut_payload_0_11070;
  reg        [7:0]    _zz_dataOut_payload_0_11071;
  reg        [7:0]    _zz_dataOut_payload_0_11072;
  reg        [7:0]    _zz_dataOut_payload_0_11073;
  reg        [7:0]    _zz_dataOut_payload_0_11074;
  reg        [7:0]    _zz_dataOut_payload_0_11075;
  reg        [7:0]    _zz_dataOut_payload_0_11076;
  reg        [7:0]    _zz_dataOut_payload_0_11077;
  reg        [7:0]    _zz_dataOut_payload_0_11078;
  reg        [7:0]    _zz_dataOut_payload_0_11079;
  reg        [7:0]    _zz_dataOut_payload_0_11080;
  reg        [7:0]    _zz_dataOut_payload_0_11081;
  reg        [7:0]    _zz_dataOut_payload_0_11082;
  reg        [7:0]    _zz_dataOut_payload_0_11083;
  reg        [7:0]    _zz_dataOut_payload_0_11084;
  reg        [7:0]    _zz_dataOut_payload_0_11085;
  reg        [7:0]    _zz_dataOut_payload_0_11086;
  reg        [7:0]    _zz_dataOut_payload_0_11087;
  wire                _zz_dataOut_payload_0_11088;
  wire       [7:0]    _zz_dataOut_payload_0_11089;
  wire       [7:0]    _zz_dataOut_payload_0_11090;
  wire                _zz_dataOut_payload_0_11091;
  wire       [7:0]    _zz_dataOut_payload_0_11092;
  wire       [7:0]    _zz_dataOut_payload_0_11093;
  wire                _zz_dataOut_payload_0_11094;
  wire       [7:0]    _zz_dataOut_payload_0_11095;
  wire       [7:0]    _zz_dataOut_payload_0_11096;
  wire                _zz_dataOut_payload_0_11097;
  wire       [7:0]    _zz_dataOut_payload_0_11098;
  wire       [7:0]    _zz_dataOut_payload_0_11099;
  wire                _zz_dataOut_payload_0_11100;
  wire       [7:0]    _zz_dataOut_payload_0_11101;
  wire       [7:0]    _zz_dataOut_payload_0_11102;
  wire                _zz_dataOut_payload_0_11103;
  wire       [7:0]    _zz_dataOut_payload_0_11104;
  wire       [7:0]    _zz_dataOut_payload_0_11105;
  wire                _zz_dataOut_payload_0_11106;
  wire       [7:0]    _zz_dataOut_payload_0_11107;
  wire       [7:0]    _zz_dataOut_payload_0_11108;
  wire                _zz_dataOut_payload_0_11109;
  wire       [7:0]    _zz_dataOut_payload_0_11110;
  wire       [7:0]    _zz_dataOut_payload_0_11111;
  wire                _zz_dataOut_payload_0_11112;
  wire       [7:0]    _zz_dataOut_payload_0_11113;
  wire       [7:0]    _zz_dataOut_payload_0_11114;
  wire                _zz_dataOut_payload_0_11115;
  wire       [7:0]    _zz_dataOut_payload_0_11116;
  wire       [7:0]    _zz_dataOut_payload_0_11117;
  wire                _zz_dataOut_payload_0_11118;
  wire       [7:0]    _zz_dataOut_payload_0_11119;
  wire       [7:0]    _zz_dataOut_payload_0_11120;
  wire                _zz_dataOut_payload_0_11121;
  wire       [7:0]    _zz_dataOut_payload_0_11122;
  wire       [7:0]    _zz_dataOut_payload_0_11123;
  wire                _zz_dataOut_payload_0_11124;
  wire       [7:0]    _zz_dataOut_payload_0_11125;
  wire       [7:0]    _zz_dataOut_payload_0_11126;
  wire                _zz_dataOut_payload_0_11127;
  wire       [7:0]    _zz_dataOut_payload_0_11128;
  wire       [7:0]    _zz_dataOut_payload_0_11129;
  wire                _zz_dataOut_payload_0_11130;
  wire                _zz_dataOut_payload_0_11131;
  reg        [7:0]    _zz_dataOut_payload_0_11132;
  reg        [7:0]    _zz_dataOut_payload_0_11133;
  reg        [7:0]    _zz_dataOut_payload_0_11134;
  reg        [7:0]    _zz_dataOut_payload_0_11135;
  wire                _zz_dataOut_payload_0_11136;
  wire       [7:0]    _zz_dataOut_payload_0_11137;
  wire       [7:0]    _zz_dataOut_payload_0_11138;
  wire                _zz_dataOut_payload_0_11139;
  wire       [7:0]    _zz_dataOut_payload_0_11140;
  wire       [7:0]    _zz_dataOut_payload_0_11141;
  wire                _zz_dataOut_payload_0_11142;
  wire                _zz_dataOut_payload_0_11143;
  reg        [7:0]    _zz_dataOut_payload_0_11144;
  reg        [7:0]    _zz_dataOut_payload_0_11145;
  reg        [7:0]    _zz_dataOut_payload_0_11146;
  reg        [7:0]    _zz_dataOut_payload_0_11147;
  reg        [7:0]    _zz_dataOut_payload_0_11148;
  reg        [7:0]    _zz_dataOut_payload_0_11149;
  reg        [7:0]    _zz_dataOut_payload_0_11150;
  reg        [7:0]    _zz_dataOut_payload_0_11151;
  reg        [7:0]    _zz_dataOut_payload_0_11152;
  reg        [7:0]    _zz_dataOut_payload_0_11153;
  reg        [7:0]    _zz_dataOut_payload_0_11154;
  reg        [7:0]    _zz_dataOut_payload_0_11155;
  wire                _zz_dataOut_payload_0_11156;
  wire       [7:0]    _zz_dataOut_payload_0_11157;
  wire       [7:0]    _zz_dataOut_payload_0_11158;
  wire                _zz_dataOut_payload_0_11159;
  wire       [7:0]    _zz_dataOut_payload_0_11160;
  wire       [7:0]    _zz_dataOut_payload_0_11161;
  wire                _zz_dataOut_payload_0_11162;
  wire       [7:0]    _zz_dataOut_payload_0_11163;
  wire       [7:0]    _zz_dataOut_payload_0_11164;
  wire                _zz_dataOut_payload_0_11165;
  wire       [7:0]    _zz_dataOut_payload_0_11166;
  wire       [7:0]    _zz_dataOut_payload_0_11167;
  wire                _zz_dataOut_payload_0_11168;
  wire       [7:0]    _zz_dataOut_payload_0_11169;
  wire       [7:0]    _zz_dataOut_payload_0_11170;
  wire                _zz_dataOut_payload_0_11171;
  wire       [7:0]    _zz_dataOut_payload_0_11172;
  wire       [7:0]    _zz_dataOut_payload_0_11173;
  wire                _zz_dataOut_payload_0_11174;
  wire                _zz_dataOut_payload_0_11175;
  reg        [7:0]    _zz_dataOut_payload_0_11176;
  reg        [7:0]    _zz_dataOut_payload_0_11177;
  reg        [7:0]    _zz_dataOut_payload_0_11178;
  reg        [7:0]    _zz_dataOut_payload_0_11179;
  wire                _zz_dataOut_payload_0_11180;
  wire       [7:0]    _zz_dataOut_payload_0_11181;
  wire       [7:0]    _zz_dataOut_payload_0_11182;
  wire                _zz_dataOut_payload_0_11183;
  wire       [7:0]    _zz_dataOut_payload_0_11184;
  wire       [7:0]    _zz_dataOut_payload_0_11185;
  wire                _zz_dataOut_payload_0_11186;
  wire                _zz_dataOut_payload_0_11187;
  reg        [7:0]    _zz_dataOut_payload_0_11188;
  reg        [7:0]    _zz_dataOut_payload_0_11189;
  reg        [7:0]    _zz_dataOut_payload_0_11190;
  reg        [7:0]    _zz_dataOut_payload_0_11191;
  reg        [7:0]    _zz_dataOut_payload_0_11192;
  reg        [7:0]    _zz_dataOut_payload_0_11193;
  reg        [7:0]    _zz_dataOut_payload_0_11194;
  reg        [7:0]    _zz_dataOut_payload_0_11195;
  reg        [7:0]    _zz_dataOut_payload_0_11196;
  reg        [7:0]    _zz_dataOut_payload_0_11197;
  reg        [7:0]    _zz_dataOut_payload_0_11198;
  reg        [7:0]    _zz_dataOut_payload_0_11199;
  reg        [7:0]    _zz_dataOut_payload_0_11200;
  reg        [7:0]    _zz_dataOut_payload_0_11201;
  reg        [7:0]    _zz_dataOut_payload_0_11202;
  reg        [7:0]    _zz_dataOut_payload_0_11203;
  reg        [7:0]    _zz_dataOut_payload_0_11204;
  reg        [7:0]    _zz_dataOut_payload_0_11205;
  reg        [7:0]    _zz_dataOut_payload_0_11206;
  reg        [7:0]    _zz_dataOut_payload_0_11207;
  reg        [7:0]    _zz_dataOut_payload_0_11208;
  reg        [7:0]    _zz_dataOut_payload_0_11209;
  reg        [7:0]    _zz_dataOut_payload_0_11210;
  reg        [7:0]    _zz_dataOut_payload_0_11211;
  reg        [7:0]    _zz_dataOut_payload_0_11212;
  reg        [7:0]    _zz_dataOut_payload_0_11213;
  reg        [7:0]    _zz_dataOut_payload_0_11214;
  reg        [7:0]    _zz_dataOut_payload_0_11215;
  reg        [7:0]    _zz_dataOut_payload_0_11216;
  reg        [7:0]    _zz_dataOut_payload_0_11217;
  reg        [7:0]    _zz_dataOut_payload_0_11218;
  reg        [7:0]    _zz_dataOut_payload_0_11219;
  reg        [7:0]    _zz_dataOut_payload_0_11220;
  reg        [7:0]    _zz_dataOut_payload_0_11221;
  reg        [7:0]    _zz_dataOut_payload_0_11222;
  reg        [7:0]    _zz_dataOut_payload_0_11223;
  reg        [7:0]    _zz_dataOut_payload_0_11224;
  reg        [7:0]    _zz_dataOut_payload_0_11225;
  reg        [7:0]    _zz_dataOut_payload_0_11226;
  reg        [7:0]    _zz_dataOut_payload_0_11227;
  reg        [7:0]    _zz_dataOut_payload_0_11228;
  reg        [7:0]    _zz_dataOut_payload_0_11229;
  reg        [7:0]    _zz_dataOut_payload_0_11230;
  reg        [7:0]    _zz_dataOut_payload_0_11231;
  reg        [7:0]    _zz_dataOut_payload_0_11232;
  reg        [7:0]    _zz_dataOut_payload_0_11233;
  reg        [7:0]    _zz_dataOut_payload_0_11234;
  reg        [7:0]    _zz_dataOut_payload_0_11235;
  reg        [7:0]    _zz_dataOut_payload_0_11236;
  reg        [7:0]    _zz_dataOut_payload_0_11237;
  reg        [7:0]    _zz_dataOut_payload_0_11238;
  reg        [7:0]    _zz_dataOut_payload_0_11239;
  reg        [7:0]    _zz_dataOut_payload_0_11240;
  reg        [7:0]    _zz_dataOut_payload_0_11241;
  reg        [7:0]    _zz_dataOut_payload_0_11242;
  reg        [7:0]    _zz_dataOut_payload_0_11243;
  reg        [7:0]    _zz_dataOut_payload_0_11244;
  reg        [7:0]    _zz_dataOut_payload_0_11245;
  reg        [7:0]    _zz_dataOut_payload_0_11246;
  reg        [7:0]    _zz_dataOut_payload_0_11247;
  wire                _zz_dataOut_payload_0_11248;
  wire       [7:0]    _zz_dataOut_payload_0_11249;
  wire       [7:0]    _zz_dataOut_payload_0_11250;
  wire                _zz_dataOut_payload_0_11251;
  wire       [7:0]    _zz_dataOut_payload_0_11252;
  wire       [7:0]    _zz_dataOut_payload_0_11253;
  wire                _zz_dataOut_payload_0_11254;
  wire       [7:0]    _zz_dataOut_payload_0_11255;
  wire       [7:0]    _zz_dataOut_payload_0_11256;
  wire                _zz_dataOut_payload_0_11257;
  wire       [7:0]    _zz_dataOut_payload_0_11258;
  wire       [7:0]    _zz_dataOut_payload_0_11259;
  wire                _zz_dataOut_payload_0_11260;
  wire       [7:0]    _zz_dataOut_payload_0_11261;
  wire       [7:0]    _zz_dataOut_payload_0_11262;
  wire                _zz_dataOut_payload_0_11263;
  wire       [7:0]    _zz_dataOut_payload_0_11264;
  wire       [7:0]    _zz_dataOut_payload_0_11265;
  wire                _zz_dataOut_payload_0_11266;
  wire       [7:0]    _zz_dataOut_payload_0_11267;
  wire       [7:0]    _zz_dataOut_payload_0_11268;
  wire                _zz_dataOut_payload_0_11269;
  wire       [7:0]    _zz_dataOut_payload_0_11270;
  wire       [7:0]    _zz_dataOut_payload_0_11271;
  wire                _zz_dataOut_payload_0_11272;
  wire       [7:0]    _zz_dataOut_payload_0_11273;
  wire       [7:0]    _zz_dataOut_payload_0_11274;
  wire                _zz_dataOut_payload_0_11275;
  wire       [7:0]    _zz_dataOut_payload_0_11276;
  wire       [7:0]    _zz_dataOut_payload_0_11277;
  wire                _zz_dataOut_payload_0_11278;
  wire       [7:0]    _zz_dataOut_payload_0_11279;
  wire       [7:0]    _zz_dataOut_payload_0_11280;
  wire                _zz_dataOut_payload_0_11281;
  wire       [7:0]    _zz_dataOut_payload_0_11282;
  wire       [7:0]    _zz_dataOut_payload_0_11283;
  wire                _zz_dataOut_payload_0_11284;
  wire       [7:0]    _zz_dataOut_payload_0_11285;
  wire       [7:0]    _zz_dataOut_payload_0_11286;
  wire                _zz_dataOut_payload_0_11287;
  wire       [7:0]    _zz_dataOut_payload_0_11288;
  wire       [7:0]    _zz_dataOut_payload_0_11289;
  wire                _zz_dataOut_payload_0_11290;
  wire       [7:0]    _zz_dataOut_payload_0_11291;
  wire       [7:0]    _zz_dataOut_payload_0_11292;
  wire                _zz_dataOut_payload_0_11293;
  wire       [7:0]    _zz_dataOut_payload_0_11294;
  wire       [7:0]    _zz_dataOut_payload_0_11295;
  wire                _zz_dataOut_payload_0_11296;
  wire       [7:0]    _zz_dataOut_payload_0_11297;
  wire       [7:0]    _zz_dataOut_payload_0_11298;
  wire                _zz_dataOut_payload_0_11299;
  wire       [7:0]    _zz_dataOut_payload_0_11300;
  wire       [7:0]    _zz_dataOut_payload_0_11301;
  wire                _zz_dataOut_payload_0_11302;
  wire       [7:0]    _zz_dataOut_payload_0_11303;
  wire       [7:0]    _zz_dataOut_payload_0_11304;
  wire                _zz_dataOut_payload_0_11305;
  wire       [7:0]    _zz_dataOut_payload_0_11306;
  wire       [7:0]    _zz_dataOut_payload_0_11307;
  wire                _zz_dataOut_payload_0_11308;
  wire       [7:0]    _zz_dataOut_payload_0_11309;
  wire       [7:0]    _zz_dataOut_payload_0_11310;
  wire                _zz_dataOut_payload_0_11311;
  wire       [7:0]    _zz_dataOut_payload_0_11312;
  wire       [7:0]    _zz_dataOut_payload_0_11313;
  wire                _zz_dataOut_payload_0_11314;
  wire       [7:0]    _zz_dataOut_payload_0_11315;
  wire       [7:0]    _zz_dataOut_payload_0_11316;
  wire                _zz_dataOut_payload_0_11317;
  wire       [7:0]    _zz_dataOut_payload_0_11318;
  wire       [7:0]    _zz_dataOut_payload_0_11319;
  wire                _zz_dataOut_payload_0_11320;
  wire       [7:0]    _zz_dataOut_payload_0_11321;
  wire       [7:0]    _zz_dataOut_payload_0_11322;
  wire                _zz_dataOut_payload_0_11323;
  wire       [7:0]    _zz_dataOut_payload_0_11324;
  wire       [7:0]    _zz_dataOut_payload_0_11325;
  wire                _zz_dataOut_payload_0_11326;
  wire       [7:0]    _zz_dataOut_payload_0_11327;
  wire       [7:0]    _zz_dataOut_payload_0_11328;
  wire                _zz_dataOut_payload_0_11329;
  wire       [7:0]    _zz_dataOut_payload_0_11330;
  wire       [7:0]    _zz_dataOut_payload_0_11331;
  wire                _zz_dataOut_payload_0_11332;
  wire       [7:0]    _zz_dataOut_payload_0_11333;
  wire       [7:0]    _zz_dataOut_payload_0_11334;
  wire                _zz_dataOut_payload_0_11335;
  wire       [7:0]    _zz_dataOut_payload_0_11336;
  wire       [7:0]    _zz_dataOut_payload_0_11337;
  wire                _zz_dataOut_payload_0_11338;
  wire                _zz_dataOut_payload_0_11339;
  reg        [7:0]    _zz_dataOut_payload_0_11340;
  reg        [7:0]    _zz_dataOut_payload_0_11341;
  reg        [7:0]    _zz_dataOut_payload_0_11342;
  reg        [7:0]    _zz_dataOut_payload_0_11343;
  wire                _zz_dataOut_payload_0_11344;
  wire       [7:0]    _zz_dataOut_payload_0_11345;
  wire       [7:0]    _zz_dataOut_payload_0_11346;
  wire                _zz_dataOut_payload_0_11347;
  wire       [7:0]    _zz_dataOut_payload_0_11348;
  wire       [7:0]    _zz_dataOut_payload_0_11349;
  wire                _zz_dataOut_payload_0_11350;
  wire                _zz_dataOut_payload_0_11351;
  reg        [7:0]    _zz_dataOut_payload_0_11352;
  reg        [7:0]    _zz_dataOut_payload_0_11353;
  reg        [7:0]    _zz_dataOut_payload_0_11354;
  reg        [7:0]    _zz_dataOut_payload_0_11355;
  reg        [7:0]    _zz_dataOut_payload_0_11356;
  reg        [7:0]    _zz_dataOut_payload_0_11357;
  reg        [7:0]    _zz_dataOut_payload_0_11358;
  reg        [7:0]    _zz_dataOut_payload_0_11359;
  reg        [7:0]    _zz_dataOut_payload_0_11360;
  reg        [7:0]    _zz_dataOut_payload_0_11361;
  reg        [7:0]    _zz_dataOut_payload_0_11362;
  reg        [7:0]    _zz_dataOut_payload_0_11363;
  wire                _zz_dataOut_payload_0_11364;
  wire       [7:0]    _zz_dataOut_payload_0_11365;
  wire       [7:0]    _zz_dataOut_payload_0_11366;
  wire                _zz_dataOut_payload_0_11367;
  wire       [7:0]    _zz_dataOut_payload_0_11368;
  wire       [7:0]    _zz_dataOut_payload_0_11369;
  wire                _zz_dataOut_payload_0_11370;
  wire       [7:0]    _zz_dataOut_payload_0_11371;
  wire       [7:0]    _zz_dataOut_payload_0_11372;
  wire                _zz_dataOut_payload_0_11373;
  wire       [7:0]    _zz_dataOut_payload_0_11374;
  wire       [7:0]    _zz_dataOut_payload_0_11375;
  wire                _zz_dataOut_payload_0_11376;
  wire       [7:0]    _zz_dataOut_payload_0_11377;
  wire       [7:0]    _zz_dataOut_payload_0_11378;
  wire                _zz_dataOut_payload_0_11379;
  wire       [7:0]    _zz_dataOut_payload_0_11380;
  wire       [7:0]    _zz_dataOut_payload_0_11381;
  wire                _zz_dataOut_payload_0_11382;
  wire                _zz_dataOut_payload_0_11383;
  reg        [7:0]    _zz_dataOut_payload_0_11384;
  reg        [7:0]    _zz_dataOut_payload_0_11385;
  reg        [7:0]    _zz_dataOut_payload_0_11386;
  reg        [7:0]    _zz_dataOut_payload_0_11387;
  wire                _zz_dataOut_payload_0_11388;
  wire       [7:0]    _zz_dataOut_payload_0_11389;
  wire       [7:0]    _zz_dataOut_payload_0_11390;
  wire                _zz_dataOut_payload_0_11391;
  wire       [7:0]    _zz_dataOut_payload_0_11392;
  wire       [7:0]    _zz_dataOut_payload_0_11393;
  wire                _zz_dataOut_payload_0_11394;
  wire                _zz_dataOut_payload_0_11395;
  reg        [7:0]    _zz_dataOut_payload_0_11396;
  reg        [7:0]    _zz_dataOut_payload_0_11397;
  reg        [7:0]    _zz_dataOut_payload_0_11398;
  reg        [7:0]    _zz_dataOut_payload_0_11399;
  reg        [7:0]    _zz_dataOut_payload_0_11400;
  reg        [7:0]    _zz_dataOut_payload_0_11401;
  reg        [7:0]    _zz_dataOut_payload_0_11402;
  reg        [7:0]    _zz_dataOut_payload_0_11403;
  reg        [7:0]    _zz_dataOut_payload_0_11404;
  reg        [7:0]    _zz_dataOut_payload_0_11405;
  reg        [7:0]    _zz_dataOut_payload_0_11406;
  reg        [7:0]    _zz_dataOut_payload_0_11407;
  reg        [7:0]    _zz_dataOut_payload_0_11408;
  reg        [7:0]    _zz_dataOut_payload_0_11409;
  reg        [7:0]    _zz_dataOut_payload_0_11410;
  reg        [7:0]    _zz_dataOut_payload_0_11411;
  reg        [7:0]    _zz_dataOut_payload_0_11412;
  reg        [7:0]    _zz_dataOut_payload_0_11413;
  reg        [7:0]    _zz_dataOut_payload_0_11414;
  reg        [7:0]    _zz_dataOut_payload_0_11415;
  reg        [7:0]    _zz_dataOut_payload_0_11416;
  reg        [7:0]    _zz_dataOut_payload_0_11417;
  reg        [7:0]    _zz_dataOut_payload_0_11418;
  reg        [7:0]    _zz_dataOut_payload_0_11419;
  reg        [7:0]    _zz_dataOut_payload_0_11420;
  reg        [7:0]    _zz_dataOut_payload_0_11421;
  reg        [7:0]    _zz_dataOut_payload_0_11422;
  reg        [7:0]    _zz_dataOut_payload_0_11423;
  wire                _zz_dataOut_payload_0_11424;
  wire       [7:0]    _zz_dataOut_payload_0_11425;
  wire       [7:0]    _zz_dataOut_payload_0_11426;
  wire                _zz_dataOut_payload_0_11427;
  wire       [7:0]    _zz_dataOut_payload_0_11428;
  wire       [7:0]    _zz_dataOut_payload_0_11429;
  wire                _zz_dataOut_payload_0_11430;
  wire       [7:0]    _zz_dataOut_payload_0_11431;
  wire       [7:0]    _zz_dataOut_payload_0_11432;
  wire                _zz_dataOut_payload_0_11433;
  wire       [7:0]    _zz_dataOut_payload_0_11434;
  wire       [7:0]    _zz_dataOut_payload_0_11435;
  wire                _zz_dataOut_payload_0_11436;
  wire       [7:0]    _zz_dataOut_payload_0_11437;
  wire       [7:0]    _zz_dataOut_payload_0_11438;
  wire                _zz_dataOut_payload_0_11439;
  wire       [7:0]    _zz_dataOut_payload_0_11440;
  wire       [7:0]    _zz_dataOut_payload_0_11441;
  wire                _zz_dataOut_payload_0_11442;
  wire       [7:0]    _zz_dataOut_payload_0_11443;
  wire       [7:0]    _zz_dataOut_payload_0_11444;
  wire                _zz_dataOut_payload_0_11445;
  wire       [7:0]    _zz_dataOut_payload_0_11446;
  wire       [7:0]    _zz_dataOut_payload_0_11447;
  wire                _zz_dataOut_payload_0_11448;
  wire       [7:0]    _zz_dataOut_payload_0_11449;
  wire       [7:0]    _zz_dataOut_payload_0_11450;
  wire                _zz_dataOut_payload_0_11451;
  wire       [7:0]    _zz_dataOut_payload_0_11452;
  wire       [7:0]    _zz_dataOut_payload_0_11453;
  wire                _zz_dataOut_payload_0_11454;
  wire       [7:0]    _zz_dataOut_payload_0_11455;
  wire       [7:0]    _zz_dataOut_payload_0_11456;
  wire                _zz_dataOut_payload_0_11457;
  wire       [7:0]    _zz_dataOut_payload_0_11458;
  wire       [7:0]    _zz_dataOut_payload_0_11459;
  wire                _zz_dataOut_payload_0_11460;
  wire       [7:0]    _zz_dataOut_payload_0_11461;
  wire       [7:0]    _zz_dataOut_payload_0_11462;
  wire                _zz_dataOut_payload_0_11463;
  wire       [7:0]    _zz_dataOut_payload_0_11464;
  wire       [7:0]    _zz_dataOut_payload_0_11465;
  wire                _zz_dataOut_payload_0_11466;
  wire                _zz_dataOut_payload_0_11467;
  reg        [7:0]    _zz_dataOut_payload_0_11468;
  reg        [7:0]    _zz_dataOut_payload_0_11469;
  reg        [7:0]    _zz_dataOut_payload_0_11470;
  reg        [7:0]    _zz_dataOut_payload_0_11471;
  wire                _zz_dataOut_payload_0_11472;
  wire       [7:0]    _zz_dataOut_payload_0_11473;
  wire       [7:0]    _zz_dataOut_payload_0_11474;
  wire                _zz_dataOut_payload_0_11475;
  wire       [7:0]    _zz_dataOut_payload_0_11476;
  wire       [7:0]    _zz_dataOut_payload_0_11477;
  wire                _zz_dataOut_payload_0_11478;
  wire                _zz_dataOut_payload_0_11479;
  reg        [7:0]    _zz_dataOut_payload_0_11480;
  reg        [7:0]    _zz_dataOut_payload_0_11481;
  reg        [7:0]    _zz_dataOut_payload_0_11482;
  reg        [7:0]    _zz_dataOut_payload_0_11483;
  reg        [7:0]    _zz_dataOut_payload_0_11484;
  reg        [7:0]    _zz_dataOut_payload_0_11485;
  reg        [7:0]    _zz_dataOut_payload_0_11486;
  reg        [7:0]    _zz_dataOut_payload_0_11487;
  reg        [7:0]    _zz_dataOut_payload_0_11488;
  reg        [7:0]    _zz_dataOut_payload_0_11489;
  reg        [7:0]    _zz_dataOut_payload_0_11490;
  reg        [7:0]    _zz_dataOut_payload_0_11491;
  wire                _zz_dataOut_payload_0_11492;
  wire       [7:0]    _zz_dataOut_payload_0_11493;
  wire       [7:0]    _zz_dataOut_payload_0_11494;
  wire                _zz_dataOut_payload_0_11495;
  wire       [7:0]    _zz_dataOut_payload_0_11496;
  wire       [7:0]    _zz_dataOut_payload_0_11497;
  wire                _zz_dataOut_payload_0_11498;
  wire       [7:0]    _zz_dataOut_payload_0_11499;
  wire       [7:0]    _zz_dataOut_payload_0_11500;
  wire                _zz_dataOut_payload_0_11501;
  wire       [7:0]    _zz_dataOut_payload_0_11502;
  wire       [7:0]    _zz_dataOut_payload_0_11503;
  wire                _zz_dataOut_payload_0_11504;
  wire       [7:0]    _zz_dataOut_payload_0_11505;
  wire       [7:0]    _zz_dataOut_payload_0_11506;
  wire                _zz_dataOut_payload_0_11507;
  wire       [7:0]    _zz_dataOut_payload_0_11508;
  wire       [7:0]    _zz_dataOut_payload_0_11509;
  wire                _zz_dataOut_payload_0_11510;
  wire                _zz_dataOut_payload_0_11511;
  reg        [7:0]    _zz_dataOut_payload_0_11512;
  reg        [7:0]    _zz_dataOut_payload_0_11513;
  reg        [7:0]    _zz_dataOut_payload_0_11514;
  reg        [7:0]    _zz_dataOut_payload_0_11515;
  wire                _zz_dataOut_payload_0_11516;
  wire       [7:0]    _zz_dataOut_payload_0_11517;
  wire       [7:0]    _zz_dataOut_payload_0_11518;
  wire                _zz_dataOut_payload_0_11519;
  wire       [7:0]    _zz_dataOut_payload_0_11520;
  wire       [7:0]    _zz_dataOut_payload_0_11521;
  wire                _zz_dataOut_payload_0_11522;
  wire                _zz_dataOut_payload_0_11523;
  reg        [7:0]    _zz_dataOut_payload_0_11524;
  reg        [7:0]    _zz_dataOut_payload_0_11525;
  reg        [7:0]    _zz_dataOut_payload_0_11526;
  reg        [7:0]    _zz_dataOut_payload_0_11527;
  reg        [7:0]    _zz_dataOut_payload_0_11528;
  reg        [7:0]    _zz_dataOut_payload_0_11529;
  reg        [7:0]    _zz_dataOut_payload_0_11530;
  reg        [7:0]    _zz_dataOut_payload_0_11531;
  reg        [7:0]    _zz_dataOut_payload_0_11532;
  reg        [7:0]    _zz_dataOut_payload_0_11533;
  reg        [7:0]    _zz_dataOut_payload_0_11534;
  reg        [7:0]    _zz_dataOut_payload_0_11535;
  reg        [7:0]    _zz_dataOut_payload_0_11536;
  reg        [7:0]    _zz_dataOut_payload_0_11537;
  reg        [7:0]    _zz_dataOut_payload_0_11538;
  reg        [7:0]    _zz_dataOut_payload_0_11539;
  reg        [7:0]    _zz_dataOut_payload_0_11540;
  reg        [7:0]    _zz_dataOut_payload_0_11541;
  reg        [7:0]    _zz_dataOut_payload_0_11542;
  reg        [7:0]    _zz_dataOut_payload_0_11543;
  reg        [7:0]    _zz_dataOut_payload_0_11544;
  reg        [7:0]    _zz_dataOut_payload_0_11545;
  reg        [7:0]    _zz_dataOut_payload_0_11546;
  reg        [7:0]    _zz_dataOut_payload_0_11547;
  reg        [7:0]    _zz_dataOut_payload_0_11548;
  reg        [7:0]    _zz_dataOut_payload_0_11549;
  reg        [7:0]    _zz_dataOut_payload_0_11550;
  reg        [7:0]    _zz_dataOut_payload_0_11551;
  reg        [7:0]    _zz_dataOut_payload_0_11552;
  reg        [7:0]    _zz_dataOut_payload_0_11553;
  reg        [7:0]    _zz_dataOut_payload_0_11554;
  reg        [7:0]    _zz_dataOut_payload_0_11555;
  reg        [7:0]    _zz_dataOut_payload_0_11556;
  reg        [7:0]    _zz_dataOut_payload_0_11557;
  reg        [7:0]    _zz_dataOut_payload_0_11558;
  reg        [7:0]    _zz_dataOut_payload_0_11559;
  reg        [7:0]    _zz_dataOut_payload_0_11560;
  reg        [7:0]    _zz_dataOut_payload_0_11561;
  reg        [7:0]    _zz_dataOut_payload_0_11562;
  reg        [7:0]    _zz_dataOut_payload_0_11563;
  reg        [7:0]    _zz_dataOut_payload_0_11564;
  reg        [7:0]    _zz_dataOut_payload_0_11565;
  reg        [7:0]    _zz_dataOut_payload_0_11566;
  reg        [7:0]    _zz_dataOut_payload_0_11567;
  reg        [7:0]    _zz_dataOut_payload_0_11568;
  reg        [7:0]    _zz_dataOut_payload_0_11569;
  reg        [7:0]    _zz_dataOut_payload_0_11570;
  reg        [7:0]    _zz_dataOut_payload_0_11571;
  reg        [7:0]    _zz_dataOut_payload_0_11572;
  reg        [7:0]    _zz_dataOut_payload_0_11573;
  reg        [7:0]    _zz_dataOut_payload_0_11574;
  reg        [7:0]    _zz_dataOut_payload_0_11575;
  reg        [7:0]    _zz_dataOut_payload_0_11576;
  reg        [7:0]    _zz_dataOut_payload_0_11577;
  reg        [7:0]    _zz_dataOut_payload_0_11578;
  reg        [7:0]    _zz_dataOut_payload_0_11579;
  reg        [7:0]    _zz_dataOut_payload_0_11580;
  reg        [7:0]    _zz_dataOut_payload_0_11581;
  reg        [7:0]    _zz_dataOut_payload_0_11582;
  reg        [7:0]    _zz_dataOut_payload_0_11583;
  reg        [7:0]    _zz_dataOut_payload_0_11584;
  reg        [7:0]    _zz_dataOut_payload_0_11585;
  reg        [7:0]    _zz_dataOut_payload_0_11586;
  reg        [7:0]    _zz_dataOut_payload_0_11587;
  reg        [7:0]    _zz_dataOut_payload_0_11588;
  reg        [7:0]    _zz_dataOut_payload_0_11589;
  reg        [7:0]    _zz_dataOut_payload_0_11590;
  reg        [7:0]    _zz_dataOut_payload_0_11591;
  reg        [7:0]    _zz_dataOut_payload_0_11592;
  reg        [7:0]    _zz_dataOut_payload_0_11593;
  reg        [7:0]    _zz_dataOut_payload_0_11594;
  reg        [7:0]    _zz_dataOut_payload_0_11595;
  reg        [7:0]    _zz_dataOut_payload_0_11596;
  reg        [7:0]    _zz_dataOut_payload_0_11597;
  reg        [7:0]    _zz_dataOut_payload_0_11598;
  reg        [7:0]    _zz_dataOut_payload_0_11599;
  reg        [7:0]    _zz_dataOut_payload_0_11600;
  reg        [7:0]    _zz_dataOut_payload_0_11601;
  reg        [7:0]    _zz_dataOut_payload_0_11602;
  reg        [7:0]    _zz_dataOut_payload_0_11603;
  reg        [7:0]    _zz_dataOut_payload_0_11604;
  reg        [7:0]    _zz_dataOut_payload_0_11605;
  reg        [7:0]    _zz_dataOut_payload_0_11606;
  reg        [7:0]    _zz_dataOut_payload_0_11607;
  reg        [7:0]    _zz_dataOut_payload_0_11608;
  reg        [7:0]    _zz_dataOut_payload_0_11609;
  reg        [7:0]    _zz_dataOut_payload_0_11610;
  reg        [7:0]    _zz_dataOut_payload_0_11611;
  reg        [7:0]    _zz_dataOut_payload_0_11612;
  reg        [7:0]    _zz_dataOut_payload_0_11613;
  reg        [7:0]    _zz_dataOut_payload_0_11614;
  reg        [7:0]    _zz_dataOut_payload_0_11615;
  reg        [7:0]    _zz_dataOut_payload_0_11616;
  reg        [7:0]    _zz_dataOut_payload_0_11617;
  reg        [7:0]    _zz_dataOut_payload_0_11618;
  reg        [7:0]    _zz_dataOut_payload_0_11619;
  reg        [7:0]    _zz_dataOut_payload_0_11620;
  reg        [7:0]    _zz_dataOut_payload_0_11621;
  reg        [7:0]    _zz_dataOut_payload_0_11622;
  reg        [7:0]    _zz_dataOut_payload_0_11623;
  reg        [7:0]    _zz_dataOut_payload_0_11624;
  reg        [7:0]    _zz_dataOut_payload_0_11625;
  reg        [7:0]    _zz_dataOut_payload_0_11626;
  reg        [7:0]    _zz_dataOut_payload_0_11627;
  reg        [7:0]    _zz_dataOut_payload_0_11628;
  reg        [7:0]    _zz_dataOut_payload_0_11629;
  reg        [7:0]    _zz_dataOut_payload_0_11630;
  reg        [7:0]    _zz_dataOut_payload_0_11631;
  reg        [7:0]    _zz_dataOut_payload_0_11632;
  reg        [7:0]    _zz_dataOut_payload_0_11633;
  reg        [7:0]    _zz_dataOut_payload_0_11634;
  reg        [7:0]    _zz_dataOut_payload_0_11635;
  reg        [7:0]    _zz_dataOut_payload_0_11636;
  reg        [7:0]    _zz_dataOut_payload_0_11637;
  reg        [7:0]    _zz_dataOut_payload_0_11638;
  reg        [7:0]    _zz_dataOut_payload_0_11639;
  reg        [7:0]    _zz_dataOut_payload_0_11640;
  reg        [7:0]    _zz_dataOut_payload_0_11641;
  reg        [7:0]    _zz_dataOut_payload_0_11642;
  reg        [7:0]    _zz_dataOut_payload_0_11643;
  reg        [7:0]    _zz_dataOut_payload_0_11644;
  reg        [7:0]    _zz_dataOut_payload_0_11645;
  reg        [7:0]    _zz_dataOut_payload_0_11646;
  reg        [7:0]    _zz_dataOut_payload_0_11647;
  reg        [7:0]    _zz_dataOut_payload_0_11648;
  reg        [7:0]    _zz_dataOut_payload_0_11649;
  reg        [7:0]    _zz_dataOut_payload_0_11650;
  reg        [7:0]    _zz_dataOut_payload_0_11651;
  reg        [7:0]    _zz_dataOut_payload_0_11652;
  reg        [7:0]    _zz_dataOut_payload_0_11653;
  reg        [7:0]    _zz_dataOut_payload_0_11654;
  reg        [7:0]    _zz_dataOut_payload_0_11655;
  reg        [7:0]    _zz_dataOut_payload_0_11656;
  reg        [7:0]    _zz_dataOut_payload_0_11657;
  reg        [7:0]    _zz_dataOut_payload_0_11658;
  reg        [7:0]    _zz_dataOut_payload_0_11659;
  reg        [7:0]    _zz_dataOut_payload_0_11660;
  reg        [7:0]    _zz_dataOut_payload_0_11661;
  reg        [7:0]    _zz_dataOut_payload_0_11662;
  reg        [7:0]    _zz_dataOut_payload_0_11663;
  reg        [7:0]    _zz_dataOut_payload_0_11664;
  reg        [7:0]    _zz_dataOut_payload_0_11665;
  reg        [7:0]    _zz_dataOut_payload_0_11666;
  reg        [7:0]    _zz_dataOut_payload_0_11667;
  reg        [7:0]    _zz_dataOut_payload_0_11668;
  reg        [7:0]    _zz_dataOut_payload_0_11669;
  reg        [7:0]    _zz_dataOut_payload_0_11670;
  reg        [7:0]    _zz_dataOut_payload_0_11671;
  reg        [7:0]    _zz_dataOut_payload_0_11672;
  reg        [7:0]    _zz_dataOut_payload_0_11673;
  reg        [7:0]    _zz_dataOut_payload_0_11674;
  reg        [7:0]    _zz_dataOut_payload_0_11675;
  reg        [7:0]    _zz_dataOut_payload_0_11676;
  reg        [7:0]    _zz_dataOut_payload_0_11677;
  reg        [7:0]    _zz_dataOut_payload_0_11678;
  reg        [7:0]    _zz_dataOut_payload_0_11679;
  reg        [7:0]    _zz_dataOut_payload_0_11680;
  reg        [7:0]    _zz_dataOut_payload_0_11681;
  reg        [7:0]    _zz_dataOut_payload_0_11682;
  reg        [7:0]    _zz_dataOut_payload_0_11683;
  reg        [7:0]    _zz_dataOut_payload_0_11684;
  reg        [7:0]    _zz_dataOut_payload_0_11685;
  reg        [7:0]    _zz_dataOut_payload_0_11686;
  reg        [7:0]    _zz_dataOut_payload_0_11687;
  reg        [7:0]    _zz_dataOut_payload_0_11688;
  reg        [7:0]    _zz_dataOut_payload_0_11689;
  reg        [7:0]    _zz_dataOut_payload_0_11690;
  reg        [7:0]    _zz_dataOut_payload_0_11691;
  reg        [7:0]    _zz_dataOut_payload_0_11692;
  reg        [7:0]    _zz_dataOut_payload_0_11693;
  reg        [7:0]    _zz_dataOut_payload_0_11694;
  reg        [7:0]    _zz_dataOut_payload_0_11695;
  reg        [7:0]    _zz_dataOut_payload_0_11696;
  reg        [7:0]    _zz_dataOut_payload_0_11697;
  reg        [7:0]    _zz_dataOut_payload_0_11698;
  reg        [7:0]    _zz_dataOut_payload_0_11699;
  reg        [7:0]    _zz_dataOut_payload_0_11700;
  reg        [7:0]    _zz_dataOut_payload_0_11701;
  reg        [7:0]    _zz_dataOut_payload_0_11702;
  reg        [7:0]    _zz_dataOut_payload_0_11703;
  reg        [7:0]    _zz_dataOut_payload_0_11704;
  reg        [7:0]    _zz_dataOut_payload_0_11705;
  reg        [7:0]    _zz_dataOut_payload_0_11706;
  reg        [7:0]    _zz_dataOut_payload_0_11707;
  reg        [7:0]    _zz_dataOut_payload_0_11708;
  reg        [7:0]    _zz_dataOut_payload_0_11709;
  reg        [7:0]    _zz_dataOut_payload_0_11710;
  reg        [7:0]    _zz_dataOut_payload_0_11711;
  reg        [7:0]    _zz_dataOut_payload_0_11712;
  reg        [7:0]    _zz_dataOut_payload_0_11713;
  reg        [7:0]    _zz_dataOut_payload_0_11714;
  reg        [7:0]    _zz_dataOut_payload_0_11715;
  reg        [7:0]    _zz_dataOut_payload_0_11716;
  reg        [7:0]    _zz_dataOut_payload_0_11717;
  reg        [7:0]    _zz_dataOut_payload_0_11718;
  reg        [7:0]    _zz_dataOut_payload_0_11719;
  reg        [7:0]    _zz_dataOut_payload_0_11720;
  reg        [7:0]    _zz_dataOut_payload_0_11721;
  reg        [7:0]    _zz_dataOut_payload_0_11722;
  reg        [7:0]    _zz_dataOut_payload_0_11723;
  reg        [7:0]    _zz_dataOut_payload_0_11724;
  reg        [7:0]    _zz_dataOut_payload_0_11725;
  reg        [7:0]    _zz_dataOut_payload_0_11726;
  reg        [7:0]    _zz_dataOut_payload_0_11727;
  reg        [7:0]    _zz_dataOut_payload_0_11728;
  reg        [7:0]    _zz_dataOut_payload_0_11729;
  reg        [7:0]    _zz_dataOut_payload_0_11730;
  reg        [7:0]    _zz_dataOut_payload_0_11731;
  reg        [7:0]    _zz_dataOut_payload_0_11732;
  reg        [7:0]    _zz_dataOut_payload_0_11733;
  reg        [7:0]    _zz_dataOut_payload_0_11734;
  reg        [7:0]    _zz_dataOut_payload_0_11735;
  reg        [7:0]    _zz_dataOut_payload_0_11736;
  reg        [7:0]    _zz_dataOut_payload_0_11737;
  reg        [7:0]    _zz_dataOut_payload_0_11738;
  reg        [7:0]    _zz_dataOut_payload_0_11739;
  reg        [7:0]    _zz_dataOut_payload_0_11740;
  reg        [7:0]    _zz_dataOut_payload_0_11741;
  reg        [7:0]    _zz_dataOut_payload_0_11742;
  reg        [7:0]    _zz_dataOut_payload_0_11743;
  reg        [7:0]    _zz_dataOut_payload_0_11744;
  reg        [7:0]    _zz_dataOut_payload_0_11745;
  reg        [7:0]    _zz_dataOut_payload_0_11746;
  reg        [7:0]    _zz_dataOut_payload_0_11747;
  reg        [7:0]    _zz_dataOut_payload_0_11748;
  reg        [7:0]    _zz_dataOut_payload_0_11749;
  reg        [7:0]    _zz_dataOut_payload_0_11750;
  reg        [7:0]    _zz_dataOut_payload_0_11751;
  reg        [7:0]    _zz_dataOut_payload_0_11752;
  reg        [7:0]    _zz_dataOut_payload_0_11753;
  reg        [7:0]    _zz_dataOut_payload_0_11754;
  reg        [7:0]    _zz_dataOut_payload_0_11755;
  reg        [7:0]    _zz_dataOut_payload_0_11756;
  reg        [7:0]    _zz_dataOut_payload_0_11757;
  reg        [7:0]    _zz_dataOut_payload_0_11758;
  reg        [7:0]    _zz_dataOut_payload_0_11759;
  reg        [7:0]    _zz_dataOut_payload_0_11760;
  reg        [7:0]    _zz_dataOut_payload_0_11761;
  reg        [7:0]    _zz_dataOut_payload_0_11762;
  reg        [7:0]    _zz_dataOut_payload_0_11763;
  reg        [7:0]    _zz_dataOut_payload_0_11764;
  reg        [7:0]    _zz_dataOut_payload_0_11765;
  reg        [7:0]    _zz_dataOut_payload_0_11766;
  reg        [7:0]    _zz_dataOut_payload_0_11767;
  reg        [7:0]    _zz_dataOut_payload_0_11768;
  reg        [7:0]    _zz_dataOut_payload_0_11769;
  reg        [7:0]    _zz_dataOut_payload_0_11770;
  reg        [7:0]    _zz_dataOut_payload_0_11771;
  reg        [7:0]    _zz_dataOut_payload_0_11772;
  reg        [7:0]    _zz_dataOut_payload_0_11773;
  reg        [7:0]    _zz_dataOut_payload_0_11774;
  reg        [7:0]    _zz_dataOut_payload_0_11775;
  reg        [7:0]    _zz_dataOut_payload_0_11776;
  reg        [7:0]    _zz_dataOut_payload_0_11777;
  reg        [7:0]    _zz_dataOut_payload_0_11778;
  reg        [7:0]    _zz_dataOut_payload_0_11779;
  reg        [7:0]    _zz_dataOut_payload_0_11780;
  reg        [7:0]    _zz_dataOut_payload_0_11781;
  reg        [7:0]    _zz_dataOut_payload_0_11782;
  reg        [7:0]    _zz_dataOut_payload_0_11783;
  reg        [7:0]    _zz_dataOut_payload_0_11784;
  reg        [7:0]    _zz_dataOut_payload_0_11785;
  reg        [7:0]    _zz_dataOut_payload_0_11786;
  reg        [7:0]    _zz_dataOut_payload_0_11787;
  reg        [7:0]    _zz_dataOut_payload_0_11788;
  reg        [7:0]    _zz_dataOut_payload_0_11789;
  reg        [7:0]    _zz_dataOut_payload_0_11790;
  reg        [7:0]    _zz_dataOut_payload_0_11791;
  reg        [7:0]    _zz_dataOut_payload_0_11792;
  reg        [7:0]    _zz_dataOut_payload_0_11793;
  reg        [7:0]    _zz_dataOut_payload_0_11794;
  reg        [7:0]    _zz_dataOut_payload_0_11795;
  reg        [7:0]    _zz_dataOut_payload_0_11796;
  reg        [7:0]    _zz_dataOut_payload_0_11797;
  reg        [7:0]    _zz_dataOut_payload_0_11798;
  reg        [7:0]    _zz_dataOut_payload_0_11799;
  reg        [7:0]    _zz_dataOut_payload_0_11800;
  reg        [7:0]    _zz_dataOut_payload_0_11801;
  reg        [7:0]    _zz_dataOut_payload_0_11802;
  reg        [7:0]    _zz_dataOut_payload_0_11803;
  reg        [7:0]    _zz_dataOut_payload_0_11804;
  reg        [7:0]    _zz_dataOut_payload_0_11805;
  reg        [7:0]    _zz_dataOut_payload_0_11806;
  reg        [7:0]    _zz_dataOut_payload_0_11807;
  reg        [7:0]    _zz_dataOut_payload_0_11808;
  reg        [7:0]    _zz_dataOut_payload_0_11809;
  reg        [7:0]    _zz_dataOut_payload_0_11810;
  reg        [7:0]    _zz_dataOut_payload_0_11811;
  reg        [7:0]    _zz_dataOut_payload_0_11812;
  reg        [7:0]    _zz_dataOut_payload_0_11813;
  reg        [7:0]    _zz_dataOut_payload_0_11814;
  reg        [7:0]    _zz_dataOut_payload_0_11815;
  reg        [7:0]    _zz_dataOut_payload_0_11816;
  reg        [7:0]    _zz_dataOut_payload_0_11817;
  reg        [7:0]    _zz_dataOut_payload_0_11818;
  reg        [7:0]    _zz_dataOut_payload_0_11819;
  reg        [7:0]    _zz_dataOut_payload_0_11820;
  reg        [7:0]    _zz_dataOut_payload_0_11821;
  reg        [7:0]    _zz_dataOut_payload_0_11822;
  reg        [7:0]    _zz_dataOut_payload_0_11823;
  reg        [7:0]    _zz_dataOut_payload_0_11824;
  reg        [7:0]    _zz_dataOut_payload_0_11825;
  reg        [7:0]    _zz_dataOut_payload_0_11826;
  reg        [7:0]    _zz_dataOut_payload_0_11827;
  reg        [7:0]    _zz_dataOut_payload_0_11828;
  reg        [7:0]    _zz_dataOut_payload_0_11829;
  reg        [7:0]    _zz_dataOut_payload_0_11830;
  reg        [7:0]    _zz_dataOut_payload_0_11831;
  reg        [7:0]    _zz_dataOut_payload_0_11832;
  reg        [7:0]    _zz_dataOut_payload_0_11833;
  reg        [7:0]    _zz_dataOut_payload_0_11834;
  reg        [7:0]    _zz_dataOut_payload_0_11835;
  reg        [7:0]    _zz_dataOut_payload_0_11836;
  reg        [7:0]    _zz_dataOut_payload_0_11837;
  reg        [7:0]    _zz_dataOut_payload_0_11838;
  reg        [7:0]    _zz_dataOut_payload_0_11839;
  reg        [7:0]    _zz_dataOut_payload_0_11840;
  reg        [7:0]    _zz_dataOut_payload_0_11841;
  reg        [7:0]    _zz_dataOut_payload_0_11842;
  reg        [7:0]    _zz_dataOut_payload_0_11843;
  reg        [7:0]    _zz_dataOut_payload_0_11844;
  reg        [7:0]    _zz_dataOut_payload_0_11845;
  reg        [7:0]    _zz_dataOut_payload_0_11846;
  reg        [7:0]    _zz_dataOut_payload_0_11847;
  reg        [7:0]    _zz_dataOut_payload_0_11848;
  reg        [7:0]    _zz_dataOut_payload_0_11849;
  reg        [7:0]    _zz_dataOut_payload_0_11850;
  reg        [7:0]    _zz_dataOut_payload_0_11851;
  reg        [7:0]    _zz_dataOut_payload_0_11852;
  reg        [7:0]    _zz_dataOut_payload_0_11853;
  reg        [7:0]    _zz_dataOut_payload_0_11854;
  reg        [7:0]    _zz_dataOut_payload_0_11855;
  reg        [7:0]    _zz_dataOut_payload_0_11856;
  reg        [7:0]    _zz_dataOut_payload_0_11857;
  reg        [7:0]    _zz_dataOut_payload_0_11858;
  reg        [7:0]    _zz_dataOut_payload_0_11859;
  reg        [7:0]    _zz_dataOut_payload_0_11860;
  reg        [7:0]    _zz_dataOut_payload_0_11861;
  reg        [7:0]    _zz_dataOut_payload_0_11862;
  reg        [7:0]    _zz_dataOut_payload_0_11863;
  reg        [7:0]    _zz_dataOut_payload_0_11864;
  reg        [7:0]    _zz_dataOut_payload_0_11865;
  reg        [7:0]    _zz_dataOut_payload_0_11866;
  reg        [7:0]    _zz_dataOut_payload_0_11867;
  reg        [7:0]    _zz_dataOut_payload_0_11868;
  reg        [7:0]    _zz_dataOut_payload_0_11869;
  reg        [7:0]    _zz_dataOut_payload_0_11870;
  reg        [7:0]    _zz_dataOut_payload_0_11871;
  reg        [7:0]    _zz_dataOut_payload_0_11872;
  reg        [7:0]    _zz_dataOut_payload_0_11873;
  reg        [7:0]    _zz_dataOut_payload_0_11874;
  reg        [7:0]    _zz_dataOut_payload_0_11875;
  reg        [7:0]    _zz_dataOut_payload_0_11876;
  reg        [7:0]    _zz_dataOut_payload_0_11877;
  reg        [7:0]    _zz_dataOut_payload_0_11878;
  reg        [7:0]    _zz_dataOut_payload_0_11879;
  reg        [7:0]    _zz_dataOut_payload_0_11880;
  reg        [7:0]    _zz_dataOut_payload_0_11881;
  reg        [7:0]    _zz_dataOut_payload_0_11882;
  reg        [7:0]    _zz_dataOut_payload_0_11883;
  reg        [7:0]    _zz_dataOut_payload_0_11884;
  reg        [7:0]    _zz_dataOut_payload_0_11885;
  reg        [7:0]    _zz_dataOut_payload_0_11886;
  reg        [7:0]    _zz_dataOut_payload_0_11887;
  reg        [7:0]    _zz_dataOut_payload_0_11888;
  reg        [7:0]    _zz_dataOut_payload_0_11889;
  reg        [7:0]    _zz_dataOut_payload_0_11890;
  reg        [7:0]    _zz_dataOut_payload_0_11891;
  reg        [7:0]    _zz_dataOut_payload_0_11892;
  reg        [7:0]    _zz_dataOut_payload_0_11893;
  reg        [7:0]    _zz_dataOut_payload_0_11894;
  reg        [7:0]    _zz_dataOut_payload_0_11895;
  reg        [7:0]    _zz_dataOut_payload_0_11896;
  reg        [7:0]    _zz_dataOut_payload_0_11897;
  reg        [7:0]    _zz_dataOut_payload_0_11898;
  reg        [7:0]    _zz_dataOut_payload_0_11899;
  reg        [7:0]    _zz_dataOut_payload_0_11900;
  reg        [7:0]    _zz_dataOut_payload_0_11901;
  reg        [7:0]    _zz_dataOut_payload_0_11902;
  reg        [7:0]    _zz_dataOut_payload_0_11903;
  wire                _zz_dataOut_payload_0_11904;
  wire       [7:0]    _zz_dataOut_payload_0_11905;
  wire       [7:0]    _zz_dataOut_payload_0_11906;
  wire                _zz_dataOut_payload_0_11907;
  wire       [7:0]    _zz_dataOut_payload_0_11908;
  wire       [7:0]    _zz_dataOut_payload_0_11909;
  wire                _zz_dataOut_payload_0_11910;
  wire       [7:0]    _zz_dataOut_payload_0_11911;
  wire       [7:0]    _zz_dataOut_payload_0_11912;
  wire                _zz_dataOut_payload_0_11913;
  wire       [7:0]    _zz_dataOut_payload_0_11914;
  wire       [7:0]    _zz_dataOut_payload_0_11915;
  wire                _zz_dataOut_payload_0_11916;
  wire       [7:0]    _zz_dataOut_payload_0_11917;
  wire       [7:0]    _zz_dataOut_payload_0_11918;
  wire                _zz_dataOut_payload_0_11919;
  wire       [7:0]    _zz_dataOut_payload_0_11920;
  wire       [7:0]    _zz_dataOut_payload_0_11921;
  wire                _zz_dataOut_payload_0_11922;
  wire       [7:0]    _zz_dataOut_payload_0_11923;
  wire       [7:0]    _zz_dataOut_payload_0_11924;
  wire                _zz_dataOut_payload_0_11925;
  wire       [7:0]    _zz_dataOut_payload_0_11926;
  wire       [7:0]    _zz_dataOut_payload_0_11927;
  wire                _zz_dataOut_payload_0_11928;
  wire       [7:0]    _zz_dataOut_payload_0_11929;
  wire       [7:0]    _zz_dataOut_payload_0_11930;
  wire                _zz_dataOut_payload_0_11931;
  wire       [7:0]    _zz_dataOut_payload_0_11932;
  wire       [7:0]    _zz_dataOut_payload_0_11933;
  wire                _zz_dataOut_payload_0_11934;
  wire       [7:0]    _zz_dataOut_payload_0_11935;
  wire       [7:0]    _zz_dataOut_payload_0_11936;
  wire                _zz_dataOut_payload_0_11937;
  wire       [7:0]    _zz_dataOut_payload_0_11938;
  wire       [7:0]    _zz_dataOut_payload_0_11939;
  wire                _zz_dataOut_payload_0_11940;
  wire       [7:0]    _zz_dataOut_payload_0_11941;
  wire       [7:0]    _zz_dataOut_payload_0_11942;
  wire                _zz_dataOut_payload_0_11943;
  wire       [7:0]    _zz_dataOut_payload_0_11944;
  wire       [7:0]    _zz_dataOut_payload_0_11945;
  wire                _zz_dataOut_payload_0_11946;
  wire       [7:0]    _zz_dataOut_payload_0_11947;
  wire       [7:0]    _zz_dataOut_payload_0_11948;
  wire                _zz_dataOut_payload_0_11949;
  wire       [7:0]    _zz_dataOut_payload_0_11950;
  wire       [7:0]    _zz_dataOut_payload_0_11951;
  wire                _zz_dataOut_payload_0_11952;
  wire       [7:0]    _zz_dataOut_payload_0_11953;
  wire       [7:0]    _zz_dataOut_payload_0_11954;
  wire                _zz_dataOut_payload_0_11955;
  wire       [7:0]    _zz_dataOut_payload_0_11956;
  wire       [7:0]    _zz_dataOut_payload_0_11957;
  wire                _zz_dataOut_payload_0_11958;
  wire       [7:0]    _zz_dataOut_payload_0_11959;
  wire       [7:0]    _zz_dataOut_payload_0_11960;
  wire                _zz_dataOut_payload_0_11961;
  wire       [7:0]    _zz_dataOut_payload_0_11962;
  wire       [7:0]    _zz_dataOut_payload_0_11963;
  wire                _zz_dataOut_payload_0_11964;
  wire       [7:0]    _zz_dataOut_payload_0_11965;
  wire       [7:0]    _zz_dataOut_payload_0_11966;
  wire                _zz_dataOut_payload_0_11967;
  wire       [7:0]    _zz_dataOut_payload_0_11968;
  wire       [7:0]    _zz_dataOut_payload_0_11969;
  wire                _zz_dataOut_payload_0_11970;
  wire       [7:0]    _zz_dataOut_payload_0_11971;
  wire       [7:0]    _zz_dataOut_payload_0_11972;
  wire                _zz_dataOut_payload_0_11973;
  wire       [7:0]    _zz_dataOut_payload_0_11974;
  wire       [7:0]    _zz_dataOut_payload_0_11975;
  wire                _zz_dataOut_payload_0_11976;
  wire       [7:0]    _zz_dataOut_payload_0_11977;
  wire       [7:0]    _zz_dataOut_payload_0_11978;
  wire                _zz_dataOut_payload_0_11979;
  wire       [7:0]    _zz_dataOut_payload_0_11980;
  wire       [7:0]    _zz_dataOut_payload_0_11981;
  wire                _zz_dataOut_payload_0_11982;
  wire       [7:0]    _zz_dataOut_payload_0_11983;
  wire       [7:0]    _zz_dataOut_payload_0_11984;
  wire                _zz_dataOut_payload_0_11985;
  wire       [7:0]    _zz_dataOut_payload_0_11986;
  wire       [7:0]    _zz_dataOut_payload_0_11987;
  wire                _zz_dataOut_payload_0_11988;
  wire       [7:0]    _zz_dataOut_payload_0_11989;
  wire       [7:0]    _zz_dataOut_payload_0_11990;
  wire                _zz_dataOut_payload_0_11991;
  wire       [7:0]    _zz_dataOut_payload_0_11992;
  wire       [7:0]    _zz_dataOut_payload_0_11993;
  wire                _zz_dataOut_payload_0_11994;
  wire       [7:0]    _zz_dataOut_payload_0_11995;
  wire       [7:0]    _zz_dataOut_payload_0_11996;
  wire                _zz_dataOut_payload_0_11997;
  wire       [7:0]    _zz_dataOut_payload_0_11998;
  wire       [7:0]    _zz_dataOut_payload_0_11999;
  wire                _zz_dataOut_payload_0_12000;
  wire       [7:0]    _zz_dataOut_payload_0_12001;
  wire       [7:0]    _zz_dataOut_payload_0_12002;
  wire                _zz_dataOut_payload_0_12003;
  wire       [7:0]    _zz_dataOut_payload_0_12004;
  wire       [7:0]    _zz_dataOut_payload_0_12005;
  wire                _zz_dataOut_payload_0_12006;
  wire       [7:0]    _zz_dataOut_payload_0_12007;
  wire       [7:0]    _zz_dataOut_payload_0_12008;
  wire                _zz_dataOut_payload_0_12009;
  wire       [7:0]    _zz_dataOut_payload_0_12010;
  wire       [7:0]    _zz_dataOut_payload_0_12011;
  wire                _zz_dataOut_payload_0_12012;
  wire       [7:0]    _zz_dataOut_payload_0_12013;
  wire       [7:0]    _zz_dataOut_payload_0_12014;
  wire                _zz_dataOut_payload_0_12015;
  wire       [7:0]    _zz_dataOut_payload_0_12016;
  wire       [7:0]    _zz_dataOut_payload_0_12017;
  wire                _zz_dataOut_payload_0_12018;
  wire       [7:0]    _zz_dataOut_payload_0_12019;
  wire       [7:0]    _zz_dataOut_payload_0_12020;
  wire                _zz_dataOut_payload_0_12021;
  wire       [7:0]    _zz_dataOut_payload_0_12022;
  wire       [7:0]    _zz_dataOut_payload_0_12023;
  wire                _zz_dataOut_payload_0_12024;
  wire       [7:0]    _zz_dataOut_payload_0_12025;
  wire       [7:0]    _zz_dataOut_payload_0_12026;
  wire                _zz_dataOut_payload_0_12027;
  wire       [7:0]    _zz_dataOut_payload_0_12028;
  wire       [7:0]    _zz_dataOut_payload_0_12029;
  wire                _zz_dataOut_payload_0_12030;
  wire       [7:0]    _zz_dataOut_payload_0_12031;
  wire       [7:0]    _zz_dataOut_payload_0_12032;
  wire                _zz_dataOut_payload_0_12033;
  wire       [7:0]    _zz_dataOut_payload_0_12034;
  wire       [7:0]    _zz_dataOut_payload_0_12035;
  wire                _zz_dataOut_payload_0_12036;
  wire       [7:0]    _zz_dataOut_payload_0_12037;
  wire       [7:0]    _zz_dataOut_payload_0_12038;
  wire                _zz_dataOut_payload_0_12039;
  wire       [7:0]    _zz_dataOut_payload_0_12040;
  wire       [7:0]    _zz_dataOut_payload_0_12041;
  wire                _zz_dataOut_payload_0_12042;
  wire       [7:0]    _zz_dataOut_payload_0_12043;
  wire       [7:0]    _zz_dataOut_payload_0_12044;
  wire                _zz_dataOut_payload_0_12045;
  wire       [7:0]    _zz_dataOut_payload_0_12046;
  wire       [7:0]    _zz_dataOut_payload_0_12047;
  wire                _zz_dataOut_payload_0_12048;
  wire       [7:0]    _zz_dataOut_payload_0_12049;
  wire       [7:0]    _zz_dataOut_payload_0_12050;
  wire                _zz_dataOut_payload_0_12051;
  wire       [7:0]    _zz_dataOut_payload_0_12052;
  wire       [7:0]    _zz_dataOut_payload_0_12053;
  wire                _zz_dataOut_payload_0_12054;
  wire       [7:0]    _zz_dataOut_payload_0_12055;
  wire       [7:0]    _zz_dataOut_payload_0_12056;
  wire                _zz_dataOut_payload_0_12057;
  wire       [7:0]    _zz_dataOut_payload_0_12058;
  wire       [7:0]    _zz_dataOut_payload_0_12059;
  wire                _zz_dataOut_payload_0_12060;
  wire       [7:0]    _zz_dataOut_payload_0_12061;
  wire       [7:0]    _zz_dataOut_payload_0_12062;
  wire                _zz_dataOut_payload_0_12063;
  wire       [7:0]    _zz_dataOut_payload_0_12064;
  wire       [7:0]    _zz_dataOut_payload_0_12065;
  wire                _zz_dataOut_payload_0_12066;
  wire       [7:0]    _zz_dataOut_payload_0_12067;
  wire       [7:0]    _zz_dataOut_payload_0_12068;
  wire                _zz_dataOut_payload_0_12069;
  wire       [7:0]    _zz_dataOut_payload_0_12070;
  wire       [7:0]    _zz_dataOut_payload_0_12071;
  wire                _zz_dataOut_payload_0_12072;
  wire       [7:0]    _zz_dataOut_payload_0_12073;
  wire       [7:0]    _zz_dataOut_payload_0_12074;
  wire                _zz_dataOut_payload_0_12075;
  wire       [7:0]    _zz_dataOut_payload_0_12076;
  wire       [7:0]    _zz_dataOut_payload_0_12077;
  wire                _zz_dataOut_payload_0_12078;
  wire       [7:0]    _zz_dataOut_payload_0_12079;
  wire       [7:0]    _zz_dataOut_payload_0_12080;
  wire                _zz_dataOut_payload_0_12081;
  wire       [7:0]    _zz_dataOut_payload_0_12082;
  wire       [7:0]    _zz_dataOut_payload_0_12083;
  wire                _zz_dataOut_payload_0_12084;
  wire       [7:0]    _zz_dataOut_payload_0_12085;
  wire       [7:0]    _zz_dataOut_payload_0_12086;
  wire                _zz_dataOut_payload_0_12087;
  wire       [7:0]    _zz_dataOut_payload_0_12088;
  wire       [7:0]    _zz_dataOut_payload_0_12089;
  wire                _zz_dataOut_payload_0_12090;
  wire       [7:0]    _zz_dataOut_payload_0_12091;
  wire       [7:0]    _zz_dataOut_payload_0_12092;
  wire                _zz_dataOut_payload_0_12093;
  wire       [7:0]    _zz_dataOut_payload_0_12094;
  wire       [7:0]    _zz_dataOut_payload_0_12095;
  wire                _zz_dataOut_payload_0_12096;
  wire       [7:0]    _zz_dataOut_payload_0_12097;
  wire       [7:0]    _zz_dataOut_payload_0_12098;
  wire                _zz_dataOut_payload_0_12099;
  wire       [7:0]    _zz_dataOut_payload_0_12100;
  wire       [7:0]    _zz_dataOut_payload_0_12101;
  wire                _zz_dataOut_payload_0_12102;
  wire       [7:0]    _zz_dataOut_payload_0_12103;
  wire       [7:0]    _zz_dataOut_payload_0_12104;
  wire                _zz_dataOut_payload_0_12105;
  wire       [7:0]    _zz_dataOut_payload_0_12106;
  wire       [7:0]    _zz_dataOut_payload_0_12107;
  wire                _zz_dataOut_payload_0_12108;
  wire       [7:0]    _zz_dataOut_payload_0_12109;
  wire       [7:0]    _zz_dataOut_payload_0_12110;
  wire                _zz_dataOut_payload_0_12111;
  wire       [7:0]    _zz_dataOut_payload_0_12112;
  wire       [7:0]    _zz_dataOut_payload_0_12113;
  wire                _zz_dataOut_payload_0_12114;
  wire       [7:0]    _zz_dataOut_payload_0_12115;
  wire       [7:0]    _zz_dataOut_payload_0_12116;
  wire                _zz_dataOut_payload_0_12117;
  wire       [7:0]    _zz_dataOut_payload_0_12118;
  wire       [7:0]    _zz_dataOut_payload_0_12119;
  wire                _zz_dataOut_payload_0_12120;
  wire       [7:0]    _zz_dataOut_payload_0_12121;
  wire       [7:0]    _zz_dataOut_payload_0_12122;
  wire                _zz_dataOut_payload_0_12123;
  wire       [7:0]    _zz_dataOut_payload_0_12124;
  wire       [7:0]    _zz_dataOut_payload_0_12125;
  wire                _zz_dataOut_payload_0_12126;
  wire       [7:0]    _zz_dataOut_payload_0_12127;
  wire       [7:0]    _zz_dataOut_payload_0_12128;
  wire                _zz_dataOut_payload_0_12129;
  wire       [7:0]    _zz_dataOut_payload_0_12130;
  wire       [7:0]    _zz_dataOut_payload_0_12131;
  wire                _zz_dataOut_payload_0_12132;
  wire       [7:0]    _zz_dataOut_payload_0_12133;
  wire       [7:0]    _zz_dataOut_payload_0_12134;
  wire                _zz_dataOut_payload_0_12135;
  wire       [7:0]    _zz_dataOut_payload_0_12136;
  wire       [7:0]    _zz_dataOut_payload_0_12137;
  wire                _zz_dataOut_payload_0_12138;
  wire       [7:0]    _zz_dataOut_payload_0_12139;
  wire       [7:0]    _zz_dataOut_payload_0_12140;
  wire                _zz_dataOut_payload_0_12141;
  wire       [7:0]    _zz_dataOut_payload_0_12142;
  wire       [7:0]    _zz_dataOut_payload_0_12143;
  wire                _zz_dataOut_payload_0_12144;
  wire       [7:0]    _zz_dataOut_payload_0_12145;
  wire       [7:0]    _zz_dataOut_payload_0_12146;
  wire                _zz_dataOut_payload_0_12147;
  wire       [7:0]    _zz_dataOut_payload_0_12148;
  wire       [7:0]    _zz_dataOut_payload_0_12149;
  wire                _zz_dataOut_payload_0_12150;
  wire       [7:0]    _zz_dataOut_payload_0_12151;
  wire       [7:0]    _zz_dataOut_payload_0_12152;
  wire                _zz_dataOut_payload_0_12153;
  wire       [7:0]    _zz_dataOut_payload_0_12154;
  wire       [7:0]    _zz_dataOut_payload_0_12155;
  wire                _zz_dataOut_payload_0_12156;
  wire       [7:0]    _zz_dataOut_payload_0_12157;
  wire       [7:0]    _zz_dataOut_payload_0_12158;
  wire                _zz_dataOut_payload_0_12159;
  wire       [7:0]    _zz_dataOut_payload_0_12160;
  wire       [7:0]    _zz_dataOut_payload_0_12161;
  wire                _zz_dataOut_payload_0_12162;
  wire       [7:0]    _zz_dataOut_payload_0_12163;
  wire       [7:0]    _zz_dataOut_payload_0_12164;
  wire                _zz_dataOut_payload_0_12165;
  wire       [7:0]    _zz_dataOut_payload_0_12166;
  wire       [7:0]    _zz_dataOut_payload_0_12167;
  wire                _zz_dataOut_payload_0_12168;
  wire       [7:0]    _zz_dataOut_payload_0_12169;
  wire       [7:0]    _zz_dataOut_payload_0_12170;
  wire                _zz_dataOut_payload_0_12171;
  wire       [7:0]    _zz_dataOut_payload_0_12172;
  wire       [7:0]    _zz_dataOut_payload_0_12173;
  wire                _zz_dataOut_payload_0_12174;
  wire       [7:0]    _zz_dataOut_payload_0_12175;
  wire       [7:0]    _zz_dataOut_payload_0_12176;
  wire                _zz_dataOut_payload_0_12177;
  wire       [7:0]    _zz_dataOut_payload_0_12178;
  wire       [7:0]    _zz_dataOut_payload_0_12179;
  wire                _zz_dataOut_payload_0_12180;
  wire       [7:0]    _zz_dataOut_payload_0_12181;
  wire       [7:0]    _zz_dataOut_payload_0_12182;
  wire                _zz_dataOut_payload_0_12183;
  wire       [7:0]    _zz_dataOut_payload_0_12184;
  wire       [7:0]    _zz_dataOut_payload_0_12185;
  wire                _zz_dataOut_payload_0_12186;
  wire       [7:0]    _zz_dataOut_payload_0_12187;
  wire       [7:0]    _zz_dataOut_payload_0_12188;
  wire                _zz_dataOut_payload_0_12189;
  wire       [7:0]    _zz_dataOut_payload_0_12190;
  wire       [7:0]    _zz_dataOut_payload_0_12191;
  wire                _zz_dataOut_payload_0_12192;
  wire       [7:0]    _zz_dataOut_payload_0_12193;
  wire       [7:0]    _zz_dataOut_payload_0_12194;
  wire                _zz_dataOut_payload_0_12195;
  wire       [7:0]    _zz_dataOut_payload_0_12196;
  wire       [7:0]    _zz_dataOut_payload_0_12197;
  wire                _zz_dataOut_payload_0_12198;
  wire       [7:0]    _zz_dataOut_payload_0_12199;
  wire       [7:0]    _zz_dataOut_payload_0_12200;
  wire                _zz_dataOut_payload_0_12201;
  wire       [7:0]    _zz_dataOut_payload_0_12202;
  wire       [7:0]    _zz_dataOut_payload_0_12203;
  wire                _zz_dataOut_payload_0_12204;
  wire       [7:0]    _zz_dataOut_payload_0_12205;
  wire       [7:0]    _zz_dataOut_payload_0_12206;
  wire                _zz_dataOut_payload_0_12207;
  wire       [7:0]    _zz_dataOut_payload_0_12208;
  wire       [7:0]    _zz_dataOut_payload_0_12209;
  wire                _zz_dataOut_payload_0_12210;
  wire       [7:0]    _zz_dataOut_payload_0_12211;
  wire       [7:0]    _zz_dataOut_payload_0_12212;
  wire                _zz_dataOut_payload_0_12213;
  wire       [7:0]    _zz_dataOut_payload_0_12214;
  wire       [7:0]    _zz_dataOut_payload_0_12215;
  wire                _zz_dataOut_payload_0_12216;
  wire       [7:0]    _zz_dataOut_payload_0_12217;
  wire       [7:0]    _zz_dataOut_payload_0_12218;
  wire                _zz_dataOut_payload_0_12219;
  wire       [7:0]    _zz_dataOut_payload_0_12220;
  wire       [7:0]    _zz_dataOut_payload_0_12221;
  wire                _zz_dataOut_payload_0_12222;
  wire       [7:0]    _zz_dataOut_payload_0_12223;
  wire       [7:0]    _zz_dataOut_payload_0_12224;
  wire                _zz_dataOut_payload_0_12225;
  wire       [7:0]    _zz_dataOut_payload_0_12226;
  wire       [7:0]    _zz_dataOut_payload_0_12227;
  wire                _zz_dataOut_payload_0_12228;
  wire       [7:0]    _zz_dataOut_payload_0_12229;
  wire       [7:0]    _zz_dataOut_payload_0_12230;
  wire                _zz_dataOut_payload_0_12231;
  wire       [7:0]    _zz_dataOut_payload_0_12232;
  wire       [7:0]    _zz_dataOut_payload_0_12233;
  wire                _zz_dataOut_payload_0_12234;
  wire       [7:0]    _zz_dataOut_payload_0_12235;
  wire       [7:0]    _zz_dataOut_payload_0_12236;
  wire                _zz_dataOut_payload_0_12237;
  wire       [7:0]    _zz_dataOut_payload_0_12238;
  wire       [7:0]    _zz_dataOut_payload_0_12239;
  wire                _zz_dataOut_payload_0_12240;
  wire       [7:0]    _zz_dataOut_payload_0_12241;
  wire       [7:0]    _zz_dataOut_payload_0_12242;
  wire                _zz_dataOut_payload_0_12243;
  wire       [7:0]    _zz_dataOut_payload_0_12244;
  wire       [7:0]    _zz_dataOut_payload_0_12245;
  wire                _zz_dataOut_payload_0_12246;
  wire       [7:0]    _zz_dataOut_payload_0_12247;
  wire       [7:0]    _zz_dataOut_payload_0_12248;
  wire                _zz_dataOut_payload_0_12249;
  wire       [7:0]    _zz_dataOut_payload_0_12250;
  wire       [7:0]    _zz_dataOut_payload_0_12251;
  wire                _zz_dataOut_payload_0_12252;
  wire       [7:0]    _zz_dataOut_payload_0_12253;
  wire       [7:0]    _zz_dataOut_payload_0_12254;
  wire                _zz_dataOut_payload_0_12255;
  wire       [7:0]    _zz_dataOut_payload_0_12256;
  wire       [7:0]    _zz_dataOut_payload_0_12257;
  wire                _zz_dataOut_payload_0_12258;
  wire       [7:0]    _zz_dataOut_payload_0_12259;
  wire       [7:0]    _zz_dataOut_payload_0_12260;
  wire                _zz_dataOut_payload_0_12261;
  wire       [7:0]    _zz_dataOut_payload_0_12262;
  wire       [7:0]    _zz_dataOut_payload_0_12263;
  wire                _zz_dataOut_payload_0_12264;
  wire       [7:0]    _zz_dataOut_payload_0_12265;
  wire       [7:0]    _zz_dataOut_payload_0_12266;
  wire                _zz_dataOut_payload_0_12267;
  wire       [7:0]    _zz_dataOut_payload_0_12268;
  wire       [7:0]    _zz_dataOut_payload_0_12269;
  wire                _zz_dataOut_payload_0_12270;
  wire       [7:0]    _zz_dataOut_payload_0_12271;
  wire       [7:0]    _zz_dataOut_payload_0_12272;
  wire                _zz_dataOut_payload_0_12273;
  wire       [7:0]    _zz_dataOut_payload_0_12274;
  wire       [7:0]    _zz_dataOut_payload_0_12275;
  wire                _zz_dataOut_payload_0_12276;
  wire       [7:0]    _zz_dataOut_payload_0_12277;
  wire       [7:0]    _zz_dataOut_payload_0_12278;
  wire                _zz_dataOut_payload_0_12279;
  wire       [7:0]    _zz_dataOut_payload_0_12280;
  wire       [7:0]    _zz_dataOut_payload_0_12281;
  wire                _zz_dataOut_payload_0_12282;
  wire                _zz_dataOut_payload_0_12283;
  reg        [7:0]    _zz_dataOut_payload_0_12284;
  reg        [7:0]    _zz_dataOut_payload_0_12285;
  reg        [7:0]    _zz_dataOut_payload_0_12286;
  reg        [7:0]    _zz_dataOut_payload_0_12287;
  wire                _zz_dataOut_payload_0_12288;
  wire       [7:0]    _zz_dataOut_payload_0_12289;
  wire       [7:0]    _zz_dataOut_payload_0_12290;
  wire                _zz_dataOut_payload_0_12291;
  wire       [7:0]    _zz_dataOut_payload_0_12292;
  wire       [7:0]    _zz_dataOut_payload_0_12293;
  wire                _zz_dataOut_payload_0_12294;
  wire                _zz_dataOut_payload_0_12295;
  reg        [7:0]    _zz_dataOut_payload_0_12296;
  reg        [7:0]    _zz_dataOut_payload_0_12297;
  reg        [7:0]    _zz_dataOut_payload_0_12298;
  reg        [7:0]    _zz_dataOut_payload_0_12299;
  reg        [7:0]    _zz_dataOut_payload_0_12300;
  reg        [7:0]    _zz_dataOut_payload_0_12301;
  reg        [7:0]    _zz_dataOut_payload_0_12302;
  reg        [7:0]    _zz_dataOut_payload_0_12303;
  reg        [7:0]    _zz_dataOut_payload_0_12304;
  reg        [7:0]    _zz_dataOut_payload_0_12305;
  reg        [7:0]    _zz_dataOut_payload_0_12306;
  reg        [7:0]    _zz_dataOut_payload_0_12307;
  wire                _zz_dataOut_payload_0_12308;
  wire       [7:0]    _zz_dataOut_payload_0_12309;
  wire       [7:0]    _zz_dataOut_payload_0_12310;
  wire                _zz_dataOut_payload_0_12311;
  wire       [7:0]    _zz_dataOut_payload_0_12312;
  wire       [7:0]    _zz_dataOut_payload_0_12313;
  wire                _zz_dataOut_payload_0_12314;
  wire       [7:0]    _zz_dataOut_payload_0_12315;
  wire       [7:0]    _zz_dataOut_payload_0_12316;
  wire                _zz_dataOut_payload_0_12317;
  wire       [7:0]    _zz_dataOut_payload_0_12318;
  wire       [7:0]    _zz_dataOut_payload_0_12319;
  wire                _zz_dataOut_payload_0_12320;
  wire       [7:0]    _zz_dataOut_payload_0_12321;
  wire       [7:0]    _zz_dataOut_payload_0_12322;
  wire                _zz_dataOut_payload_0_12323;
  wire       [7:0]    _zz_dataOut_payload_0_12324;
  wire       [7:0]    _zz_dataOut_payload_0_12325;
  wire                _zz_dataOut_payload_0_12326;
  wire                _zz_dataOut_payload_0_12327;
  reg        [7:0]    _zz_dataOut_payload_0_12328;
  reg        [7:0]    _zz_dataOut_payload_0_12329;
  reg        [7:0]    _zz_dataOut_payload_0_12330;
  reg        [7:0]    _zz_dataOut_payload_0_12331;
  wire                _zz_dataOut_payload_0_12332;
  wire       [7:0]    _zz_dataOut_payload_0_12333;
  wire       [7:0]    _zz_dataOut_payload_0_12334;
  wire                _zz_dataOut_payload_0_12335;
  wire       [7:0]    _zz_dataOut_payload_0_12336;
  wire       [7:0]    _zz_dataOut_payload_0_12337;
  wire                _zz_dataOut_payload_0_12338;
  wire                _zz_dataOut_payload_0_12339;
  reg        [7:0]    _zz_dataOut_payload_0_12340;
  reg        [7:0]    _zz_dataOut_payload_0_12341;
  reg        [7:0]    _zz_dataOut_payload_0_12342;
  reg        [7:0]    _zz_dataOut_payload_0_12343;
  reg        [7:0]    _zz_dataOut_payload_0_12344;
  reg        [7:0]    _zz_dataOut_payload_0_12345;
  reg        [7:0]    _zz_dataOut_payload_0_12346;
  reg        [7:0]    _zz_dataOut_payload_0_12347;
  reg        [7:0]    _zz_dataOut_payload_0_12348;
  reg        [7:0]    _zz_dataOut_payload_0_12349;
  reg        [7:0]    _zz_dataOut_payload_0_12350;
  reg        [7:0]    _zz_dataOut_payload_0_12351;
  reg        [7:0]    _zz_dataOut_payload_0_12352;
  reg        [7:0]    _zz_dataOut_payload_0_12353;
  reg        [7:0]    _zz_dataOut_payload_0_12354;
  reg        [7:0]    _zz_dataOut_payload_0_12355;
  reg        [7:0]    _zz_dataOut_payload_0_12356;
  reg        [7:0]    _zz_dataOut_payload_0_12357;
  reg        [7:0]    _zz_dataOut_payload_0_12358;
  reg        [7:0]    _zz_dataOut_payload_0_12359;
  reg        [7:0]    _zz_dataOut_payload_0_12360;
  reg        [7:0]    _zz_dataOut_payload_0_12361;
  reg        [7:0]    _zz_dataOut_payload_0_12362;
  reg        [7:0]    _zz_dataOut_payload_0_12363;
  reg        [7:0]    _zz_dataOut_payload_0_12364;
  reg        [7:0]    _zz_dataOut_payload_0_12365;
  reg        [7:0]    _zz_dataOut_payload_0_12366;
  reg        [7:0]    _zz_dataOut_payload_0_12367;
  wire                _zz_dataOut_payload_0_12368;
  wire       [7:0]    _zz_dataOut_payload_0_12369;
  wire       [7:0]    _zz_dataOut_payload_0_12370;
  wire                _zz_dataOut_payload_0_12371;
  wire       [7:0]    _zz_dataOut_payload_0_12372;
  wire       [7:0]    _zz_dataOut_payload_0_12373;
  wire                _zz_dataOut_payload_0_12374;
  wire       [7:0]    _zz_dataOut_payload_0_12375;
  wire       [7:0]    _zz_dataOut_payload_0_12376;
  wire                _zz_dataOut_payload_0_12377;
  wire       [7:0]    _zz_dataOut_payload_0_12378;
  wire       [7:0]    _zz_dataOut_payload_0_12379;
  wire                _zz_dataOut_payload_0_12380;
  wire       [7:0]    _zz_dataOut_payload_0_12381;
  wire       [7:0]    _zz_dataOut_payload_0_12382;
  wire                _zz_dataOut_payload_0_12383;
  wire       [7:0]    _zz_dataOut_payload_0_12384;
  wire       [7:0]    _zz_dataOut_payload_0_12385;
  wire                _zz_dataOut_payload_0_12386;
  wire       [7:0]    _zz_dataOut_payload_0_12387;
  wire       [7:0]    _zz_dataOut_payload_0_12388;
  wire                _zz_dataOut_payload_0_12389;
  wire       [7:0]    _zz_dataOut_payload_0_12390;
  wire       [7:0]    _zz_dataOut_payload_0_12391;
  wire                _zz_dataOut_payload_0_12392;
  wire       [7:0]    _zz_dataOut_payload_0_12393;
  wire       [7:0]    _zz_dataOut_payload_0_12394;
  wire                _zz_dataOut_payload_0_12395;
  wire       [7:0]    _zz_dataOut_payload_0_12396;
  wire       [7:0]    _zz_dataOut_payload_0_12397;
  wire                _zz_dataOut_payload_0_12398;
  wire       [7:0]    _zz_dataOut_payload_0_12399;
  wire       [7:0]    _zz_dataOut_payload_0_12400;
  wire                _zz_dataOut_payload_0_12401;
  wire       [7:0]    _zz_dataOut_payload_0_12402;
  wire       [7:0]    _zz_dataOut_payload_0_12403;
  wire                _zz_dataOut_payload_0_12404;
  wire       [7:0]    _zz_dataOut_payload_0_12405;
  wire       [7:0]    _zz_dataOut_payload_0_12406;
  wire                _zz_dataOut_payload_0_12407;
  wire       [7:0]    _zz_dataOut_payload_0_12408;
  wire       [7:0]    _zz_dataOut_payload_0_12409;
  wire                _zz_dataOut_payload_0_12410;
  wire                _zz_dataOut_payload_0_12411;
  reg        [7:0]    _zz_dataOut_payload_0_12412;
  reg        [7:0]    _zz_dataOut_payload_0_12413;
  reg        [7:0]    _zz_dataOut_payload_0_12414;
  reg        [7:0]    _zz_dataOut_payload_0_12415;
  wire                _zz_dataOut_payload_0_12416;
  wire       [7:0]    _zz_dataOut_payload_0_12417;
  wire       [7:0]    _zz_dataOut_payload_0_12418;
  wire                _zz_dataOut_payload_0_12419;
  wire       [7:0]    _zz_dataOut_payload_0_12420;
  wire       [7:0]    _zz_dataOut_payload_0_12421;
  wire                _zz_dataOut_payload_0_12422;
  wire                _zz_dataOut_payload_0_12423;
  reg        [7:0]    _zz_dataOut_payload_0_12424;
  reg        [7:0]    _zz_dataOut_payload_0_12425;
  reg        [7:0]    _zz_dataOut_payload_0_12426;
  reg        [7:0]    _zz_dataOut_payload_0_12427;
  reg        [7:0]    _zz_dataOut_payload_0_12428;
  reg        [7:0]    _zz_dataOut_payload_0_12429;
  reg        [7:0]    _zz_dataOut_payload_0_12430;
  reg        [7:0]    _zz_dataOut_payload_0_12431;
  reg        [7:0]    _zz_dataOut_payload_0_12432;
  reg        [7:0]    _zz_dataOut_payload_0_12433;
  reg        [7:0]    _zz_dataOut_payload_0_12434;
  reg        [7:0]    _zz_dataOut_payload_0_12435;
  wire                _zz_dataOut_payload_0_12436;
  wire       [7:0]    _zz_dataOut_payload_0_12437;
  wire       [7:0]    _zz_dataOut_payload_0_12438;
  wire                _zz_dataOut_payload_0_12439;
  wire       [7:0]    _zz_dataOut_payload_0_12440;
  wire       [7:0]    _zz_dataOut_payload_0_12441;
  wire                _zz_dataOut_payload_0_12442;
  wire       [7:0]    _zz_dataOut_payload_0_12443;
  wire       [7:0]    _zz_dataOut_payload_0_12444;
  wire                _zz_dataOut_payload_0_12445;
  wire       [7:0]    _zz_dataOut_payload_0_12446;
  wire       [7:0]    _zz_dataOut_payload_0_12447;
  wire                _zz_dataOut_payload_0_12448;
  wire       [7:0]    _zz_dataOut_payload_0_12449;
  wire       [7:0]    _zz_dataOut_payload_0_12450;
  wire                _zz_dataOut_payload_0_12451;
  wire       [7:0]    _zz_dataOut_payload_0_12452;
  wire       [7:0]    _zz_dataOut_payload_0_12453;
  wire                _zz_dataOut_payload_0_12454;
  wire                _zz_dataOut_payload_0_12455;
  reg        [7:0]    _zz_dataOut_payload_0_12456;
  reg        [7:0]    _zz_dataOut_payload_0_12457;
  reg        [7:0]    _zz_dataOut_payload_0_12458;
  reg        [7:0]    _zz_dataOut_payload_0_12459;
  wire                _zz_dataOut_payload_0_12460;
  wire       [7:0]    _zz_dataOut_payload_0_12461;
  wire       [7:0]    _zz_dataOut_payload_0_12462;
  wire                _zz_dataOut_payload_0_12463;
  wire       [7:0]    _zz_dataOut_payload_0_12464;
  wire       [7:0]    _zz_dataOut_payload_0_12465;
  wire                _zz_dataOut_payload_0_12466;
  wire                _zz_dataOut_payload_0_12467;
  reg        [7:0]    _zz_dataOut_payload_0_12468;
  reg        [7:0]    _zz_dataOut_payload_0_12469;
  reg        [7:0]    _zz_dataOut_payload_0_12470;
  reg        [7:0]    _zz_dataOut_payload_0_12471;
  reg        [7:0]    _zz_dataOut_payload_0_12472;
  reg        [7:0]    _zz_dataOut_payload_0_12473;
  reg        [7:0]    _zz_dataOut_payload_0_12474;
  reg        [7:0]    _zz_dataOut_payload_0_12475;
  reg        [7:0]    _zz_dataOut_payload_0_12476;
  reg        [7:0]    _zz_dataOut_payload_0_12477;
  reg        [7:0]    _zz_dataOut_payload_0_12478;
  reg        [7:0]    _zz_dataOut_payload_0_12479;
  reg        [7:0]    _zz_dataOut_payload_0_12480;
  reg        [7:0]    _zz_dataOut_payload_0_12481;
  reg        [7:0]    _zz_dataOut_payload_0_12482;
  reg        [7:0]    _zz_dataOut_payload_0_12483;
  reg        [7:0]    _zz_dataOut_payload_0_12484;
  reg        [7:0]    _zz_dataOut_payload_0_12485;
  reg        [7:0]    _zz_dataOut_payload_0_12486;
  reg        [7:0]    _zz_dataOut_payload_0_12487;
  reg        [7:0]    _zz_dataOut_payload_0_12488;
  reg        [7:0]    _zz_dataOut_payload_0_12489;
  reg        [7:0]    _zz_dataOut_payload_0_12490;
  reg        [7:0]    _zz_dataOut_payload_0_12491;
  reg        [7:0]    _zz_dataOut_payload_0_12492;
  reg        [7:0]    _zz_dataOut_payload_0_12493;
  reg        [7:0]    _zz_dataOut_payload_0_12494;
  reg        [7:0]    _zz_dataOut_payload_0_12495;
  reg        [7:0]    _zz_dataOut_payload_0_12496;
  reg        [7:0]    _zz_dataOut_payload_0_12497;
  reg        [7:0]    _zz_dataOut_payload_0_12498;
  reg        [7:0]    _zz_dataOut_payload_0_12499;
  reg        [7:0]    _zz_dataOut_payload_0_12500;
  reg        [7:0]    _zz_dataOut_payload_0_12501;
  reg        [7:0]    _zz_dataOut_payload_0_12502;
  reg        [7:0]    _zz_dataOut_payload_0_12503;
  reg        [7:0]    _zz_dataOut_payload_0_12504;
  reg        [7:0]    _zz_dataOut_payload_0_12505;
  reg        [7:0]    _zz_dataOut_payload_0_12506;
  reg        [7:0]    _zz_dataOut_payload_0_12507;
  reg        [7:0]    _zz_dataOut_payload_0_12508;
  reg        [7:0]    _zz_dataOut_payload_0_12509;
  reg        [7:0]    _zz_dataOut_payload_0_12510;
  reg        [7:0]    _zz_dataOut_payload_0_12511;
  reg        [7:0]    _zz_dataOut_payload_0_12512;
  reg        [7:0]    _zz_dataOut_payload_0_12513;
  reg        [7:0]    _zz_dataOut_payload_0_12514;
  reg        [7:0]    _zz_dataOut_payload_0_12515;
  reg        [7:0]    _zz_dataOut_payload_0_12516;
  reg        [7:0]    _zz_dataOut_payload_0_12517;
  reg        [7:0]    _zz_dataOut_payload_0_12518;
  reg        [7:0]    _zz_dataOut_payload_0_12519;
  reg        [7:0]    _zz_dataOut_payload_0_12520;
  reg        [7:0]    _zz_dataOut_payload_0_12521;
  reg        [7:0]    _zz_dataOut_payload_0_12522;
  reg        [7:0]    _zz_dataOut_payload_0_12523;
  reg        [7:0]    _zz_dataOut_payload_0_12524;
  reg        [7:0]    _zz_dataOut_payload_0_12525;
  reg        [7:0]    _zz_dataOut_payload_0_12526;
  reg        [7:0]    _zz_dataOut_payload_0_12527;
  wire                _zz_dataOut_payload_0_12528;
  wire       [7:0]    _zz_dataOut_payload_0_12529;
  wire       [7:0]    _zz_dataOut_payload_0_12530;
  wire                _zz_dataOut_payload_0_12531;
  wire       [7:0]    _zz_dataOut_payload_0_12532;
  wire       [7:0]    _zz_dataOut_payload_0_12533;
  wire                _zz_dataOut_payload_0_12534;
  wire       [7:0]    _zz_dataOut_payload_0_12535;
  wire       [7:0]    _zz_dataOut_payload_0_12536;
  wire                _zz_dataOut_payload_0_12537;
  wire       [7:0]    _zz_dataOut_payload_0_12538;
  wire       [7:0]    _zz_dataOut_payload_0_12539;
  wire                _zz_dataOut_payload_0_12540;
  wire       [7:0]    _zz_dataOut_payload_0_12541;
  wire       [7:0]    _zz_dataOut_payload_0_12542;
  wire                _zz_dataOut_payload_0_12543;
  wire       [7:0]    _zz_dataOut_payload_0_12544;
  wire       [7:0]    _zz_dataOut_payload_0_12545;
  wire                _zz_dataOut_payload_0_12546;
  wire       [7:0]    _zz_dataOut_payload_0_12547;
  wire       [7:0]    _zz_dataOut_payload_0_12548;
  wire                _zz_dataOut_payload_0_12549;
  wire       [7:0]    _zz_dataOut_payload_0_12550;
  wire       [7:0]    _zz_dataOut_payload_0_12551;
  wire                _zz_dataOut_payload_0_12552;
  wire       [7:0]    _zz_dataOut_payload_0_12553;
  wire       [7:0]    _zz_dataOut_payload_0_12554;
  wire                _zz_dataOut_payload_0_12555;
  wire       [7:0]    _zz_dataOut_payload_0_12556;
  wire       [7:0]    _zz_dataOut_payload_0_12557;
  wire                _zz_dataOut_payload_0_12558;
  wire       [7:0]    _zz_dataOut_payload_0_12559;
  wire       [7:0]    _zz_dataOut_payload_0_12560;
  wire                _zz_dataOut_payload_0_12561;
  wire       [7:0]    _zz_dataOut_payload_0_12562;
  wire       [7:0]    _zz_dataOut_payload_0_12563;
  wire                _zz_dataOut_payload_0_12564;
  wire       [7:0]    _zz_dataOut_payload_0_12565;
  wire       [7:0]    _zz_dataOut_payload_0_12566;
  wire                _zz_dataOut_payload_0_12567;
  wire       [7:0]    _zz_dataOut_payload_0_12568;
  wire       [7:0]    _zz_dataOut_payload_0_12569;
  wire                _zz_dataOut_payload_0_12570;
  wire       [7:0]    _zz_dataOut_payload_0_12571;
  wire       [7:0]    _zz_dataOut_payload_0_12572;
  wire                _zz_dataOut_payload_0_12573;
  wire       [7:0]    _zz_dataOut_payload_0_12574;
  wire       [7:0]    _zz_dataOut_payload_0_12575;
  wire                _zz_dataOut_payload_0_12576;
  wire       [7:0]    _zz_dataOut_payload_0_12577;
  wire       [7:0]    _zz_dataOut_payload_0_12578;
  wire                _zz_dataOut_payload_0_12579;
  wire       [7:0]    _zz_dataOut_payload_0_12580;
  wire       [7:0]    _zz_dataOut_payload_0_12581;
  wire                _zz_dataOut_payload_0_12582;
  wire       [7:0]    _zz_dataOut_payload_0_12583;
  wire       [7:0]    _zz_dataOut_payload_0_12584;
  wire                _zz_dataOut_payload_0_12585;
  wire       [7:0]    _zz_dataOut_payload_0_12586;
  wire       [7:0]    _zz_dataOut_payload_0_12587;
  wire                _zz_dataOut_payload_0_12588;
  wire       [7:0]    _zz_dataOut_payload_0_12589;
  wire       [7:0]    _zz_dataOut_payload_0_12590;
  wire                _zz_dataOut_payload_0_12591;
  wire       [7:0]    _zz_dataOut_payload_0_12592;
  wire       [7:0]    _zz_dataOut_payload_0_12593;
  wire                _zz_dataOut_payload_0_12594;
  wire       [7:0]    _zz_dataOut_payload_0_12595;
  wire       [7:0]    _zz_dataOut_payload_0_12596;
  wire                _zz_dataOut_payload_0_12597;
  wire       [7:0]    _zz_dataOut_payload_0_12598;
  wire       [7:0]    _zz_dataOut_payload_0_12599;
  wire                _zz_dataOut_payload_0_12600;
  wire       [7:0]    _zz_dataOut_payload_0_12601;
  wire       [7:0]    _zz_dataOut_payload_0_12602;
  wire                _zz_dataOut_payload_0_12603;
  wire       [7:0]    _zz_dataOut_payload_0_12604;
  wire       [7:0]    _zz_dataOut_payload_0_12605;
  wire                _zz_dataOut_payload_0_12606;
  wire       [7:0]    _zz_dataOut_payload_0_12607;
  wire       [7:0]    _zz_dataOut_payload_0_12608;
  wire                _zz_dataOut_payload_0_12609;
  wire       [7:0]    _zz_dataOut_payload_0_12610;
  wire       [7:0]    _zz_dataOut_payload_0_12611;
  wire                _zz_dataOut_payload_0_12612;
  wire       [7:0]    _zz_dataOut_payload_0_12613;
  wire       [7:0]    _zz_dataOut_payload_0_12614;
  wire                _zz_dataOut_payload_0_12615;
  wire       [7:0]    _zz_dataOut_payload_0_12616;
  wire       [7:0]    _zz_dataOut_payload_0_12617;
  wire                _zz_dataOut_payload_0_12618;
  wire                _zz_dataOut_payload_0_12619;
  reg        [7:0]    _zz_dataOut_payload_0_12620;
  reg        [7:0]    _zz_dataOut_payload_0_12621;
  reg        [7:0]    _zz_dataOut_payload_0_12622;
  reg        [7:0]    _zz_dataOut_payload_0_12623;
  wire                _zz_dataOut_payload_0_12624;
  wire       [7:0]    _zz_dataOut_payload_0_12625;
  wire       [7:0]    _zz_dataOut_payload_0_12626;
  wire                _zz_dataOut_payload_0_12627;
  wire       [7:0]    _zz_dataOut_payload_0_12628;
  wire       [7:0]    _zz_dataOut_payload_0_12629;
  wire                _zz_dataOut_payload_0_12630;
  wire                _zz_dataOut_payload_0_12631;
  reg        [7:0]    _zz_dataOut_payload_0_12632;
  reg        [7:0]    _zz_dataOut_payload_0_12633;
  reg        [7:0]    _zz_dataOut_payload_0_12634;
  reg        [7:0]    _zz_dataOut_payload_0_12635;
  reg        [7:0]    _zz_dataOut_payload_0_12636;
  reg        [7:0]    _zz_dataOut_payload_0_12637;
  reg        [7:0]    _zz_dataOut_payload_0_12638;
  reg        [7:0]    _zz_dataOut_payload_0_12639;
  reg        [7:0]    _zz_dataOut_payload_0_12640;
  reg        [7:0]    _zz_dataOut_payload_0_12641;
  reg        [7:0]    _zz_dataOut_payload_0_12642;
  reg        [7:0]    _zz_dataOut_payload_0_12643;
  wire                _zz_dataOut_payload_0_12644;
  wire       [7:0]    _zz_dataOut_payload_0_12645;
  wire       [7:0]    _zz_dataOut_payload_0_12646;
  wire                _zz_dataOut_payload_0_12647;
  wire       [7:0]    _zz_dataOut_payload_0_12648;
  wire       [7:0]    _zz_dataOut_payload_0_12649;
  wire                _zz_dataOut_payload_0_12650;
  wire       [7:0]    _zz_dataOut_payload_0_12651;
  wire       [7:0]    _zz_dataOut_payload_0_12652;
  wire                _zz_dataOut_payload_0_12653;
  wire       [7:0]    _zz_dataOut_payload_0_12654;
  wire       [7:0]    _zz_dataOut_payload_0_12655;
  wire                _zz_dataOut_payload_0_12656;
  wire       [7:0]    _zz_dataOut_payload_0_12657;
  wire       [7:0]    _zz_dataOut_payload_0_12658;
  wire                _zz_dataOut_payload_0_12659;
  wire       [7:0]    _zz_dataOut_payload_0_12660;
  wire       [7:0]    _zz_dataOut_payload_0_12661;
  wire                _zz_dataOut_payload_0_12662;
  wire                _zz_dataOut_payload_0_12663;
  reg        [7:0]    _zz_dataOut_payload_0_12664;
  reg        [7:0]    _zz_dataOut_payload_0_12665;
  reg        [7:0]    _zz_dataOut_payload_0_12666;
  reg        [7:0]    _zz_dataOut_payload_0_12667;
  wire                _zz_dataOut_payload_0_12668;
  wire       [7:0]    _zz_dataOut_payload_0_12669;
  wire       [7:0]    _zz_dataOut_payload_0_12670;
  wire                _zz_dataOut_payload_0_12671;
  wire       [7:0]    _zz_dataOut_payload_0_12672;
  wire       [7:0]    _zz_dataOut_payload_0_12673;
  wire                _zz_dataOut_payload_0_12674;
  wire                _zz_dataOut_payload_0_12675;
  reg        [7:0]    _zz_dataOut_payload_0_12676;
  reg        [7:0]    _zz_dataOut_payload_0_12677;
  reg        [7:0]    _zz_dataOut_payload_0_12678;
  reg        [7:0]    _zz_dataOut_payload_0_12679;
  reg        [7:0]    _zz_dataOut_payload_0_12680;
  reg        [7:0]    _zz_dataOut_payload_0_12681;
  reg        [7:0]    _zz_dataOut_payload_0_12682;
  reg        [7:0]    _zz_dataOut_payload_0_12683;
  reg        [7:0]    _zz_dataOut_payload_0_12684;
  reg        [7:0]    _zz_dataOut_payload_0_12685;
  reg        [7:0]    _zz_dataOut_payload_0_12686;
  reg        [7:0]    _zz_dataOut_payload_0_12687;
  reg        [7:0]    _zz_dataOut_payload_0_12688;
  reg        [7:0]    _zz_dataOut_payload_0_12689;
  reg        [7:0]    _zz_dataOut_payload_0_12690;
  reg        [7:0]    _zz_dataOut_payload_0_12691;
  reg        [7:0]    _zz_dataOut_payload_0_12692;
  reg        [7:0]    _zz_dataOut_payload_0_12693;
  reg        [7:0]    _zz_dataOut_payload_0_12694;
  reg        [7:0]    _zz_dataOut_payload_0_12695;
  reg        [7:0]    _zz_dataOut_payload_0_12696;
  reg        [7:0]    _zz_dataOut_payload_0_12697;
  reg        [7:0]    _zz_dataOut_payload_0_12698;
  reg        [7:0]    _zz_dataOut_payload_0_12699;
  reg        [7:0]    _zz_dataOut_payload_0_12700;
  reg        [7:0]    _zz_dataOut_payload_0_12701;
  reg        [7:0]    _zz_dataOut_payload_0_12702;
  reg        [7:0]    _zz_dataOut_payload_0_12703;
  wire                _zz_dataOut_payload_0_12704;
  wire       [7:0]    _zz_dataOut_payload_0_12705;
  wire       [7:0]    _zz_dataOut_payload_0_12706;
  wire                _zz_dataOut_payload_0_12707;
  wire       [7:0]    _zz_dataOut_payload_0_12708;
  wire       [7:0]    _zz_dataOut_payload_0_12709;
  wire                _zz_dataOut_payload_0_12710;
  wire       [7:0]    _zz_dataOut_payload_0_12711;
  wire       [7:0]    _zz_dataOut_payload_0_12712;
  wire                _zz_dataOut_payload_0_12713;
  wire       [7:0]    _zz_dataOut_payload_0_12714;
  wire       [7:0]    _zz_dataOut_payload_0_12715;
  wire                _zz_dataOut_payload_0_12716;
  wire       [7:0]    _zz_dataOut_payload_0_12717;
  wire       [7:0]    _zz_dataOut_payload_0_12718;
  wire                _zz_dataOut_payload_0_12719;
  wire       [7:0]    _zz_dataOut_payload_0_12720;
  wire       [7:0]    _zz_dataOut_payload_0_12721;
  wire                _zz_dataOut_payload_0_12722;
  wire       [7:0]    _zz_dataOut_payload_0_12723;
  wire       [7:0]    _zz_dataOut_payload_0_12724;
  wire                _zz_dataOut_payload_0_12725;
  wire       [7:0]    _zz_dataOut_payload_0_12726;
  wire       [7:0]    _zz_dataOut_payload_0_12727;
  wire                _zz_dataOut_payload_0_12728;
  wire       [7:0]    _zz_dataOut_payload_0_12729;
  wire       [7:0]    _zz_dataOut_payload_0_12730;
  wire                _zz_dataOut_payload_0_12731;
  wire       [7:0]    _zz_dataOut_payload_0_12732;
  wire       [7:0]    _zz_dataOut_payload_0_12733;
  wire                _zz_dataOut_payload_0_12734;
  wire       [7:0]    _zz_dataOut_payload_0_12735;
  wire       [7:0]    _zz_dataOut_payload_0_12736;
  wire                _zz_dataOut_payload_0_12737;
  wire       [7:0]    _zz_dataOut_payload_0_12738;
  wire       [7:0]    _zz_dataOut_payload_0_12739;
  wire                _zz_dataOut_payload_0_12740;
  wire       [7:0]    _zz_dataOut_payload_0_12741;
  wire       [7:0]    _zz_dataOut_payload_0_12742;
  wire                _zz_dataOut_payload_0_12743;
  wire       [7:0]    _zz_dataOut_payload_0_12744;
  wire       [7:0]    _zz_dataOut_payload_0_12745;
  wire                _zz_dataOut_payload_0_12746;
  wire                _zz_dataOut_payload_0_12747;
  reg        [7:0]    _zz_dataOut_payload_0_12748;
  reg        [7:0]    _zz_dataOut_payload_0_12749;
  reg        [7:0]    _zz_dataOut_payload_0_12750;
  reg        [7:0]    _zz_dataOut_payload_0_12751;
  wire                _zz_dataOut_payload_0_12752;
  wire       [7:0]    _zz_dataOut_payload_0_12753;
  wire       [7:0]    _zz_dataOut_payload_0_12754;
  wire                _zz_dataOut_payload_0_12755;
  wire       [7:0]    _zz_dataOut_payload_0_12756;
  wire       [7:0]    _zz_dataOut_payload_0_12757;
  wire                _zz_dataOut_payload_0_12758;
  wire                _zz_dataOut_payload_0_12759;
  reg        [7:0]    _zz_dataOut_payload_0_12760;
  reg        [7:0]    _zz_dataOut_payload_0_12761;
  reg        [7:0]    _zz_dataOut_payload_0_12762;
  reg        [7:0]    _zz_dataOut_payload_0_12763;
  reg        [7:0]    _zz_dataOut_payload_0_12764;
  reg        [7:0]    _zz_dataOut_payload_0_12765;
  reg        [7:0]    _zz_dataOut_payload_0_12766;
  reg        [7:0]    _zz_dataOut_payload_0_12767;
  reg        [7:0]    _zz_dataOut_payload_0_12768;
  reg        [7:0]    _zz_dataOut_payload_0_12769;
  reg        [7:0]    _zz_dataOut_payload_0_12770;
  reg        [7:0]    _zz_dataOut_payload_0_12771;
  wire                _zz_dataOut_payload_0_12772;
  wire       [7:0]    _zz_dataOut_payload_0_12773;
  wire       [7:0]    _zz_dataOut_payload_0_12774;
  wire                _zz_dataOut_payload_0_12775;
  wire       [7:0]    _zz_dataOut_payload_0_12776;
  wire       [7:0]    _zz_dataOut_payload_0_12777;
  wire                _zz_dataOut_payload_0_12778;
  wire       [7:0]    _zz_dataOut_payload_0_12779;
  wire       [7:0]    _zz_dataOut_payload_0_12780;
  wire                _zz_dataOut_payload_0_12781;
  wire       [7:0]    _zz_dataOut_payload_0_12782;
  wire       [7:0]    _zz_dataOut_payload_0_12783;
  wire                _zz_dataOut_payload_0_12784;
  wire       [7:0]    _zz_dataOut_payload_0_12785;
  wire       [7:0]    _zz_dataOut_payload_0_12786;
  wire                _zz_dataOut_payload_0_12787;
  wire       [7:0]    _zz_dataOut_payload_0_12788;
  wire       [7:0]    _zz_dataOut_payload_0_12789;
  wire                _zz_dataOut_payload_0_12790;
  wire                _zz_dataOut_payload_0_12791;
  reg        [7:0]    _zz_dataOut_payload_0_12792;
  reg        [7:0]    _zz_dataOut_payload_0_12793;
  reg        [7:0]    _zz_dataOut_payload_0_12794;
  reg        [7:0]    _zz_dataOut_payload_0_12795;
  wire                _zz_dataOut_payload_0_12796;
  wire       [7:0]    _zz_dataOut_payload_0_12797;
  wire       [7:0]    _zz_dataOut_payload_0_12798;
  wire                _zz_dataOut_payload_0_12799;
  wire       [7:0]    _zz_dataOut_payload_0_12800;
  wire       [7:0]    _zz_dataOut_payload_0_12801;
  wire                _zz_dataOut_payload_0_12802;
  wire                _zz_dataOut_payload_0_12803;
  reg        [7:0]    _zz_dataOut_payload_0_12804;
  reg        [7:0]    _zz_dataOut_payload_0_12805;
  reg        [7:0]    _zz_dataOut_payload_0_12806;
  reg        [7:0]    _zz_dataOut_payload_0_12807;
  reg        [7:0]    _zz_dataOut_payload_0_12808;
  reg        [7:0]    _zz_dataOut_payload_0_12809;
  reg        [7:0]    _zz_dataOut_payload_0_12810;
  reg        [7:0]    _zz_dataOut_payload_0_12811;
  reg        [7:0]    _zz_dataOut_payload_0_12812;
  reg        [7:0]    _zz_dataOut_payload_0_12813;
  reg        [7:0]    _zz_dataOut_payload_0_12814;
  reg        [7:0]    _zz_dataOut_payload_0_12815;
  reg        [7:0]    _zz_dataOut_payload_0_12816;
  reg        [7:0]    _zz_dataOut_payload_0_12817;
  reg        [7:0]    _zz_dataOut_payload_0_12818;
  reg        [7:0]    _zz_dataOut_payload_0_12819;
  reg        [7:0]    _zz_dataOut_payload_0_12820;
  reg        [7:0]    _zz_dataOut_payload_0_12821;
  reg        [7:0]    _zz_dataOut_payload_0_12822;
  reg        [7:0]    _zz_dataOut_payload_0_12823;
  reg        [7:0]    _zz_dataOut_payload_0_12824;
  reg        [7:0]    _zz_dataOut_payload_0_12825;
  reg        [7:0]    _zz_dataOut_payload_0_12826;
  reg        [7:0]    _zz_dataOut_payload_0_12827;
  reg        [7:0]    _zz_dataOut_payload_0_12828;
  reg        [7:0]    _zz_dataOut_payload_0_12829;
  reg        [7:0]    _zz_dataOut_payload_0_12830;
  reg        [7:0]    _zz_dataOut_payload_0_12831;
  reg        [7:0]    _zz_dataOut_payload_0_12832;
  reg        [7:0]    _zz_dataOut_payload_0_12833;
  reg        [7:0]    _zz_dataOut_payload_0_12834;
  reg        [7:0]    _zz_dataOut_payload_0_12835;
  reg        [7:0]    _zz_dataOut_payload_0_12836;
  reg        [7:0]    _zz_dataOut_payload_0_12837;
  reg        [7:0]    _zz_dataOut_payload_0_12838;
  reg        [7:0]    _zz_dataOut_payload_0_12839;
  reg        [7:0]    _zz_dataOut_payload_0_12840;
  reg        [7:0]    _zz_dataOut_payload_0_12841;
  reg        [7:0]    _zz_dataOut_payload_0_12842;
  reg        [7:0]    _zz_dataOut_payload_0_12843;
  reg        [7:0]    _zz_dataOut_payload_0_12844;
  reg        [7:0]    _zz_dataOut_payload_0_12845;
  reg        [7:0]    _zz_dataOut_payload_0_12846;
  reg        [7:0]    _zz_dataOut_payload_0_12847;
  reg        [7:0]    _zz_dataOut_payload_0_12848;
  reg        [7:0]    _zz_dataOut_payload_0_12849;
  reg        [7:0]    _zz_dataOut_payload_0_12850;
  reg        [7:0]    _zz_dataOut_payload_0_12851;
  reg        [7:0]    _zz_dataOut_payload_0_12852;
  reg        [7:0]    _zz_dataOut_payload_0_12853;
  reg        [7:0]    _zz_dataOut_payload_0_12854;
  reg        [7:0]    _zz_dataOut_payload_0_12855;
  reg        [7:0]    _zz_dataOut_payload_0_12856;
  reg        [7:0]    _zz_dataOut_payload_0_12857;
  reg        [7:0]    _zz_dataOut_payload_0_12858;
  reg        [7:0]    _zz_dataOut_payload_0_12859;
  reg        [7:0]    _zz_dataOut_payload_0_12860;
  reg        [7:0]    _zz_dataOut_payload_0_12861;
  reg        [7:0]    _zz_dataOut_payload_0_12862;
  reg        [7:0]    _zz_dataOut_payload_0_12863;
  reg        [7:0]    _zz_dataOut_payload_0_12864;
  reg        [7:0]    _zz_dataOut_payload_0_12865;
  reg        [7:0]    _zz_dataOut_payload_0_12866;
  reg        [7:0]    _zz_dataOut_payload_0_12867;
  reg        [7:0]    _zz_dataOut_payload_0_12868;
  reg        [7:0]    _zz_dataOut_payload_0_12869;
  reg        [7:0]    _zz_dataOut_payload_0_12870;
  reg        [7:0]    _zz_dataOut_payload_0_12871;
  reg        [7:0]    _zz_dataOut_payload_0_12872;
  reg        [7:0]    _zz_dataOut_payload_0_12873;
  reg        [7:0]    _zz_dataOut_payload_0_12874;
  reg        [7:0]    _zz_dataOut_payload_0_12875;
  reg        [7:0]    _zz_dataOut_payload_0_12876;
  reg        [7:0]    _zz_dataOut_payload_0_12877;
  reg        [7:0]    _zz_dataOut_payload_0_12878;
  reg        [7:0]    _zz_dataOut_payload_0_12879;
  reg        [7:0]    _zz_dataOut_payload_0_12880;
  reg        [7:0]    _zz_dataOut_payload_0_12881;
  reg        [7:0]    _zz_dataOut_payload_0_12882;
  reg        [7:0]    _zz_dataOut_payload_0_12883;
  reg        [7:0]    _zz_dataOut_payload_0_12884;
  reg        [7:0]    _zz_dataOut_payload_0_12885;
  reg        [7:0]    _zz_dataOut_payload_0_12886;
  reg        [7:0]    _zz_dataOut_payload_0_12887;
  reg        [7:0]    _zz_dataOut_payload_0_12888;
  reg        [7:0]    _zz_dataOut_payload_0_12889;
  reg        [7:0]    _zz_dataOut_payload_0_12890;
  reg        [7:0]    _zz_dataOut_payload_0_12891;
  reg        [7:0]    _zz_dataOut_payload_0_12892;
  reg        [7:0]    _zz_dataOut_payload_0_12893;
  reg        [7:0]    _zz_dataOut_payload_0_12894;
  reg        [7:0]    _zz_dataOut_payload_0_12895;
  reg        [7:0]    _zz_dataOut_payload_0_12896;
  reg        [7:0]    _zz_dataOut_payload_0_12897;
  reg        [7:0]    _zz_dataOut_payload_0_12898;
  reg        [7:0]    _zz_dataOut_payload_0_12899;
  reg        [7:0]    _zz_dataOut_payload_0_12900;
  reg        [7:0]    _zz_dataOut_payload_0_12901;
  reg        [7:0]    _zz_dataOut_payload_0_12902;
  reg        [7:0]    _zz_dataOut_payload_0_12903;
  reg        [7:0]    _zz_dataOut_payload_0_12904;
  reg        [7:0]    _zz_dataOut_payload_0_12905;
  reg        [7:0]    _zz_dataOut_payload_0_12906;
  reg        [7:0]    _zz_dataOut_payload_0_12907;
  reg        [7:0]    _zz_dataOut_payload_0_12908;
  reg        [7:0]    _zz_dataOut_payload_0_12909;
  reg        [7:0]    _zz_dataOut_payload_0_12910;
  reg        [7:0]    _zz_dataOut_payload_0_12911;
  reg        [7:0]    _zz_dataOut_payload_0_12912;
  reg        [7:0]    _zz_dataOut_payload_0_12913;
  reg        [7:0]    _zz_dataOut_payload_0_12914;
  reg        [7:0]    _zz_dataOut_payload_0_12915;
  reg        [7:0]    _zz_dataOut_payload_0_12916;
  reg        [7:0]    _zz_dataOut_payload_0_12917;
  reg        [7:0]    _zz_dataOut_payload_0_12918;
  reg        [7:0]    _zz_dataOut_payload_0_12919;
  reg        [7:0]    _zz_dataOut_payload_0_12920;
  reg        [7:0]    _zz_dataOut_payload_0_12921;
  reg        [7:0]    _zz_dataOut_payload_0_12922;
  reg        [7:0]    _zz_dataOut_payload_0_12923;
  reg        [7:0]    _zz_dataOut_payload_0_12924;
  reg        [7:0]    _zz_dataOut_payload_0_12925;
  reg        [7:0]    _zz_dataOut_payload_0_12926;
  reg        [7:0]    _zz_dataOut_payload_0_12927;
  wire                _zz_dataOut_payload_0_12928;
  wire       [7:0]    _zz_dataOut_payload_0_12929;
  wire       [7:0]    _zz_dataOut_payload_0_12930;
  wire                _zz_dataOut_payload_0_12931;
  wire       [7:0]    _zz_dataOut_payload_0_12932;
  wire       [7:0]    _zz_dataOut_payload_0_12933;
  wire                _zz_dataOut_payload_0_12934;
  wire       [7:0]    _zz_dataOut_payload_0_12935;
  wire       [7:0]    _zz_dataOut_payload_0_12936;
  wire                _zz_dataOut_payload_0_12937;
  wire       [7:0]    _zz_dataOut_payload_0_12938;
  wire       [7:0]    _zz_dataOut_payload_0_12939;
  wire                _zz_dataOut_payload_0_12940;
  wire       [7:0]    _zz_dataOut_payload_0_12941;
  wire       [7:0]    _zz_dataOut_payload_0_12942;
  wire                _zz_dataOut_payload_0_12943;
  wire       [7:0]    _zz_dataOut_payload_0_12944;
  wire       [7:0]    _zz_dataOut_payload_0_12945;
  wire                _zz_dataOut_payload_0_12946;
  wire       [7:0]    _zz_dataOut_payload_0_12947;
  wire       [7:0]    _zz_dataOut_payload_0_12948;
  wire                _zz_dataOut_payload_0_12949;
  wire       [7:0]    _zz_dataOut_payload_0_12950;
  wire       [7:0]    _zz_dataOut_payload_0_12951;
  wire                _zz_dataOut_payload_0_12952;
  wire       [7:0]    _zz_dataOut_payload_0_12953;
  wire       [7:0]    _zz_dataOut_payload_0_12954;
  wire                _zz_dataOut_payload_0_12955;
  wire       [7:0]    _zz_dataOut_payload_0_12956;
  wire       [7:0]    _zz_dataOut_payload_0_12957;
  wire                _zz_dataOut_payload_0_12958;
  wire       [7:0]    _zz_dataOut_payload_0_12959;
  wire       [7:0]    _zz_dataOut_payload_0_12960;
  wire                _zz_dataOut_payload_0_12961;
  wire       [7:0]    _zz_dataOut_payload_0_12962;
  wire       [7:0]    _zz_dataOut_payload_0_12963;
  wire                _zz_dataOut_payload_0_12964;
  wire       [7:0]    _zz_dataOut_payload_0_12965;
  wire       [7:0]    _zz_dataOut_payload_0_12966;
  wire                _zz_dataOut_payload_0_12967;
  wire       [7:0]    _zz_dataOut_payload_0_12968;
  wire       [7:0]    _zz_dataOut_payload_0_12969;
  wire                _zz_dataOut_payload_0_12970;
  wire       [7:0]    _zz_dataOut_payload_0_12971;
  wire       [7:0]    _zz_dataOut_payload_0_12972;
  wire                _zz_dataOut_payload_0_12973;
  wire       [7:0]    _zz_dataOut_payload_0_12974;
  wire       [7:0]    _zz_dataOut_payload_0_12975;
  wire                _zz_dataOut_payload_0_12976;
  wire       [7:0]    _zz_dataOut_payload_0_12977;
  wire       [7:0]    _zz_dataOut_payload_0_12978;
  wire                _zz_dataOut_payload_0_12979;
  wire       [7:0]    _zz_dataOut_payload_0_12980;
  wire       [7:0]    _zz_dataOut_payload_0_12981;
  wire                _zz_dataOut_payload_0_12982;
  wire       [7:0]    _zz_dataOut_payload_0_12983;
  wire       [7:0]    _zz_dataOut_payload_0_12984;
  wire                _zz_dataOut_payload_0_12985;
  wire       [7:0]    _zz_dataOut_payload_0_12986;
  wire       [7:0]    _zz_dataOut_payload_0_12987;
  wire                _zz_dataOut_payload_0_12988;
  wire       [7:0]    _zz_dataOut_payload_0_12989;
  wire       [7:0]    _zz_dataOut_payload_0_12990;
  wire                _zz_dataOut_payload_0_12991;
  wire       [7:0]    _zz_dataOut_payload_0_12992;
  wire       [7:0]    _zz_dataOut_payload_0_12993;
  wire                _zz_dataOut_payload_0_12994;
  wire       [7:0]    _zz_dataOut_payload_0_12995;
  wire       [7:0]    _zz_dataOut_payload_0_12996;
  wire                _zz_dataOut_payload_0_12997;
  wire       [7:0]    _zz_dataOut_payload_0_12998;
  wire       [7:0]    _zz_dataOut_payload_0_12999;
  wire                _zz_dataOut_payload_0_13000;
  wire       [7:0]    _zz_dataOut_payload_0_13001;
  wire       [7:0]    _zz_dataOut_payload_0_13002;
  wire                _zz_dataOut_payload_0_13003;
  wire       [7:0]    _zz_dataOut_payload_0_13004;
  wire       [7:0]    _zz_dataOut_payload_0_13005;
  wire                _zz_dataOut_payload_0_13006;
  wire       [7:0]    _zz_dataOut_payload_0_13007;
  wire       [7:0]    _zz_dataOut_payload_0_13008;
  wire                _zz_dataOut_payload_0_13009;
  wire       [7:0]    _zz_dataOut_payload_0_13010;
  wire       [7:0]    _zz_dataOut_payload_0_13011;
  wire                _zz_dataOut_payload_0_13012;
  wire       [7:0]    _zz_dataOut_payload_0_13013;
  wire       [7:0]    _zz_dataOut_payload_0_13014;
  wire                _zz_dataOut_payload_0_13015;
  wire       [7:0]    _zz_dataOut_payload_0_13016;
  wire       [7:0]    _zz_dataOut_payload_0_13017;
  wire                _zz_dataOut_payload_0_13018;
  wire       [7:0]    _zz_dataOut_payload_0_13019;
  wire       [7:0]    _zz_dataOut_payload_0_13020;
  wire                _zz_dataOut_payload_0_13021;
  wire       [7:0]    _zz_dataOut_payload_0_13022;
  wire       [7:0]    _zz_dataOut_payload_0_13023;
  wire                _zz_dataOut_payload_0_13024;
  wire       [7:0]    _zz_dataOut_payload_0_13025;
  wire       [7:0]    _zz_dataOut_payload_0_13026;
  wire                _zz_dataOut_payload_0_13027;
  wire       [7:0]    _zz_dataOut_payload_0_13028;
  wire       [7:0]    _zz_dataOut_payload_0_13029;
  wire                _zz_dataOut_payload_0_13030;
  wire       [7:0]    _zz_dataOut_payload_0_13031;
  wire       [7:0]    _zz_dataOut_payload_0_13032;
  wire                _zz_dataOut_payload_0_13033;
  wire       [7:0]    _zz_dataOut_payload_0_13034;
  wire       [7:0]    _zz_dataOut_payload_0_13035;
  wire                _zz_dataOut_payload_0_13036;
  wire       [7:0]    _zz_dataOut_payload_0_13037;
  wire       [7:0]    _zz_dataOut_payload_0_13038;
  wire                _zz_dataOut_payload_0_13039;
  wire       [7:0]    _zz_dataOut_payload_0_13040;
  wire       [7:0]    _zz_dataOut_payload_0_13041;
  wire                _zz_dataOut_payload_0_13042;
  wire       [7:0]    _zz_dataOut_payload_0_13043;
  wire       [7:0]    _zz_dataOut_payload_0_13044;
  wire                _zz_dataOut_payload_0_13045;
  wire       [7:0]    _zz_dataOut_payload_0_13046;
  wire       [7:0]    _zz_dataOut_payload_0_13047;
  wire                _zz_dataOut_payload_0_13048;
  wire       [7:0]    _zz_dataOut_payload_0_13049;
  wire       [7:0]    _zz_dataOut_payload_0_13050;
  wire                _zz_dataOut_payload_0_13051;
  wire       [7:0]    _zz_dataOut_payload_0_13052;
  wire       [7:0]    _zz_dataOut_payload_0_13053;
  wire                _zz_dataOut_payload_0_13054;
  wire       [7:0]    _zz_dataOut_payload_0_13055;
  wire       [7:0]    _zz_dataOut_payload_0_13056;
  wire                _zz_dataOut_payload_0_13057;
  wire       [7:0]    _zz_dataOut_payload_0_13058;
  wire       [7:0]    _zz_dataOut_payload_0_13059;
  wire                _zz_dataOut_payload_0_13060;
  wire       [7:0]    _zz_dataOut_payload_0_13061;
  wire       [7:0]    _zz_dataOut_payload_0_13062;
  wire                _zz_dataOut_payload_0_13063;
  wire       [7:0]    _zz_dataOut_payload_0_13064;
  wire       [7:0]    _zz_dataOut_payload_0_13065;
  wire                _zz_dataOut_payload_0_13066;
  wire       [7:0]    _zz_dataOut_payload_0_13067;
  wire       [7:0]    _zz_dataOut_payload_0_13068;
  wire                _zz_dataOut_payload_0_13069;
  wire       [7:0]    _zz_dataOut_payload_0_13070;
  wire       [7:0]    _zz_dataOut_payload_0_13071;
  wire                _zz_dataOut_payload_0_13072;
  wire       [7:0]    _zz_dataOut_payload_0_13073;
  wire       [7:0]    _zz_dataOut_payload_0_13074;
  wire                _zz_dataOut_payload_0_13075;
  wire       [7:0]    _zz_dataOut_payload_0_13076;
  wire       [7:0]    _zz_dataOut_payload_0_13077;
  wire                _zz_dataOut_payload_0_13078;
  wire       [7:0]    _zz_dataOut_payload_0_13079;
  wire       [7:0]    _zz_dataOut_payload_0_13080;
  wire                _zz_dataOut_payload_0_13081;
  wire       [7:0]    _zz_dataOut_payload_0_13082;
  wire       [7:0]    _zz_dataOut_payload_0_13083;
  wire                _zz_dataOut_payload_0_13084;
  wire       [7:0]    _zz_dataOut_payload_0_13085;
  wire       [7:0]    _zz_dataOut_payload_0_13086;
  wire                _zz_dataOut_payload_0_13087;
  wire       [7:0]    _zz_dataOut_payload_0_13088;
  wire       [7:0]    _zz_dataOut_payload_0_13089;
  wire                _zz_dataOut_payload_0_13090;
  wire       [7:0]    _zz_dataOut_payload_0_13091;
  wire       [7:0]    _zz_dataOut_payload_0_13092;
  wire                _zz_dataOut_payload_0_13093;
  wire       [7:0]    _zz_dataOut_payload_0_13094;
  wire       [7:0]    _zz_dataOut_payload_0_13095;
  wire                _zz_dataOut_payload_0_13096;
  wire       [7:0]    _zz_dataOut_payload_0_13097;
  wire       [7:0]    _zz_dataOut_payload_0_13098;
  wire                _zz_dataOut_payload_0_13099;
  wire       [7:0]    _zz_dataOut_payload_0_13100;
  wire       [7:0]    _zz_dataOut_payload_0_13101;
  wire                _zz_dataOut_payload_0_13102;
  wire       [7:0]    _zz_dataOut_payload_0_13103;
  wire       [7:0]    _zz_dataOut_payload_0_13104;
  wire                _zz_dataOut_payload_0_13105;
  wire       [7:0]    _zz_dataOut_payload_0_13106;
  wire       [7:0]    _zz_dataOut_payload_0_13107;
  wire                _zz_dataOut_payload_0_13108;
  wire       [7:0]    _zz_dataOut_payload_0_13109;
  wire       [7:0]    _zz_dataOut_payload_0_13110;
  wire                _zz_dataOut_payload_0_13111;
  wire       [7:0]    _zz_dataOut_payload_0_13112;
  wire       [7:0]    _zz_dataOut_payload_0_13113;
  wire                _zz_dataOut_payload_0_13114;
  wire                _zz_dataOut_payload_0_13115;
  reg        [7:0]    _zz_dataOut_payload_0_13116;
  reg        [7:0]    _zz_dataOut_payload_0_13117;
  reg        [7:0]    _zz_dataOut_payload_0_13118;
  reg        [7:0]    _zz_dataOut_payload_0_13119;
  wire                _zz_dataOut_payload_0_13120;
  wire       [7:0]    _zz_dataOut_payload_0_13121;
  wire       [7:0]    _zz_dataOut_payload_0_13122;
  wire                _zz_dataOut_payload_0_13123;
  wire       [7:0]    _zz_dataOut_payload_0_13124;
  wire       [7:0]    _zz_dataOut_payload_0_13125;
  wire                _zz_dataOut_payload_0_13126;
  wire                _zz_dataOut_payload_0_13127;
  reg        [7:0]    _zz_dataOut_payload_0_13128;
  reg        [7:0]    _zz_dataOut_payload_0_13129;
  reg        [7:0]    _zz_dataOut_payload_0_13130;
  reg        [7:0]    _zz_dataOut_payload_0_13131;
  reg        [7:0]    _zz_dataOut_payload_0_13132;
  reg        [7:0]    _zz_dataOut_payload_0_13133;
  reg        [7:0]    _zz_dataOut_payload_0_13134;
  reg        [7:0]    _zz_dataOut_payload_0_13135;
  reg        [7:0]    _zz_dataOut_payload_0_13136;
  reg        [7:0]    _zz_dataOut_payload_0_13137;
  reg        [7:0]    _zz_dataOut_payload_0_13138;
  reg        [7:0]    _zz_dataOut_payload_0_13139;
  wire                _zz_dataOut_payload_0_13140;
  wire       [7:0]    _zz_dataOut_payload_0_13141;
  wire       [7:0]    _zz_dataOut_payload_0_13142;
  wire                _zz_dataOut_payload_0_13143;
  wire       [7:0]    _zz_dataOut_payload_0_13144;
  wire       [7:0]    _zz_dataOut_payload_0_13145;
  wire                _zz_dataOut_payload_0_13146;
  wire       [7:0]    _zz_dataOut_payload_0_13147;
  wire       [7:0]    _zz_dataOut_payload_0_13148;
  wire                _zz_dataOut_payload_0_13149;
  wire       [7:0]    _zz_dataOut_payload_0_13150;
  wire       [7:0]    _zz_dataOut_payload_0_13151;
  wire                _zz_dataOut_payload_0_13152;
  wire       [7:0]    _zz_dataOut_payload_0_13153;
  wire       [7:0]    _zz_dataOut_payload_0_13154;
  wire                _zz_dataOut_payload_0_13155;
  wire       [7:0]    _zz_dataOut_payload_0_13156;
  wire       [7:0]    _zz_dataOut_payload_0_13157;
  wire                _zz_dataOut_payload_0_13158;
  wire                _zz_dataOut_payload_0_13159;
  reg        [7:0]    _zz_dataOut_payload_0_13160;
  reg        [7:0]    _zz_dataOut_payload_0_13161;
  reg        [7:0]    _zz_dataOut_payload_0_13162;
  reg        [7:0]    _zz_dataOut_payload_0_13163;
  wire                _zz_dataOut_payload_0_13164;
  wire       [7:0]    _zz_dataOut_payload_0_13165;
  wire       [7:0]    _zz_dataOut_payload_0_13166;
  wire                _zz_dataOut_payload_0_13167;
  wire       [7:0]    _zz_dataOut_payload_0_13168;
  wire       [7:0]    _zz_dataOut_payload_0_13169;
  wire                _zz_dataOut_payload_0_13170;
  wire                _zz_dataOut_payload_0_13171;
  reg        [7:0]    _zz_dataOut_payload_0_13172;
  reg        [7:0]    _zz_dataOut_payload_0_13173;
  reg        [7:0]    _zz_dataOut_payload_0_13174;
  reg        [7:0]    _zz_dataOut_payload_0_13175;
  reg        [7:0]    _zz_dataOut_payload_0_13176;
  reg        [7:0]    _zz_dataOut_payload_0_13177;
  reg        [7:0]    _zz_dataOut_payload_0_13178;
  reg        [7:0]    _zz_dataOut_payload_0_13179;
  reg        [7:0]    _zz_dataOut_payload_0_13180;
  reg        [7:0]    _zz_dataOut_payload_0_13181;
  reg        [7:0]    _zz_dataOut_payload_0_13182;
  reg        [7:0]    _zz_dataOut_payload_0_13183;
  reg        [7:0]    _zz_dataOut_payload_0_13184;
  reg        [7:0]    _zz_dataOut_payload_0_13185;
  reg        [7:0]    _zz_dataOut_payload_0_13186;
  reg        [7:0]    _zz_dataOut_payload_0_13187;
  reg        [7:0]    _zz_dataOut_payload_0_13188;
  reg        [7:0]    _zz_dataOut_payload_0_13189;
  reg        [7:0]    _zz_dataOut_payload_0_13190;
  reg        [7:0]    _zz_dataOut_payload_0_13191;
  reg        [7:0]    _zz_dataOut_payload_0_13192;
  reg        [7:0]    _zz_dataOut_payload_0_13193;
  reg        [7:0]    _zz_dataOut_payload_0_13194;
  reg        [7:0]    _zz_dataOut_payload_0_13195;
  reg        [7:0]    _zz_dataOut_payload_0_13196;
  reg        [7:0]    _zz_dataOut_payload_0_13197;
  reg        [7:0]    _zz_dataOut_payload_0_13198;
  reg        [7:0]    _zz_dataOut_payload_0_13199;
  wire                _zz_dataOut_payload_0_13200;
  wire       [7:0]    _zz_dataOut_payload_0_13201;
  wire       [7:0]    _zz_dataOut_payload_0_13202;
  wire                _zz_dataOut_payload_0_13203;
  wire       [7:0]    _zz_dataOut_payload_0_13204;
  wire       [7:0]    _zz_dataOut_payload_0_13205;
  wire                _zz_dataOut_payload_0_13206;
  wire       [7:0]    _zz_dataOut_payload_0_13207;
  wire       [7:0]    _zz_dataOut_payload_0_13208;
  wire                _zz_dataOut_payload_0_13209;
  wire       [7:0]    _zz_dataOut_payload_0_13210;
  wire       [7:0]    _zz_dataOut_payload_0_13211;
  wire                _zz_dataOut_payload_0_13212;
  wire       [7:0]    _zz_dataOut_payload_0_13213;
  wire       [7:0]    _zz_dataOut_payload_0_13214;
  wire                _zz_dataOut_payload_0_13215;
  wire       [7:0]    _zz_dataOut_payload_0_13216;
  wire       [7:0]    _zz_dataOut_payload_0_13217;
  wire                _zz_dataOut_payload_0_13218;
  wire       [7:0]    _zz_dataOut_payload_0_13219;
  wire       [7:0]    _zz_dataOut_payload_0_13220;
  wire                _zz_dataOut_payload_0_13221;
  wire       [7:0]    _zz_dataOut_payload_0_13222;
  wire       [7:0]    _zz_dataOut_payload_0_13223;
  wire                _zz_dataOut_payload_0_13224;
  wire       [7:0]    _zz_dataOut_payload_0_13225;
  wire       [7:0]    _zz_dataOut_payload_0_13226;
  wire                _zz_dataOut_payload_0_13227;
  wire       [7:0]    _zz_dataOut_payload_0_13228;
  wire       [7:0]    _zz_dataOut_payload_0_13229;
  wire                _zz_dataOut_payload_0_13230;
  wire       [7:0]    _zz_dataOut_payload_0_13231;
  wire       [7:0]    _zz_dataOut_payload_0_13232;
  wire                _zz_dataOut_payload_0_13233;
  wire       [7:0]    _zz_dataOut_payload_0_13234;
  wire       [7:0]    _zz_dataOut_payload_0_13235;
  wire                _zz_dataOut_payload_0_13236;
  wire       [7:0]    _zz_dataOut_payload_0_13237;
  wire       [7:0]    _zz_dataOut_payload_0_13238;
  wire                _zz_dataOut_payload_0_13239;
  wire       [7:0]    _zz_dataOut_payload_0_13240;
  wire       [7:0]    _zz_dataOut_payload_0_13241;
  wire                _zz_dataOut_payload_0_13242;
  wire                _zz_dataOut_payload_0_13243;
  reg        [7:0]    _zz_dataOut_payload_0_13244;
  reg        [7:0]    _zz_dataOut_payload_0_13245;
  reg        [7:0]    _zz_dataOut_payload_0_13246;
  reg        [7:0]    _zz_dataOut_payload_0_13247;
  wire                _zz_dataOut_payload_0_13248;
  wire       [7:0]    _zz_dataOut_payload_0_13249;
  wire       [7:0]    _zz_dataOut_payload_0_13250;
  wire                _zz_dataOut_payload_0_13251;
  wire       [7:0]    _zz_dataOut_payload_0_13252;
  wire       [7:0]    _zz_dataOut_payload_0_13253;
  wire                _zz_dataOut_payload_0_13254;
  wire                _zz_dataOut_payload_0_13255;
  reg        [7:0]    _zz_dataOut_payload_0_13256;
  reg        [7:0]    _zz_dataOut_payload_0_13257;
  reg        [7:0]    _zz_dataOut_payload_0_13258;
  reg        [7:0]    _zz_dataOut_payload_0_13259;
  reg        [7:0]    _zz_dataOut_payload_0_13260;
  reg        [7:0]    _zz_dataOut_payload_0_13261;
  reg        [7:0]    _zz_dataOut_payload_0_13262;
  reg        [7:0]    _zz_dataOut_payload_0_13263;
  reg        [7:0]    _zz_dataOut_payload_0_13264;
  reg        [7:0]    _zz_dataOut_payload_0_13265;
  reg        [7:0]    _zz_dataOut_payload_0_13266;
  reg        [7:0]    _zz_dataOut_payload_0_13267;
  wire                _zz_dataOut_payload_0_13268;
  wire       [7:0]    _zz_dataOut_payload_0_13269;
  wire       [7:0]    _zz_dataOut_payload_0_13270;
  wire                _zz_dataOut_payload_0_13271;
  wire       [7:0]    _zz_dataOut_payload_0_13272;
  wire       [7:0]    _zz_dataOut_payload_0_13273;
  wire                _zz_dataOut_payload_0_13274;
  wire       [7:0]    _zz_dataOut_payload_0_13275;
  wire       [7:0]    _zz_dataOut_payload_0_13276;
  wire                _zz_dataOut_payload_0_13277;
  wire       [7:0]    _zz_dataOut_payload_0_13278;
  wire       [7:0]    _zz_dataOut_payload_0_13279;
  wire                _zz_dataOut_payload_0_13280;
  wire       [7:0]    _zz_dataOut_payload_0_13281;
  wire       [7:0]    _zz_dataOut_payload_0_13282;
  wire                _zz_dataOut_payload_0_13283;
  wire       [7:0]    _zz_dataOut_payload_0_13284;
  wire       [7:0]    _zz_dataOut_payload_0_13285;
  wire                _zz_dataOut_payload_0_13286;
  wire                _zz_dataOut_payload_0_13287;
  reg        [7:0]    _zz_dataOut_payload_0_13288;
  reg        [7:0]    _zz_dataOut_payload_0_13289;
  reg        [7:0]    _zz_dataOut_payload_0_13290;
  reg        [7:0]    _zz_dataOut_payload_0_13291;
  wire                _zz_dataOut_payload_0_13292;
  wire       [7:0]    _zz_dataOut_payload_0_13293;
  wire       [7:0]    _zz_dataOut_payload_0_13294;
  wire                _zz_dataOut_payload_0_13295;
  wire       [7:0]    _zz_dataOut_payload_0_13296;
  wire       [7:0]    _zz_dataOut_payload_0_13297;
  wire                _zz_dataOut_payload_0_13298;
  wire                _zz_dataOut_payload_0_13299;
  reg        [7:0]    _zz_dataOut_payload_0_13300;
  reg        [7:0]    _zz_dataOut_payload_0_13301;
  reg        [7:0]    _zz_dataOut_payload_0_13302;
  reg        [7:0]    _zz_dataOut_payload_0_13303;
  reg        [7:0]    _zz_dataOut_payload_0_13304;
  reg        [7:0]    _zz_dataOut_payload_0_13305;
  reg        [7:0]    _zz_dataOut_payload_0_13306;
  reg        [7:0]    _zz_dataOut_payload_0_13307;
  reg        [7:0]    _zz_dataOut_payload_0_13308;
  reg        [7:0]    _zz_dataOut_payload_0_13309;
  reg        [7:0]    _zz_dataOut_payload_0_13310;
  reg        [7:0]    _zz_dataOut_payload_0_13311;
  reg        [7:0]    _zz_dataOut_payload_0_13312;
  reg        [7:0]    _zz_dataOut_payload_0_13313;
  reg        [7:0]    _zz_dataOut_payload_0_13314;
  reg        [7:0]    _zz_dataOut_payload_0_13315;
  reg        [7:0]    _zz_dataOut_payload_0_13316;
  reg        [7:0]    _zz_dataOut_payload_0_13317;
  reg        [7:0]    _zz_dataOut_payload_0_13318;
  reg        [7:0]    _zz_dataOut_payload_0_13319;
  reg        [7:0]    _zz_dataOut_payload_0_13320;
  reg        [7:0]    _zz_dataOut_payload_0_13321;
  reg        [7:0]    _zz_dataOut_payload_0_13322;
  reg        [7:0]    _zz_dataOut_payload_0_13323;
  reg        [7:0]    _zz_dataOut_payload_0_13324;
  reg        [7:0]    _zz_dataOut_payload_0_13325;
  reg        [7:0]    _zz_dataOut_payload_0_13326;
  reg        [7:0]    _zz_dataOut_payload_0_13327;
  reg        [7:0]    _zz_dataOut_payload_0_13328;
  reg        [7:0]    _zz_dataOut_payload_0_13329;
  reg        [7:0]    _zz_dataOut_payload_0_13330;
  reg        [7:0]    _zz_dataOut_payload_0_13331;
  reg        [7:0]    _zz_dataOut_payload_0_13332;
  reg        [7:0]    _zz_dataOut_payload_0_13333;
  reg        [7:0]    _zz_dataOut_payload_0_13334;
  reg        [7:0]    _zz_dataOut_payload_0_13335;
  reg        [7:0]    _zz_dataOut_payload_0_13336;
  reg        [7:0]    _zz_dataOut_payload_0_13337;
  reg        [7:0]    _zz_dataOut_payload_0_13338;
  reg        [7:0]    _zz_dataOut_payload_0_13339;
  reg        [7:0]    _zz_dataOut_payload_0_13340;
  reg        [7:0]    _zz_dataOut_payload_0_13341;
  reg        [7:0]    _zz_dataOut_payload_0_13342;
  reg        [7:0]    _zz_dataOut_payload_0_13343;
  reg        [7:0]    _zz_dataOut_payload_0_13344;
  reg        [7:0]    _zz_dataOut_payload_0_13345;
  reg        [7:0]    _zz_dataOut_payload_0_13346;
  reg        [7:0]    _zz_dataOut_payload_0_13347;
  reg        [7:0]    _zz_dataOut_payload_0_13348;
  reg        [7:0]    _zz_dataOut_payload_0_13349;
  reg        [7:0]    _zz_dataOut_payload_0_13350;
  reg        [7:0]    _zz_dataOut_payload_0_13351;
  reg        [7:0]    _zz_dataOut_payload_0_13352;
  reg        [7:0]    _zz_dataOut_payload_0_13353;
  reg        [7:0]    _zz_dataOut_payload_0_13354;
  reg        [7:0]    _zz_dataOut_payload_0_13355;
  reg        [7:0]    _zz_dataOut_payload_0_13356;
  reg        [7:0]    _zz_dataOut_payload_0_13357;
  reg        [7:0]    _zz_dataOut_payload_0_13358;
  reg        [7:0]    _zz_dataOut_payload_0_13359;
  wire                _zz_dataOut_payload_0_13360;
  wire       [7:0]    _zz_dataOut_payload_0_13361;
  wire       [7:0]    _zz_dataOut_payload_0_13362;
  wire                _zz_dataOut_payload_0_13363;
  wire       [7:0]    _zz_dataOut_payload_0_13364;
  wire       [7:0]    _zz_dataOut_payload_0_13365;
  wire                _zz_dataOut_payload_0_13366;
  wire       [7:0]    _zz_dataOut_payload_0_13367;
  wire       [7:0]    _zz_dataOut_payload_0_13368;
  wire                _zz_dataOut_payload_0_13369;
  wire       [7:0]    _zz_dataOut_payload_0_13370;
  wire       [7:0]    _zz_dataOut_payload_0_13371;
  wire                _zz_dataOut_payload_0_13372;
  wire       [7:0]    _zz_dataOut_payload_0_13373;
  wire       [7:0]    _zz_dataOut_payload_0_13374;
  wire                _zz_dataOut_payload_0_13375;
  wire       [7:0]    _zz_dataOut_payload_0_13376;
  wire       [7:0]    _zz_dataOut_payload_0_13377;
  wire                _zz_dataOut_payload_0_13378;
  wire       [7:0]    _zz_dataOut_payload_0_13379;
  wire       [7:0]    _zz_dataOut_payload_0_13380;
  wire                _zz_dataOut_payload_0_13381;
  wire       [7:0]    _zz_dataOut_payload_0_13382;
  wire       [7:0]    _zz_dataOut_payload_0_13383;
  wire                _zz_dataOut_payload_0_13384;
  wire       [7:0]    _zz_dataOut_payload_0_13385;
  wire       [7:0]    _zz_dataOut_payload_0_13386;
  wire                _zz_dataOut_payload_0_13387;
  wire       [7:0]    _zz_dataOut_payload_0_13388;
  wire       [7:0]    _zz_dataOut_payload_0_13389;
  wire                _zz_dataOut_payload_0_13390;
  wire       [7:0]    _zz_dataOut_payload_0_13391;
  wire       [7:0]    _zz_dataOut_payload_0_13392;
  wire                _zz_dataOut_payload_0_13393;
  wire       [7:0]    _zz_dataOut_payload_0_13394;
  wire       [7:0]    _zz_dataOut_payload_0_13395;
  wire                _zz_dataOut_payload_0_13396;
  wire       [7:0]    _zz_dataOut_payload_0_13397;
  wire       [7:0]    _zz_dataOut_payload_0_13398;
  wire                _zz_dataOut_payload_0_13399;
  wire       [7:0]    _zz_dataOut_payload_0_13400;
  wire       [7:0]    _zz_dataOut_payload_0_13401;
  wire                _zz_dataOut_payload_0_13402;
  wire       [7:0]    _zz_dataOut_payload_0_13403;
  wire       [7:0]    _zz_dataOut_payload_0_13404;
  wire                _zz_dataOut_payload_0_13405;
  wire       [7:0]    _zz_dataOut_payload_0_13406;
  wire       [7:0]    _zz_dataOut_payload_0_13407;
  wire                _zz_dataOut_payload_0_13408;
  wire       [7:0]    _zz_dataOut_payload_0_13409;
  wire       [7:0]    _zz_dataOut_payload_0_13410;
  wire                _zz_dataOut_payload_0_13411;
  wire       [7:0]    _zz_dataOut_payload_0_13412;
  wire       [7:0]    _zz_dataOut_payload_0_13413;
  wire                _zz_dataOut_payload_0_13414;
  wire       [7:0]    _zz_dataOut_payload_0_13415;
  wire       [7:0]    _zz_dataOut_payload_0_13416;
  wire                _zz_dataOut_payload_0_13417;
  wire       [7:0]    _zz_dataOut_payload_0_13418;
  wire       [7:0]    _zz_dataOut_payload_0_13419;
  wire                _zz_dataOut_payload_0_13420;
  wire       [7:0]    _zz_dataOut_payload_0_13421;
  wire       [7:0]    _zz_dataOut_payload_0_13422;
  wire                _zz_dataOut_payload_0_13423;
  wire       [7:0]    _zz_dataOut_payload_0_13424;
  wire       [7:0]    _zz_dataOut_payload_0_13425;
  wire                _zz_dataOut_payload_0_13426;
  wire       [7:0]    _zz_dataOut_payload_0_13427;
  wire       [7:0]    _zz_dataOut_payload_0_13428;
  wire                _zz_dataOut_payload_0_13429;
  wire       [7:0]    _zz_dataOut_payload_0_13430;
  wire       [7:0]    _zz_dataOut_payload_0_13431;
  wire                _zz_dataOut_payload_0_13432;
  wire       [7:0]    _zz_dataOut_payload_0_13433;
  wire       [7:0]    _zz_dataOut_payload_0_13434;
  wire                _zz_dataOut_payload_0_13435;
  wire       [7:0]    _zz_dataOut_payload_0_13436;
  wire       [7:0]    _zz_dataOut_payload_0_13437;
  wire                _zz_dataOut_payload_0_13438;
  wire       [7:0]    _zz_dataOut_payload_0_13439;
  wire       [7:0]    _zz_dataOut_payload_0_13440;
  wire                _zz_dataOut_payload_0_13441;
  wire       [7:0]    _zz_dataOut_payload_0_13442;
  wire       [7:0]    _zz_dataOut_payload_0_13443;
  wire                _zz_dataOut_payload_0_13444;
  wire       [7:0]    _zz_dataOut_payload_0_13445;
  wire       [7:0]    _zz_dataOut_payload_0_13446;
  wire                _zz_dataOut_payload_0_13447;
  wire       [7:0]    _zz_dataOut_payload_0_13448;
  wire       [7:0]    _zz_dataOut_payload_0_13449;
  wire                _zz_dataOut_payload_0_13450;
  wire                _zz_dataOut_payload_0_13451;
  reg        [7:0]    _zz_dataOut_payload_0_13452;
  reg        [7:0]    _zz_dataOut_payload_0_13453;
  reg        [7:0]    _zz_dataOut_payload_0_13454;
  reg        [7:0]    _zz_dataOut_payload_0_13455;
  wire                _zz_dataOut_payload_0_13456;
  wire       [7:0]    _zz_dataOut_payload_0_13457;
  wire       [7:0]    _zz_dataOut_payload_0_13458;
  wire                _zz_dataOut_payload_0_13459;
  wire       [7:0]    _zz_dataOut_payload_0_13460;
  wire       [7:0]    _zz_dataOut_payload_0_13461;
  wire                _zz_dataOut_payload_0_13462;
  wire                _zz_dataOut_payload_0_13463;
  reg        [7:0]    _zz_dataOut_payload_0_13464;
  reg        [7:0]    _zz_dataOut_payload_0_13465;
  reg        [7:0]    _zz_dataOut_payload_0_13466;
  reg        [7:0]    _zz_dataOut_payload_0_13467;
  reg        [7:0]    _zz_dataOut_payload_0_13468;
  reg        [7:0]    _zz_dataOut_payload_0_13469;
  reg        [7:0]    _zz_dataOut_payload_0_13470;
  reg        [7:0]    _zz_dataOut_payload_0_13471;
  reg        [7:0]    _zz_dataOut_payload_0_13472;
  reg        [7:0]    _zz_dataOut_payload_0_13473;
  reg        [7:0]    _zz_dataOut_payload_0_13474;
  reg        [7:0]    _zz_dataOut_payload_0_13475;
  wire                _zz_dataOut_payload_0_13476;
  wire       [7:0]    _zz_dataOut_payload_0_13477;
  wire       [7:0]    _zz_dataOut_payload_0_13478;
  wire                _zz_dataOut_payload_0_13479;
  wire       [7:0]    _zz_dataOut_payload_0_13480;
  wire       [7:0]    _zz_dataOut_payload_0_13481;
  wire                _zz_dataOut_payload_0_13482;
  wire       [7:0]    _zz_dataOut_payload_0_13483;
  wire       [7:0]    _zz_dataOut_payload_0_13484;
  wire                _zz_dataOut_payload_0_13485;
  wire       [7:0]    _zz_dataOut_payload_0_13486;
  wire       [7:0]    _zz_dataOut_payload_0_13487;
  wire                _zz_dataOut_payload_0_13488;
  wire       [7:0]    _zz_dataOut_payload_0_13489;
  wire       [7:0]    _zz_dataOut_payload_0_13490;
  wire                _zz_dataOut_payload_0_13491;
  wire       [7:0]    _zz_dataOut_payload_0_13492;
  wire       [7:0]    _zz_dataOut_payload_0_13493;
  wire                _zz_dataOut_payload_0_13494;
  wire                _zz_dataOut_payload_0_13495;
  reg        [7:0]    _zz_dataOut_payload_0_13496;
  reg        [7:0]    _zz_dataOut_payload_0_13497;
  reg        [7:0]    _zz_dataOut_payload_0_13498;
  reg        [7:0]    _zz_dataOut_payload_0_13499;
  wire                _zz_dataOut_payload_0_13500;
  wire       [7:0]    _zz_dataOut_payload_0_13501;
  wire       [7:0]    _zz_dataOut_payload_0_13502;
  wire                _zz_dataOut_payload_0_13503;
  wire       [7:0]    _zz_dataOut_payload_0_13504;
  wire       [7:0]    _zz_dataOut_payload_0_13505;
  wire                _zz_dataOut_payload_0_13506;
  wire                _zz_dataOut_payload_0_13507;
  reg        [7:0]    _zz_dataOut_payload_0_13508;
  reg        [7:0]    _zz_dataOut_payload_0_13509;
  reg        [7:0]    _zz_dataOut_payload_0_13510;
  reg        [7:0]    _zz_dataOut_payload_0_13511;
  reg        [7:0]    _zz_dataOut_payload_0_13512;
  reg        [7:0]    _zz_dataOut_payload_0_13513;
  reg        [7:0]    _zz_dataOut_payload_0_13514;
  reg        [7:0]    _zz_dataOut_payload_0_13515;
  reg        [7:0]    _zz_dataOut_payload_0_13516;
  reg        [7:0]    _zz_dataOut_payload_0_13517;
  reg        [7:0]    _zz_dataOut_payload_0_13518;
  reg        [7:0]    _zz_dataOut_payload_0_13519;
  reg        [7:0]    _zz_dataOut_payload_0_13520;
  reg        [7:0]    _zz_dataOut_payload_0_13521;
  reg        [7:0]    _zz_dataOut_payload_0_13522;
  reg        [7:0]    _zz_dataOut_payload_0_13523;
  reg        [7:0]    _zz_dataOut_payload_0_13524;
  reg        [7:0]    _zz_dataOut_payload_0_13525;
  reg        [7:0]    _zz_dataOut_payload_0_13526;
  reg        [7:0]    _zz_dataOut_payload_0_13527;
  reg        [7:0]    _zz_dataOut_payload_0_13528;
  reg        [7:0]    _zz_dataOut_payload_0_13529;
  reg        [7:0]    _zz_dataOut_payload_0_13530;
  reg        [7:0]    _zz_dataOut_payload_0_13531;
  reg        [7:0]    _zz_dataOut_payload_0_13532;
  reg        [7:0]    _zz_dataOut_payload_0_13533;
  reg        [7:0]    _zz_dataOut_payload_0_13534;
  reg        [7:0]    _zz_dataOut_payload_0_13535;
  wire                _zz_dataOut_payload_0_13536;
  wire       [7:0]    _zz_dataOut_payload_0_13537;
  wire       [7:0]    _zz_dataOut_payload_0_13538;
  wire                _zz_dataOut_payload_0_13539;
  wire       [7:0]    _zz_dataOut_payload_0_13540;
  wire       [7:0]    _zz_dataOut_payload_0_13541;
  wire                _zz_dataOut_payload_0_13542;
  wire       [7:0]    _zz_dataOut_payload_0_13543;
  wire       [7:0]    _zz_dataOut_payload_0_13544;
  wire                _zz_dataOut_payload_0_13545;
  wire       [7:0]    _zz_dataOut_payload_0_13546;
  wire       [7:0]    _zz_dataOut_payload_0_13547;
  wire                _zz_dataOut_payload_0_13548;
  wire       [7:0]    _zz_dataOut_payload_0_13549;
  wire       [7:0]    _zz_dataOut_payload_0_13550;
  wire                _zz_dataOut_payload_0_13551;
  wire       [7:0]    _zz_dataOut_payload_0_13552;
  wire       [7:0]    _zz_dataOut_payload_0_13553;
  wire                _zz_dataOut_payload_0_13554;
  wire       [7:0]    _zz_dataOut_payload_0_13555;
  wire       [7:0]    _zz_dataOut_payload_0_13556;
  wire                _zz_dataOut_payload_0_13557;
  wire       [7:0]    _zz_dataOut_payload_0_13558;
  wire       [7:0]    _zz_dataOut_payload_0_13559;
  wire                _zz_dataOut_payload_0_13560;
  wire       [7:0]    _zz_dataOut_payload_0_13561;
  wire       [7:0]    _zz_dataOut_payload_0_13562;
  wire                _zz_dataOut_payload_0_13563;
  wire       [7:0]    _zz_dataOut_payload_0_13564;
  wire       [7:0]    _zz_dataOut_payload_0_13565;
  wire                _zz_dataOut_payload_0_13566;
  wire       [7:0]    _zz_dataOut_payload_0_13567;
  wire       [7:0]    _zz_dataOut_payload_0_13568;
  wire                _zz_dataOut_payload_0_13569;
  wire       [7:0]    _zz_dataOut_payload_0_13570;
  wire       [7:0]    _zz_dataOut_payload_0_13571;
  wire                _zz_dataOut_payload_0_13572;
  wire       [7:0]    _zz_dataOut_payload_0_13573;
  wire       [7:0]    _zz_dataOut_payload_0_13574;
  wire                _zz_dataOut_payload_0_13575;
  wire       [7:0]    _zz_dataOut_payload_0_13576;
  wire       [7:0]    _zz_dataOut_payload_0_13577;
  wire                _zz_dataOut_payload_0_13578;
  wire                _zz_dataOut_payload_0_13579;
  reg        [7:0]    _zz_dataOut_payload_0_13580;
  reg        [7:0]    _zz_dataOut_payload_0_13581;
  reg        [7:0]    _zz_dataOut_payload_0_13582;
  reg        [7:0]    _zz_dataOut_payload_0_13583;
  wire                _zz_dataOut_payload_0_13584;
  wire       [7:0]    _zz_dataOut_payload_0_13585;
  wire       [7:0]    _zz_dataOut_payload_0_13586;
  wire                _zz_dataOut_payload_0_13587;
  wire       [7:0]    _zz_dataOut_payload_0_13588;
  wire       [7:0]    _zz_dataOut_payload_0_13589;
  wire                _zz_dataOut_payload_0_13590;
  wire                _zz_dataOut_payload_0_13591;
  reg        [7:0]    _zz_dataOut_payload_0_13592;
  reg        [7:0]    _zz_dataOut_payload_0_13593;
  reg        [7:0]    _zz_dataOut_payload_0_13594;
  reg        [7:0]    _zz_dataOut_payload_0_13595;
  reg        [7:0]    _zz_dataOut_payload_0_13596;
  reg        [7:0]    _zz_dataOut_payload_0_13597;
  reg        [7:0]    _zz_dataOut_payload_0_13598;
  reg        [7:0]    _zz_dataOut_payload_0_13599;
  reg        [7:0]    _zz_dataOut_payload_0_13600;
  reg        [7:0]    _zz_dataOut_payload_0_13601;
  reg        [7:0]    _zz_dataOut_payload_0_13602;
  reg        [7:0]    _zz_dataOut_payload_0_13603;
  wire                _zz_dataOut_payload_0_13604;
  wire       [7:0]    _zz_dataOut_payload_0_13605;
  wire       [7:0]    _zz_dataOut_payload_0_13606;
  wire                _zz_dataOut_payload_0_13607;
  wire       [7:0]    _zz_dataOut_payload_0_13608;
  wire       [7:0]    _zz_dataOut_payload_0_13609;
  wire                _zz_dataOut_payload_0_13610;
  wire       [7:0]    _zz_dataOut_payload_0_13611;
  wire       [7:0]    _zz_dataOut_payload_0_13612;
  wire                _zz_dataOut_payload_0_13613;
  wire       [7:0]    _zz_dataOut_payload_0_13614;
  wire       [7:0]    _zz_dataOut_payload_0_13615;
  wire                _zz_dataOut_payload_0_13616;
  wire       [7:0]    _zz_dataOut_payload_0_13617;
  wire       [7:0]    _zz_dataOut_payload_0_13618;
  wire                _zz_dataOut_payload_0_13619;
  wire       [7:0]    _zz_dataOut_payload_0_13620;
  wire       [7:0]    _zz_dataOut_payload_0_13621;
  wire                _zz_dataOut_payload_0_13622;
  wire                _zz_dataOut_payload_0_13623;
  reg        [7:0]    _zz_dataOut_payload_0_13624;
  reg        [7:0]    _zz_dataOut_payload_0_13625;
  reg        [7:0]    _zz_dataOut_payload_0_13626;
  reg        [7:0]    _zz_dataOut_payload_0_13627;
  wire                _zz_dataOut_payload_0_13628;
  wire       [7:0]    _zz_dataOut_payload_0_13629;
  wire       [7:0]    _zz_dataOut_payload_0_13630;
  wire                _zz_dataOut_payload_0_13631;
  wire       [7:0]    _zz_dataOut_payload_0_13632;
  wire       [7:0]    _zz_dataOut_payload_0_13633;
  wire                _zz_dataOut_payload_0_13634;
  wire                _zz_dataOut_payload_0_13635;
  reg        [7:0]    _zz_dataOut_payload_0_13636;
  reg        [7:0]    _zz_dataOut_payload_0_13637;
  reg        [7:0]    _zz_dataOut_payload_0_13638;
  reg        [7:0]    _zz_dataOut_payload_0_13639;
  reg        [7:0]    _zz_dataOut_payload_0_13640;
  reg        [7:0]    _zz_dataOut_payload_0_13641;
  reg        [7:0]    _zz_dataOut_payload_0_13642;
  reg        [7:0]    _zz_dataOut_payload_0_13643;
  reg        [7:0]    _zz_dataOut_payload_0_13644;
  reg        [7:0]    _zz_dataOut_payload_0_13645;
  reg        [7:0]    _zz_dataOut_payload_0_13646;
  reg        [7:0]    _zz_dataOut_payload_0_13647;
  reg        [7:0]    _zz_dataOut_payload_0_13648;
  reg        [7:0]    _zz_dataOut_payload_0_13649;
  reg        [7:0]    _zz_dataOut_payload_0_13650;
  reg        [7:0]    _zz_dataOut_payload_0_13651;
  reg        [7:0]    _zz_dataOut_payload_0_13652;
  reg        [7:0]    _zz_dataOut_payload_0_13653;
  reg        [7:0]    _zz_dataOut_payload_0_13654;
  reg        [7:0]    _zz_dataOut_payload_0_13655;
  reg        [7:0]    _zz_dataOut_payload_0_13656;
  reg        [7:0]    _zz_dataOut_payload_0_13657;
  reg        [7:0]    _zz_dataOut_payload_0_13658;
  reg        [7:0]    _zz_dataOut_payload_0_13659;
  reg        [7:0]    _zz_dataOut_payload_0_13660;
  reg        [7:0]    _zz_dataOut_payload_0_13661;
  reg        [7:0]    _zz_dataOut_payload_0_13662;
  reg        [7:0]    _zz_dataOut_payload_0_13663;
  reg        [7:0]    _zz_dataOut_payload_0_13664;
  reg        [7:0]    _zz_dataOut_payload_0_13665;
  reg        [7:0]    _zz_dataOut_payload_0_13666;
  reg        [7:0]    _zz_dataOut_payload_0_13667;
  reg        [7:0]    _zz_dataOut_payload_0_13668;
  reg        [7:0]    _zz_dataOut_payload_0_13669;
  reg        [7:0]    _zz_dataOut_payload_0_13670;
  reg        [7:0]    _zz_dataOut_payload_0_13671;
  reg        [7:0]    _zz_dataOut_payload_0_13672;
  reg        [7:0]    _zz_dataOut_payload_0_13673;
  reg        [7:0]    _zz_dataOut_payload_0_13674;
  reg        [7:0]    _zz_dataOut_payload_0_13675;
  reg        [7:0]    _zz_dataOut_payload_0_13676;
  reg        [7:0]    _zz_dataOut_payload_0_13677;
  reg        [7:0]    _zz_dataOut_payload_0_13678;
  reg        [7:0]    _zz_dataOut_payload_0_13679;
  reg        [7:0]    _zz_dataOut_payload_0_13680;
  reg        [7:0]    _zz_dataOut_payload_0_13681;
  reg        [7:0]    _zz_dataOut_payload_0_13682;
  reg        [7:0]    _zz_dataOut_payload_0_13683;
  reg        [7:0]    _zz_dataOut_payload_0_13684;
  reg        [7:0]    _zz_dataOut_payload_0_13685;
  reg        [7:0]    _zz_dataOut_payload_0_13686;
  reg        [7:0]    _zz_dataOut_payload_0_13687;
  reg        [7:0]    _zz_dataOut_payload_0_13688;
  reg        [7:0]    _zz_dataOut_payload_0_13689;
  reg        [7:0]    _zz_dataOut_payload_0_13690;
  reg        [7:0]    _zz_dataOut_payload_0_13691;
  reg        [7:0]    _zz_dataOut_payload_0_13692;
  reg        [7:0]    _zz_dataOut_payload_0_13693;
  reg        [7:0]    _zz_dataOut_payload_0_13694;
  reg        [7:0]    _zz_dataOut_payload_0_13695;
  reg        [7:0]    _zz_dataOut_payload_0_13696;
  reg        [7:0]    _zz_dataOut_payload_0_13697;
  reg        [7:0]    _zz_dataOut_payload_0_13698;
  reg        [7:0]    _zz_dataOut_payload_0_13699;
  reg        [7:0]    _zz_dataOut_payload_0_13700;
  reg        [7:0]    _zz_dataOut_payload_0_13701;
  reg        [7:0]    _zz_dataOut_payload_0_13702;
  reg        [7:0]    _zz_dataOut_payload_0_13703;
  reg        [7:0]    _zz_dataOut_payload_0_13704;
  reg        [7:0]    _zz_dataOut_payload_0_13705;
  reg        [7:0]    _zz_dataOut_payload_0_13706;
  reg        [7:0]    _zz_dataOut_payload_0_13707;
  reg        [7:0]    _zz_dataOut_payload_0_13708;
  reg        [7:0]    _zz_dataOut_payload_0_13709;
  reg        [7:0]    _zz_dataOut_payload_0_13710;
  reg        [7:0]    _zz_dataOut_payload_0_13711;
  reg        [7:0]    _zz_dataOut_payload_0_13712;
  reg        [7:0]    _zz_dataOut_payload_0_13713;
  reg        [7:0]    _zz_dataOut_payload_0_13714;
  reg        [7:0]    _zz_dataOut_payload_0_13715;
  reg        [7:0]    _zz_dataOut_payload_0_13716;
  reg        [7:0]    _zz_dataOut_payload_0_13717;
  reg        [7:0]    _zz_dataOut_payload_0_13718;
  reg        [7:0]    _zz_dataOut_payload_0_13719;
  reg        [7:0]    _zz_dataOut_payload_0_13720;
  reg        [7:0]    _zz_dataOut_payload_0_13721;
  reg        [7:0]    _zz_dataOut_payload_0_13722;
  reg        [7:0]    _zz_dataOut_payload_0_13723;
  reg        [7:0]    _zz_dataOut_payload_0_13724;
  reg        [7:0]    _zz_dataOut_payload_0_13725;
  reg        [7:0]    _zz_dataOut_payload_0_13726;
  reg        [7:0]    _zz_dataOut_payload_0_13727;
  reg        [7:0]    _zz_dataOut_payload_0_13728;
  reg        [7:0]    _zz_dataOut_payload_0_13729;
  reg        [7:0]    _zz_dataOut_payload_0_13730;
  reg        [7:0]    _zz_dataOut_payload_0_13731;
  reg        [7:0]    _zz_dataOut_payload_0_13732;
  reg        [7:0]    _zz_dataOut_payload_0_13733;
  reg        [7:0]    _zz_dataOut_payload_0_13734;
  reg        [7:0]    _zz_dataOut_payload_0_13735;
  reg        [7:0]    _zz_dataOut_payload_0_13736;
  reg        [7:0]    _zz_dataOut_payload_0_13737;
  reg        [7:0]    _zz_dataOut_payload_0_13738;
  reg        [7:0]    _zz_dataOut_payload_0_13739;
  reg        [7:0]    _zz_dataOut_payload_0_13740;
  reg        [7:0]    _zz_dataOut_payload_0_13741;
  reg        [7:0]    _zz_dataOut_payload_0_13742;
  reg        [7:0]    _zz_dataOut_payload_0_13743;
  reg        [7:0]    _zz_dataOut_payload_0_13744;
  reg        [7:0]    _zz_dataOut_payload_0_13745;
  reg        [7:0]    _zz_dataOut_payload_0_13746;
  reg        [7:0]    _zz_dataOut_payload_0_13747;
  reg        [7:0]    _zz_dataOut_payload_0_13748;
  reg        [7:0]    _zz_dataOut_payload_0_13749;
  reg        [7:0]    _zz_dataOut_payload_0_13750;
  reg        [7:0]    _zz_dataOut_payload_0_13751;
  reg        [7:0]    _zz_dataOut_payload_0_13752;
  reg        [7:0]    _zz_dataOut_payload_0_13753;
  reg        [7:0]    _zz_dataOut_payload_0_13754;
  reg        [7:0]    _zz_dataOut_payload_0_13755;
  reg        [7:0]    _zz_dataOut_payload_0_13756;
  reg        [7:0]    _zz_dataOut_payload_0_13757;
  reg        [7:0]    _zz_dataOut_payload_0_13758;
  reg        [7:0]    _zz_dataOut_payload_0_13759;
  reg        [7:0]    _zz_dataOut_payload_0_13760;
  reg        [7:0]    _zz_dataOut_payload_0_13761;
  reg        [7:0]    _zz_dataOut_payload_0_13762;
  reg        [7:0]    _zz_dataOut_payload_0_13763;
  reg        [7:0]    _zz_dataOut_payload_0_13764;
  reg        [7:0]    _zz_dataOut_payload_0_13765;
  reg        [7:0]    _zz_dataOut_payload_0_13766;
  reg        [7:0]    _zz_dataOut_payload_0_13767;
  reg        [7:0]    _zz_dataOut_payload_0_13768;
  reg        [7:0]    _zz_dataOut_payload_0_13769;
  reg        [7:0]    _zz_dataOut_payload_0_13770;
  reg        [7:0]    _zz_dataOut_payload_0_13771;
  reg        [7:0]    _zz_dataOut_payload_0_13772;
  reg        [7:0]    _zz_dataOut_payload_0_13773;
  reg        [7:0]    _zz_dataOut_payload_0_13774;
  reg        [7:0]    _zz_dataOut_payload_0_13775;
  reg        [7:0]    _zz_dataOut_payload_0_13776;
  reg        [7:0]    _zz_dataOut_payload_0_13777;
  reg        [7:0]    _zz_dataOut_payload_0_13778;
  reg        [7:0]    _zz_dataOut_payload_0_13779;
  reg        [7:0]    _zz_dataOut_payload_0_13780;
  reg        [7:0]    _zz_dataOut_payload_0_13781;
  reg        [7:0]    _zz_dataOut_payload_0_13782;
  reg        [7:0]    _zz_dataOut_payload_0_13783;
  reg        [7:0]    _zz_dataOut_payload_0_13784;
  reg        [7:0]    _zz_dataOut_payload_0_13785;
  reg        [7:0]    _zz_dataOut_payload_0_13786;
  reg        [7:0]    _zz_dataOut_payload_0_13787;
  reg        [7:0]    _zz_dataOut_payload_0_13788;
  reg        [7:0]    _zz_dataOut_payload_0_13789;
  reg        [7:0]    _zz_dataOut_payload_0_13790;
  reg        [7:0]    _zz_dataOut_payload_0_13791;
  reg        [7:0]    _zz_dataOut_payload_0_13792;
  reg        [7:0]    _zz_dataOut_payload_0_13793;
  reg        [7:0]    _zz_dataOut_payload_0_13794;
  reg        [7:0]    _zz_dataOut_payload_0_13795;
  reg        [7:0]    _zz_dataOut_payload_0_13796;
  reg        [7:0]    _zz_dataOut_payload_0_13797;
  reg        [7:0]    _zz_dataOut_payload_0_13798;
  reg        [7:0]    _zz_dataOut_payload_0_13799;
  reg        [7:0]    _zz_dataOut_payload_0_13800;
  reg        [7:0]    _zz_dataOut_payload_0_13801;
  reg        [7:0]    _zz_dataOut_payload_0_13802;
  reg        [7:0]    _zz_dataOut_payload_0_13803;
  reg        [7:0]    _zz_dataOut_payload_0_13804;
  reg        [7:0]    _zz_dataOut_payload_0_13805;
  reg        [7:0]    _zz_dataOut_payload_0_13806;
  reg        [7:0]    _zz_dataOut_payload_0_13807;
  reg        [7:0]    _zz_dataOut_payload_0_13808;
  reg        [7:0]    _zz_dataOut_payload_0_13809;
  reg        [7:0]    _zz_dataOut_payload_0_13810;
  reg        [7:0]    _zz_dataOut_payload_0_13811;
  reg        [7:0]    _zz_dataOut_payload_0_13812;
  reg        [7:0]    _zz_dataOut_payload_0_13813;
  reg        [7:0]    _zz_dataOut_payload_0_13814;
  reg        [7:0]    _zz_dataOut_payload_0_13815;
  reg        [7:0]    _zz_dataOut_payload_0_13816;
  reg        [7:0]    _zz_dataOut_payload_0_13817;
  reg        [7:0]    _zz_dataOut_payload_0_13818;
  reg        [7:0]    _zz_dataOut_payload_0_13819;
  reg        [7:0]    _zz_dataOut_payload_0_13820;
  reg        [7:0]    _zz_dataOut_payload_0_13821;
  reg        [7:0]    _zz_dataOut_payload_0_13822;
  reg        [7:0]    _zz_dataOut_payload_0_13823;
  reg        [7:0]    _zz_dataOut_payload_0_13824;
  reg        [7:0]    _zz_dataOut_payload_0_13825;
  reg        [7:0]    _zz_dataOut_payload_0_13826;
  reg        [7:0]    _zz_dataOut_payload_0_13827;
  reg        [7:0]    _zz_dataOut_payload_0_13828;
  reg        [7:0]    _zz_dataOut_payload_0_13829;
  reg        [7:0]    _zz_dataOut_payload_0_13830;
  reg        [7:0]    _zz_dataOut_payload_0_13831;
  reg        [7:0]    _zz_dataOut_payload_0_13832;
  reg        [7:0]    _zz_dataOut_payload_0_13833;
  reg        [7:0]    _zz_dataOut_payload_0_13834;
  reg        [7:0]    _zz_dataOut_payload_0_13835;
  reg        [7:0]    _zz_dataOut_payload_0_13836;
  reg        [7:0]    _zz_dataOut_payload_0_13837;
  reg        [7:0]    _zz_dataOut_payload_0_13838;
  reg        [7:0]    _zz_dataOut_payload_0_13839;
  reg        [7:0]    _zz_dataOut_payload_0_13840;
  reg        [7:0]    _zz_dataOut_payload_0_13841;
  reg        [7:0]    _zz_dataOut_payload_0_13842;
  reg        [7:0]    _zz_dataOut_payload_0_13843;
  reg        [7:0]    _zz_dataOut_payload_0_13844;
  reg        [7:0]    _zz_dataOut_payload_0_13845;
  reg        [7:0]    _zz_dataOut_payload_0_13846;
  reg        [7:0]    _zz_dataOut_payload_0_13847;
  reg        [7:0]    _zz_dataOut_payload_0_13848;
  reg        [7:0]    _zz_dataOut_payload_0_13849;
  reg        [7:0]    _zz_dataOut_payload_0_13850;
  reg        [7:0]    _zz_dataOut_payload_0_13851;
  reg        [7:0]    _zz_dataOut_payload_0_13852;
  reg        [7:0]    _zz_dataOut_payload_0_13853;
  reg        [7:0]    _zz_dataOut_payload_0_13854;
  reg        [7:0]    _zz_dataOut_payload_0_13855;
  reg        [7:0]    _zz_dataOut_payload_0_13856;
  reg        [7:0]    _zz_dataOut_payload_0_13857;
  reg        [7:0]    _zz_dataOut_payload_0_13858;
  reg        [7:0]    _zz_dataOut_payload_0_13859;
  reg        [7:0]    _zz_dataOut_payload_0_13860;
  reg        [7:0]    _zz_dataOut_payload_0_13861;
  reg        [7:0]    _zz_dataOut_payload_0_13862;
  reg        [7:0]    _zz_dataOut_payload_0_13863;
  reg        [7:0]    _zz_dataOut_payload_0_13864;
  reg        [7:0]    _zz_dataOut_payload_0_13865;
  reg        [7:0]    _zz_dataOut_payload_0_13866;
  reg        [7:0]    _zz_dataOut_payload_0_13867;
  reg        [7:0]    _zz_dataOut_payload_0_13868;
  reg        [7:0]    _zz_dataOut_payload_0_13869;
  reg        [7:0]    _zz_dataOut_payload_0_13870;
  reg        [7:0]    _zz_dataOut_payload_0_13871;
  reg        [7:0]    _zz_dataOut_payload_0_13872;
  reg        [7:0]    _zz_dataOut_payload_0_13873;
  reg        [7:0]    _zz_dataOut_payload_0_13874;
  reg        [7:0]    _zz_dataOut_payload_0_13875;
  reg        [7:0]    _zz_dataOut_payload_0_13876;
  reg        [7:0]    _zz_dataOut_payload_0_13877;
  reg        [7:0]    _zz_dataOut_payload_0_13878;
  reg        [7:0]    _zz_dataOut_payload_0_13879;
  reg        [7:0]    _zz_dataOut_payload_0_13880;
  reg        [7:0]    _zz_dataOut_payload_0_13881;
  reg        [7:0]    _zz_dataOut_payload_0_13882;
  reg        [7:0]    _zz_dataOut_payload_0_13883;
  reg        [7:0]    _zz_dataOut_payload_0_13884;
  reg        [7:0]    _zz_dataOut_payload_0_13885;
  reg        [7:0]    _zz_dataOut_payload_0_13886;
  reg        [7:0]    _zz_dataOut_payload_0_13887;
  wire                _zz_dataOut_payload_0_13888;
  wire       [7:0]    _zz_dataOut_payload_0_13889;
  wire       [7:0]    _zz_dataOut_payload_0_13890;
  wire                _zz_dataOut_payload_0_13891;
  wire       [7:0]    _zz_dataOut_payload_0_13892;
  wire       [7:0]    _zz_dataOut_payload_0_13893;
  wire                _zz_dataOut_payload_0_13894;
  wire       [7:0]    _zz_dataOut_payload_0_13895;
  wire       [7:0]    _zz_dataOut_payload_0_13896;
  wire                _zz_dataOut_payload_0_13897;
  wire       [7:0]    _zz_dataOut_payload_0_13898;
  wire       [7:0]    _zz_dataOut_payload_0_13899;
  wire                _zz_dataOut_payload_0_13900;
  wire       [7:0]    _zz_dataOut_payload_0_13901;
  wire       [7:0]    _zz_dataOut_payload_0_13902;
  wire                _zz_dataOut_payload_0_13903;
  wire       [7:0]    _zz_dataOut_payload_0_13904;
  wire       [7:0]    _zz_dataOut_payload_0_13905;
  wire                _zz_dataOut_payload_0_13906;
  wire       [7:0]    _zz_dataOut_payload_0_13907;
  wire       [7:0]    _zz_dataOut_payload_0_13908;
  wire                _zz_dataOut_payload_0_13909;
  wire       [7:0]    _zz_dataOut_payload_0_13910;
  wire       [7:0]    _zz_dataOut_payload_0_13911;
  wire                _zz_dataOut_payload_0_13912;
  wire       [7:0]    _zz_dataOut_payload_0_13913;
  wire       [7:0]    _zz_dataOut_payload_0_13914;
  wire                _zz_dataOut_payload_0_13915;
  wire       [7:0]    _zz_dataOut_payload_0_13916;
  wire       [7:0]    _zz_dataOut_payload_0_13917;
  wire                _zz_dataOut_payload_0_13918;
  wire       [7:0]    _zz_dataOut_payload_0_13919;
  wire       [7:0]    _zz_dataOut_payload_0_13920;
  wire                _zz_dataOut_payload_0_13921;
  wire       [7:0]    _zz_dataOut_payload_0_13922;
  wire       [7:0]    _zz_dataOut_payload_0_13923;
  wire                _zz_dataOut_payload_0_13924;
  wire       [7:0]    _zz_dataOut_payload_0_13925;
  wire       [7:0]    _zz_dataOut_payload_0_13926;
  wire                _zz_dataOut_payload_0_13927;
  wire       [7:0]    _zz_dataOut_payload_0_13928;
  wire       [7:0]    _zz_dataOut_payload_0_13929;
  wire                _zz_dataOut_payload_0_13930;
  wire       [7:0]    _zz_dataOut_payload_0_13931;
  wire       [7:0]    _zz_dataOut_payload_0_13932;
  wire                _zz_dataOut_payload_0_13933;
  wire       [7:0]    _zz_dataOut_payload_0_13934;
  wire       [7:0]    _zz_dataOut_payload_0_13935;
  wire                _zz_dataOut_payload_0_13936;
  wire       [7:0]    _zz_dataOut_payload_0_13937;
  wire       [7:0]    _zz_dataOut_payload_0_13938;
  wire                _zz_dataOut_payload_0_13939;
  wire       [7:0]    _zz_dataOut_payload_0_13940;
  wire       [7:0]    _zz_dataOut_payload_0_13941;
  wire                _zz_dataOut_payload_0_13942;
  wire       [7:0]    _zz_dataOut_payload_0_13943;
  wire       [7:0]    _zz_dataOut_payload_0_13944;
  wire                _zz_dataOut_payload_0_13945;
  wire       [7:0]    _zz_dataOut_payload_0_13946;
  wire       [7:0]    _zz_dataOut_payload_0_13947;
  wire                _zz_dataOut_payload_0_13948;
  wire       [7:0]    _zz_dataOut_payload_0_13949;
  wire       [7:0]    _zz_dataOut_payload_0_13950;
  wire                _zz_dataOut_payload_0_13951;
  wire       [7:0]    _zz_dataOut_payload_0_13952;
  wire       [7:0]    _zz_dataOut_payload_0_13953;
  wire                _zz_dataOut_payload_0_13954;
  wire       [7:0]    _zz_dataOut_payload_0_13955;
  wire       [7:0]    _zz_dataOut_payload_0_13956;
  wire                _zz_dataOut_payload_0_13957;
  wire       [7:0]    _zz_dataOut_payload_0_13958;
  wire       [7:0]    _zz_dataOut_payload_0_13959;
  wire                _zz_dataOut_payload_0_13960;
  wire       [7:0]    _zz_dataOut_payload_0_13961;
  wire       [7:0]    _zz_dataOut_payload_0_13962;
  wire                _zz_dataOut_payload_0_13963;
  wire       [7:0]    _zz_dataOut_payload_0_13964;
  wire       [7:0]    _zz_dataOut_payload_0_13965;
  wire                _zz_dataOut_payload_0_13966;
  wire       [7:0]    _zz_dataOut_payload_0_13967;
  wire       [7:0]    _zz_dataOut_payload_0_13968;
  wire                _zz_dataOut_payload_0_13969;
  wire       [7:0]    _zz_dataOut_payload_0_13970;
  wire       [7:0]    _zz_dataOut_payload_0_13971;
  wire                _zz_dataOut_payload_0_13972;
  wire       [7:0]    _zz_dataOut_payload_0_13973;
  wire       [7:0]    _zz_dataOut_payload_0_13974;
  wire                _zz_dataOut_payload_0_13975;
  wire       [7:0]    _zz_dataOut_payload_0_13976;
  wire       [7:0]    _zz_dataOut_payload_0_13977;
  wire                _zz_dataOut_payload_0_13978;
  wire       [7:0]    _zz_dataOut_payload_0_13979;
  wire       [7:0]    _zz_dataOut_payload_0_13980;
  wire                _zz_dataOut_payload_0_13981;
  wire       [7:0]    _zz_dataOut_payload_0_13982;
  wire       [7:0]    _zz_dataOut_payload_0_13983;
  wire                _zz_dataOut_payload_0_13984;
  wire       [7:0]    _zz_dataOut_payload_0_13985;
  wire       [7:0]    _zz_dataOut_payload_0_13986;
  wire                _zz_dataOut_payload_0_13987;
  wire       [7:0]    _zz_dataOut_payload_0_13988;
  wire       [7:0]    _zz_dataOut_payload_0_13989;
  wire                _zz_dataOut_payload_0_13990;
  wire       [7:0]    _zz_dataOut_payload_0_13991;
  wire       [7:0]    _zz_dataOut_payload_0_13992;
  wire                _zz_dataOut_payload_0_13993;
  wire       [7:0]    _zz_dataOut_payload_0_13994;
  wire       [7:0]    _zz_dataOut_payload_0_13995;
  wire                _zz_dataOut_payload_0_13996;
  wire       [7:0]    _zz_dataOut_payload_0_13997;
  wire       [7:0]    _zz_dataOut_payload_0_13998;
  wire                _zz_dataOut_payload_0_13999;
  wire       [7:0]    _zz_dataOut_payload_0_14000;
  wire       [7:0]    _zz_dataOut_payload_0_14001;
  wire                _zz_dataOut_payload_0_14002;
  wire       [7:0]    _zz_dataOut_payload_0_14003;
  wire       [7:0]    _zz_dataOut_payload_0_14004;
  wire                _zz_dataOut_payload_0_14005;
  wire       [7:0]    _zz_dataOut_payload_0_14006;
  wire       [7:0]    _zz_dataOut_payload_0_14007;
  wire                _zz_dataOut_payload_0_14008;
  wire       [7:0]    _zz_dataOut_payload_0_14009;
  wire       [7:0]    _zz_dataOut_payload_0_14010;
  wire                _zz_dataOut_payload_0_14011;
  wire       [7:0]    _zz_dataOut_payload_0_14012;
  wire       [7:0]    _zz_dataOut_payload_0_14013;
  wire                _zz_dataOut_payload_0_14014;
  wire       [7:0]    _zz_dataOut_payload_0_14015;
  wire       [7:0]    _zz_dataOut_payload_0_14016;
  wire                _zz_dataOut_payload_0_14017;
  wire       [7:0]    _zz_dataOut_payload_0_14018;
  wire       [7:0]    _zz_dataOut_payload_0_14019;
  wire                _zz_dataOut_payload_0_14020;
  wire       [7:0]    _zz_dataOut_payload_0_14021;
  wire       [7:0]    _zz_dataOut_payload_0_14022;
  wire                _zz_dataOut_payload_0_14023;
  wire       [7:0]    _zz_dataOut_payload_0_14024;
  wire       [7:0]    _zz_dataOut_payload_0_14025;
  wire                _zz_dataOut_payload_0_14026;
  wire       [7:0]    _zz_dataOut_payload_0_14027;
  wire       [7:0]    _zz_dataOut_payload_0_14028;
  wire                _zz_dataOut_payload_0_14029;
  wire       [7:0]    _zz_dataOut_payload_0_14030;
  wire       [7:0]    _zz_dataOut_payload_0_14031;
  wire                _zz_dataOut_payload_0_14032;
  wire       [7:0]    _zz_dataOut_payload_0_14033;
  wire       [7:0]    _zz_dataOut_payload_0_14034;
  wire                _zz_dataOut_payload_0_14035;
  wire       [7:0]    _zz_dataOut_payload_0_14036;
  wire       [7:0]    _zz_dataOut_payload_0_14037;
  wire                _zz_dataOut_payload_0_14038;
  wire       [7:0]    _zz_dataOut_payload_0_14039;
  wire       [7:0]    _zz_dataOut_payload_0_14040;
  wire                _zz_dataOut_payload_0_14041;
  wire       [7:0]    _zz_dataOut_payload_0_14042;
  wire       [7:0]    _zz_dataOut_payload_0_14043;
  wire                _zz_dataOut_payload_0_14044;
  wire       [7:0]    _zz_dataOut_payload_0_14045;
  wire       [7:0]    _zz_dataOut_payload_0_14046;
  wire                _zz_dataOut_payload_0_14047;
  wire       [7:0]    _zz_dataOut_payload_0_14048;
  wire       [7:0]    _zz_dataOut_payload_0_14049;
  wire                _zz_dataOut_payload_0_14050;
  wire       [7:0]    _zz_dataOut_payload_0_14051;
  wire       [7:0]    _zz_dataOut_payload_0_14052;
  wire                _zz_dataOut_payload_0_14053;
  wire       [7:0]    _zz_dataOut_payload_0_14054;
  wire       [7:0]    _zz_dataOut_payload_0_14055;
  wire                _zz_dataOut_payload_0_14056;
  wire       [7:0]    _zz_dataOut_payload_0_14057;
  wire       [7:0]    _zz_dataOut_payload_0_14058;
  wire                _zz_dataOut_payload_0_14059;
  wire       [7:0]    _zz_dataOut_payload_0_14060;
  wire       [7:0]    _zz_dataOut_payload_0_14061;
  wire                _zz_dataOut_payload_0_14062;
  wire       [7:0]    _zz_dataOut_payload_0_14063;
  wire       [7:0]    _zz_dataOut_payload_0_14064;
  wire                _zz_dataOut_payload_0_14065;
  wire       [7:0]    _zz_dataOut_payload_0_14066;
  wire       [7:0]    _zz_dataOut_payload_0_14067;
  wire                _zz_dataOut_payload_0_14068;
  wire       [7:0]    _zz_dataOut_payload_0_14069;
  wire       [7:0]    _zz_dataOut_payload_0_14070;
  wire                _zz_dataOut_payload_0_14071;
  wire       [7:0]    _zz_dataOut_payload_0_14072;
  wire       [7:0]    _zz_dataOut_payload_0_14073;
  wire                _zz_dataOut_payload_0_14074;
  wire       [7:0]    _zz_dataOut_payload_0_14075;
  wire       [7:0]    _zz_dataOut_payload_0_14076;
  wire                _zz_dataOut_payload_0_14077;
  wire       [7:0]    _zz_dataOut_payload_0_14078;
  wire       [7:0]    _zz_dataOut_payload_0_14079;
  wire                _zz_dataOut_payload_0_14080;
  wire       [7:0]    _zz_dataOut_payload_0_14081;
  wire       [7:0]    _zz_dataOut_payload_0_14082;
  wire                _zz_dataOut_payload_0_14083;
  wire       [7:0]    _zz_dataOut_payload_0_14084;
  wire       [7:0]    _zz_dataOut_payload_0_14085;
  wire                _zz_dataOut_payload_0_14086;
  wire       [7:0]    _zz_dataOut_payload_0_14087;
  wire       [7:0]    _zz_dataOut_payload_0_14088;
  wire                _zz_dataOut_payload_0_14089;
  wire       [7:0]    _zz_dataOut_payload_0_14090;
  wire       [7:0]    _zz_dataOut_payload_0_14091;
  wire                _zz_dataOut_payload_0_14092;
  wire       [7:0]    _zz_dataOut_payload_0_14093;
  wire       [7:0]    _zz_dataOut_payload_0_14094;
  wire                _zz_dataOut_payload_0_14095;
  wire       [7:0]    _zz_dataOut_payload_0_14096;
  wire       [7:0]    _zz_dataOut_payload_0_14097;
  wire                _zz_dataOut_payload_0_14098;
  wire       [7:0]    _zz_dataOut_payload_0_14099;
  wire       [7:0]    _zz_dataOut_payload_0_14100;
  wire                _zz_dataOut_payload_0_14101;
  wire       [7:0]    _zz_dataOut_payload_0_14102;
  wire       [7:0]    _zz_dataOut_payload_0_14103;
  wire                _zz_dataOut_payload_0_14104;
  wire       [7:0]    _zz_dataOut_payload_0_14105;
  wire       [7:0]    _zz_dataOut_payload_0_14106;
  wire                _zz_dataOut_payload_0_14107;
  wire       [7:0]    _zz_dataOut_payload_0_14108;
  wire       [7:0]    _zz_dataOut_payload_0_14109;
  wire                _zz_dataOut_payload_0_14110;
  wire       [7:0]    _zz_dataOut_payload_0_14111;
  wire       [7:0]    _zz_dataOut_payload_0_14112;
  wire                _zz_dataOut_payload_0_14113;
  wire       [7:0]    _zz_dataOut_payload_0_14114;
  wire       [7:0]    _zz_dataOut_payload_0_14115;
  wire                _zz_dataOut_payload_0_14116;
  wire       [7:0]    _zz_dataOut_payload_0_14117;
  wire       [7:0]    _zz_dataOut_payload_0_14118;
  wire                _zz_dataOut_payload_0_14119;
  wire       [7:0]    _zz_dataOut_payload_0_14120;
  wire       [7:0]    _zz_dataOut_payload_0_14121;
  wire                _zz_dataOut_payload_0_14122;
  wire       [7:0]    _zz_dataOut_payload_0_14123;
  wire       [7:0]    _zz_dataOut_payload_0_14124;
  wire                _zz_dataOut_payload_0_14125;
  wire       [7:0]    _zz_dataOut_payload_0_14126;
  wire       [7:0]    _zz_dataOut_payload_0_14127;
  wire                _zz_dataOut_payload_0_14128;
  wire       [7:0]    _zz_dataOut_payload_0_14129;
  wire       [7:0]    _zz_dataOut_payload_0_14130;
  wire                _zz_dataOut_payload_0_14131;
  wire       [7:0]    _zz_dataOut_payload_0_14132;
  wire       [7:0]    _zz_dataOut_payload_0_14133;
  wire                _zz_dataOut_payload_0_14134;
  wire       [7:0]    _zz_dataOut_payload_0_14135;
  wire       [7:0]    _zz_dataOut_payload_0_14136;
  wire                _zz_dataOut_payload_0_14137;
  wire       [7:0]    _zz_dataOut_payload_0_14138;
  wire       [7:0]    _zz_dataOut_payload_0_14139;
  wire                _zz_dataOut_payload_0_14140;
  wire       [7:0]    _zz_dataOut_payload_0_14141;
  wire       [7:0]    _zz_dataOut_payload_0_14142;
  wire                _zz_dataOut_payload_0_14143;
  wire       [7:0]    _zz_dataOut_payload_0_14144;
  wire       [7:0]    _zz_dataOut_payload_0_14145;
  wire                _zz_dataOut_payload_0_14146;
  wire       [7:0]    _zz_dataOut_payload_0_14147;
  wire       [7:0]    _zz_dataOut_payload_0_14148;
  wire                _zz_dataOut_payload_0_14149;
  wire       [7:0]    _zz_dataOut_payload_0_14150;
  wire       [7:0]    _zz_dataOut_payload_0_14151;
  wire                _zz_dataOut_payload_0_14152;
  wire       [7:0]    _zz_dataOut_payload_0_14153;
  wire       [7:0]    _zz_dataOut_payload_0_14154;
  wire                _zz_dataOut_payload_0_14155;
  wire       [7:0]    _zz_dataOut_payload_0_14156;
  wire       [7:0]    _zz_dataOut_payload_0_14157;
  wire                _zz_dataOut_payload_0_14158;
  wire       [7:0]    _zz_dataOut_payload_0_14159;
  wire       [7:0]    _zz_dataOut_payload_0_14160;
  wire                _zz_dataOut_payload_0_14161;
  wire       [7:0]    _zz_dataOut_payload_0_14162;
  wire       [7:0]    _zz_dataOut_payload_0_14163;
  wire                _zz_dataOut_payload_0_14164;
  wire       [7:0]    _zz_dataOut_payload_0_14165;
  wire       [7:0]    _zz_dataOut_payload_0_14166;
  wire                _zz_dataOut_payload_0_14167;
  wire       [7:0]    _zz_dataOut_payload_0_14168;
  wire       [7:0]    _zz_dataOut_payload_0_14169;
  wire                _zz_dataOut_payload_0_14170;
  wire       [7:0]    _zz_dataOut_payload_0_14171;
  wire       [7:0]    _zz_dataOut_payload_0_14172;
  wire                _zz_dataOut_payload_0_14173;
  wire       [7:0]    _zz_dataOut_payload_0_14174;
  wire       [7:0]    _zz_dataOut_payload_0_14175;
  wire                _zz_dataOut_payload_0_14176;
  wire       [7:0]    _zz_dataOut_payload_0_14177;
  wire       [7:0]    _zz_dataOut_payload_0_14178;
  wire                _zz_dataOut_payload_0_14179;
  wire       [7:0]    _zz_dataOut_payload_0_14180;
  wire       [7:0]    _zz_dataOut_payload_0_14181;
  wire                _zz_dataOut_payload_0_14182;
  wire       [7:0]    _zz_dataOut_payload_0_14183;
  wire       [7:0]    _zz_dataOut_payload_0_14184;
  wire                _zz_dataOut_payload_0_14185;
  wire       [7:0]    _zz_dataOut_payload_0_14186;
  wire       [7:0]    _zz_dataOut_payload_0_14187;
  wire                _zz_dataOut_payload_0_14188;
  wire       [7:0]    _zz_dataOut_payload_0_14189;
  wire       [7:0]    _zz_dataOut_payload_0_14190;
  wire                _zz_dataOut_payload_0_14191;
  wire       [7:0]    _zz_dataOut_payload_0_14192;
  wire       [7:0]    _zz_dataOut_payload_0_14193;
  wire                _zz_dataOut_payload_0_14194;
  wire       [7:0]    _zz_dataOut_payload_0_14195;
  wire       [7:0]    _zz_dataOut_payload_0_14196;
  wire                _zz_dataOut_payload_0_14197;
  wire       [7:0]    _zz_dataOut_payload_0_14198;
  wire       [7:0]    _zz_dataOut_payload_0_14199;
  wire                _zz_dataOut_payload_0_14200;
  wire       [7:0]    _zz_dataOut_payload_0_14201;
  wire       [7:0]    _zz_dataOut_payload_0_14202;
  wire                _zz_dataOut_payload_0_14203;
  wire       [7:0]    _zz_dataOut_payload_0_14204;
  wire       [7:0]    _zz_dataOut_payload_0_14205;
  wire                _zz_dataOut_payload_0_14206;
  wire       [7:0]    _zz_dataOut_payload_0_14207;
  wire       [7:0]    _zz_dataOut_payload_0_14208;
  wire                _zz_dataOut_payload_0_14209;
  wire       [7:0]    _zz_dataOut_payload_0_14210;
  wire       [7:0]    _zz_dataOut_payload_0_14211;
  wire                _zz_dataOut_payload_0_14212;
  wire       [7:0]    _zz_dataOut_payload_0_14213;
  wire       [7:0]    _zz_dataOut_payload_0_14214;
  wire                _zz_dataOut_payload_0_14215;
  wire       [7:0]    _zz_dataOut_payload_0_14216;
  wire       [7:0]    _zz_dataOut_payload_0_14217;
  wire                _zz_dataOut_payload_0_14218;
  wire       [7:0]    _zz_dataOut_payload_0_14219;
  wire       [7:0]    _zz_dataOut_payload_0_14220;
  wire                _zz_dataOut_payload_0_14221;
  wire       [7:0]    _zz_dataOut_payload_0_14222;
  wire       [7:0]    _zz_dataOut_payload_0_14223;
  wire                _zz_dataOut_payload_0_14224;
  wire       [7:0]    _zz_dataOut_payload_0_14225;
  wire       [7:0]    _zz_dataOut_payload_0_14226;
  wire                _zz_dataOut_payload_0_14227;
  wire       [7:0]    _zz_dataOut_payload_0_14228;
  wire       [7:0]    _zz_dataOut_payload_0_14229;
  wire                _zz_dataOut_payload_0_14230;
  wire       [7:0]    _zz_dataOut_payload_0_14231;
  wire       [7:0]    _zz_dataOut_payload_0_14232;
  wire                _zz_dataOut_payload_0_14233;
  wire       [7:0]    _zz_dataOut_payload_0_14234;
  wire       [7:0]    _zz_dataOut_payload_0_14235;
  wire                _zz_dataOut_payload_0_14236;
  wire       [7:0]    _zz_dataOut_payload_0_14237;
  wire       [7:0]    _zz_dataOut_payload_0_14238;
  wire                _zz_dataOut_payload_0_14239;
  wire       [7:0]    _zz_dataOut_payload_0_14240;
  wire       [7:0]    _zz_dataOut_payload_0_14241;
  wire                _zz_dataOut_payload_0_14242;
  wire       [7:0]    _zz_dataOut_payload_0_14243;
  wire       [7:0]    _zz_dataOut_payload_0_14244;
  wire                _zz_dataOut_payload_0_14245;
  wire       [7:0]    _zz_dataOut_payload_0_14246;
  wire       [7:0]    _zz_dataOut_payload_0_14247;
  wire                _zz_dataOut_payload_0_14248;
  wire       [7:0]    _zz_dataOut_payload_0_14249;
  wire       [7:0]    _zz_dataOut_payload_0_14250;
  wire                _zz_dataOut_payload_0_14251;
  wire       [7:0]    _zz_dataOut_payload_0_14252;
  wire       [7:0]    _zz_dataOut_payload_0_14253;
  wire                _zz_dataOut_payload_0_14254;
  wire       [7:0]    _zz_dataOut_payload_0_14255;
  wire       [7:0]    _zz_dataOut_payload_0_14256;
  wire                _zz_dataOut_payload_0_14257;
  wire       [7:0]    _zz_dataOut_payload_0_14258;
  wire       [7:0]    _zz_dataOut_payload_0_14259;
  wire                _zz_dataOut_payload_0_14260;
  wire       [7:0]    _zz_dataOut_payload_0_14261;
  wire       [7:0]    _zz_dataOut_payload_0_14262;
  wire                _zz_dataOut_payload_0_14263;
  wire       [7:0]    _zz_dataOut_payload_0_14264;
  wire       [7:0]    _zz_dataOut_payload_0_14265;
  wire                _zz_dataOut_payload_0_14266;
  wire                _zz_dataOut_payload_0_14267;
  reg        [7:0]    _zz_dataOut_payload_0_14268;
  reg        [7:0]    _zz_dataOut_payload_0_14269;
  reg        [7:0]    _zz_dataOut_payload_0_14270;
  reg        [7:0]    _zz_dataOut_payload_0_14271;
  wire                _zz_dataOut_payload_0_14272;
  wire       [7:0]    _zz_dataOut_payload_0_14273;
  wire       [7:0]    _zz_dataOut_payload_0_14274;
  wire                _zz_dataOut_payload_0_14275;
  wire       [7:0]    _zz_dataOut_payload_0_14276;
  wire       [7:0]    _zz_dataOut_payload_0_14277;
  wire                _zz_dataOut_payload_0_14278;
  wire                _zz_dataOut_payload_0_14279;
  reg        [7:0]    _zz_dataOut_payload_0_14280;
  reg        [7:0]    _zz_dataOut_payload_0_14281;
  reg        [7:0]    _zz_dataOut_payload_0_14282;
  reg        [7:0]    _zz_dataOut_payload_0_14283;
  reg        [7:0]    _zz_dataOut_payload_0_14284;
  reg        [7:0]    _zz_dataOut_payload_0_14285;
  reg        [7:0]    _zz_dataOut_payload_0_14286;
  reg        [7:0]    _zz_dataOut_payload_0_14287;
  reg        [7:0]    _zz_dataOut_payload_0_14288;
  reg        [7:0]    _zz_dataOut_payload_0_14289;
  reg        [7:0]    _zz_dataOut_payload_0_14290;
  reg        [7:0]    _zz_dataOut_payload_0_14291;
  wire                _zz_dataOut_payload_0_14292;
  wire       [7:0]    _zz_dataOut_payload_0_14293;
  wire       [7:0]    _zz_dataOut_payload_0_14294;
  wire                _zz_dataOut_payload_0_14295;
  wire       [7:0]    _zz_dataOut_payload_0_14296;
  wire       [7:0]    _zz_dataOut_payload_0_14297;
  wire                _zz_dataOut_payload_0_14298;
  wire       [7:0]    _zz_dataOut_payload_0_14299;
  wire       [7:0]    _zz_dataOut_payload_0_14300;
  wire                _zz_dataOut_payload_0_14301;
  wire       [7:0]    _zz_dataOut_payload_0_14302;
  wire       [7:0]    _zz_dataOut_payload_0_14303;
  wire                _zz_dataOut_payload_0_14304;
  wire       [7:0]    _zz_dataOut_payload_0_14305;
  wire       [7:0]    _zz_dataOut_payload_0_14306;
  wire                _zz_dataOut_payload_0_14307;
  wire       [7:0]    _zz_dataOut_payload_0_14308;
  wire       [7:0]    _zz_dataOut_payload_0_14309;
  wire                _zz_dataOut_payload_0_14310;
  wire                _zz_dataOut_payload_0_14311;
  reg        [7:0]    _zz_dataOut_payload_0_14312;
  reg        [7:0]    _zz_dataOut_payload_0_14313;
  reg        [7:0]    _zz_dataOut_payload_0_14314;
  reg        [7:0]    _zz_dataOut_payload_0_14315;
  wire                _zz_dataOut_payload_0_14316;
  wire       [7:0]    _zz_dataOut_payload_0_14317;
  wire       [7:0]    _zz_dataOut_payload_0_14318;
  wire                _zz_dataOut_payload_0_14319;
  wire       [7:0]    _zz_dataOut_payload_0_14320;
  wire       [7:0]    _zz_dataOut_payload_0_14321;
  wire                _zz_dataOut_payload_0_14322;
  wire                _zz_dataOut_payload_0_14323;
  reg        [7:0]    _zz_dataOut_payload_0_14324;
  reg        [7:0]    _zz_dataOut_payload_0_14325;
  reg        [7:0]    _zz_dataOut_payload_0_14326;
  reg        [7:0]    _zz_dataOut_payload_0_14327;
  reg        [7:0]    _zz_dataOut_payload_0_14328;
  reg        [7:0]    _zz_dataOut_payload_0_14329;
  reg        [7:0]    _zz_dataOut_payload_0_14330;
  reg        [7:0]    _zz_dataOut_payload_0_14331;
  reg        [7:0]    _zz_dataOut_payload_0_14332;
  reg        [7:0]    _zz_dataOut_payload_0_14333;
  reg        [7:0]    _zz_dataOut_payload_0_14334;
  reg        [7:0]    _zz_dataOut_payload_0_14335;
  reg        [7:0]    _zz_dataOut_payload_0_14336;
  reg        [7:0]    _zz_dataOut_payload_0_14337;
  reg        [7:0]    _zz_dataOut_payload_0_14338;
  reg        [7:0]    _zz_dataOut_payload_0_14339;
  reg        [7:0]    _zz_dataOut_payload_0_14340;
  reg        [7:0]    _zz_dataOut_payload_0_14341;
  reg        [7:0]    _zz_dataOut_payload_0_14342;
  reg        [7:0]    _zz_dataOut_payload_0_14343;
  reg        [7:0]    _zz_dataOut_payload_0_14344;
  reg        [7:0]    _zz_dataOut_payload_0_14345;
  reg        [7:0]    _zz_dataOut_payload_0_14346;
  reg        [7:0]    _zz_dataOut_payload_0_14347;
  reg        [7:0]    _zz_dataOut_payload_0_14348;
  reg        [7:0]    _zz_dataOut_payload_0_14349;
  reg        [7:0]    _zz_dataOut_payload_0_14350;
  reg        [7:0]    _zz_dataOut_payload_0_14351;
  wire                _zz_dataOut_payload_0_14352;
  wire       [7:0]    _zz_dataOut_payload_0_14353;
  wire       [7:0]    _zz_dataOut_payload_0_14354;
  wire                _zz_dataOut_payload_0_14355;
  wire       [7:0]    _zz_dataOut_payload_0_14356;
  wire       [7:0]    _zz_dataOut_payload_0_14357;
  wire                _zz_dataOut_payload_0_14358;
  wire       [7:0]    _zz_dataOut_payload_0_14359;
  wire       [7:0]    _zz_dataOut_payload_0_14360;
  wire                _zz_dataOut_payload_0_14361;
  wire       [7:0]    _zz_dataOut_payload_0_14362;
  wire       [7:0]    _zz_dataOut_payload_0_14363;
  wire                _zz_dataOut_payload_0_14364;
  wire       [7:0]    _zz_dataOut_payload_0_14365;
  wire       [7:0]    _zz_dataOut_payload_0_14366;
  wire                _zz_dataOut_payload_0_14367;
  wire       [7:0]    _zz_dataOut_payload_0_14368;
  wire       [7:0]    _zz_dataOut_payload_0_14369;
  wire                _zz_dataOut_payload_0_14370;
  wire       [7:0]    _zz_dataOut_payload_0_14371;
  wire       [7:0]    _zz_dataOut_payload_0_14372;
  wire                _zz_dataOut_payload_0_14373;
  wire       [7:0]    _zz_dataOut_payload_0_14374;
  wire       [7:0]    _zz_dataOut_payload_0_14375;
  wire                _zz_dataOut_payload_0_14376;
  wire       [7:0]    _zz_dataOut_payload_0_14377;
  wire       [7:0]    _zz_dataOut_payload_0_14378;
  wire                _zz_dataOut_payload_0_14379;
  wire       [7:0]    _zz_dataOut_payload_0_14380;
  wire       [7:0]    _zz_dataOut_payload_0_14381;
  wire                _zz_dataOut_payload_0_14382;
  wire       [7:0]    _zz_dataOut_payload_0_14383;
  wire       [7:0]    _zz_dataOut_payload_0_14384;
  wire                _zz_dataOut_payload_0_14385;
  wire       [7:0]    _zz_dataOut_payload_0_14386;
  wire       [7:0]    _zz_dataOut_payload_0_14387;
  wire                _zz_dataOut_payload_0_14388;
  wire       [7:0]    _zz_dataOut_payload_0_14389;
  wire       [7:0]    _zz_dataOut_payload_0_14390;
  wire                _zz_dataOut_payload_0_14391;
  wire       [7:0]    _zz_dataOut_payload_0_14392;
  wire       [7:0]    _zz_dataOut_payload_0_14393;
  wire                _zz_dataOut_payload_0_14394;
  wire                _zz_dataOut_payload_0_14395;
  reg        [7:0]    _zz_dataOut_payload_0_14396;
  reg        [7:0]    _zz_dataOut_payload_0_14397;
  reg        [7:0]    _zz_dataOut_payload_0_14398;
  reg        [7:0]    _zz_dataOut_payload_0_14399;
  wire                _zz_dataOut_payload_0_14400;
  wire       [7:0]    _zz_dataOut_payload_0_14401;
  wire       [7:0]    _zz_dataOut_payload_0_14402;
  wire                _zz_dataOut_payload_0_14403;
  wire       [7:0]    _zz_dataOut_payload_0_14404;
  wire       [7:0]    _zz_dataOut_payload_0_14405;
  wire                _zz_dataOut_payload_0_14406;
  wire                _zz_dataOut_payload_0_14407;
  reg        [7:0]    _zz_dataOut_payload_0_14408;
  reg        [7:0]    _zz_dataOut_payload_0_14409;
  reg        [7:0]    _zz_dataOut_payload_0_14410;
  reg        [7:0]    _zz_dataOut_payload_0_14411;
  reg        [7:0]    _zz_dataOut_payload_0_14412;
  reg        [7:0]    _zz_dataOut_payload_0_14413;
  reg        [7:0]    _zz_dataOut_payload_0_14414;
  reg        [7:0]    _zz_dataOut_payload_0_14415;
  reg        [7:0]    _zz_dataOut_payload_0_14416;
  reg        [7:0]    _zz_dataOut_payload_0_14417;
  reg        [7:0]    _zz_dataOut_payload_0_14418;
  reg        [7:0]    _zz_dataOut_payload_0_14419;
  wire                _zz_dataOut_payload_0_14420;
  wire       [7:0]    _zz_dataOut_payload_0_14421;
  wire       [7:0]    _zz_dataOut_payload_0_14422;
  wire                _zz_dataOut_payload_0_14423;
  wire       [7:0]    _zz_dataOut_payload_0_14424;
  wire       [7:0]    _zz_dataOut_payload_0_14425;
  wire                _zz_dataOut_payload_0_14426;
  wire       [7:0]    _zz_dataOut_payload_0_14427;
  wire       [7:0]    _zz_dataOut_payload_0_14428;
  wire                _zz_dataOut_payload_0_14429;
  wire       [7:0]    _zz_dataOut_payload_0_14430;
  wire       [7:0]    _zz_dataOut_payload_0_14431;
  wire                _zz_dataOut_payload_0_14432;
  wire       [7:0]    _zz_dataOut_payload_0_14433;
  wire       [7:0]    _zz_dataOut_payload_0_14434;
  wire                _zz_dataOut_payload_0_14435;
  wire       [7:0]    _zz_dataOut_payload_0_14436;
  wire       [7:0]    _zz_dataOut_payload_0_14437;
  wire                _zz_dataOut_payload_0_14438;
  wire                _zz_dataOut_payload_0_14439;
  reg        [7:0]    _zz_dataOut_payload_0_14440;
  reg        [7:0]    _zz_dataOut_payload_0_14441;
  reg        [7:0]    _zz_dataOut_payload_0_14442;
  reg        [7:0]    _zz_dataOut_payload_0_14443;
  wire                _zz_dataOut_payload_0_14444;
  wire       [7:0]    _zz_dataOut_payload_0_14445;
  wire       [7:0]    _zz_dataOut_payload_0_14446;
  wire                _zz_dataOut_payload_0_14447;
  wire       [7:0]    _zz_dataOut_payload_0_14448;
  wire       [7:0]    _zz_dataOut_payload_0_14449;
  wire                _zz_dataOut_payload_0_14450;
  wire                _zz_dataOut_payload_0_14451;
  reg        [7:0]    _zz_dataOut_payload_0_14452;
  reg        [7:0]    _zz_dataOut_payload_0_14453;
  reg        [7:0]    _zz_dataOut_payload_0_14454;
  reg        [7:0]    _zz_dataOut_payload_0_14455;
  reg        [7:0]    _zz_dataOut_payload_0_14456;
  reg        [7:0]    _zz_dataOut_payload_0_14457;
  reg        [7:0]    _zz_dataOut_payload_0_14458;
  reg        [7:0]    _zz_dataOut_payload_0_14459;
  reg        [7:0]    _zz_dataOut_payload_0_14460;
  reg        [7:0]    _zz_dataOut_payload_0_14461;
  reg        [7:0]    _zz_dataOut_payload_0_14462;
  reg        [7:0]    _zz_dataOut_payload_0_14463;
  reg        [7:0]    _zz_dataOut_payload_0_14464;
  reg        [7:0]    _zz_dataOut_payload_0_14465;
  reg        [7:0]    _zz_dataOut_payload_0_14466;
  reg        [7:0]    _zz_dataOut_payload_0_14467;
  reg        [7:0]    _zz_dataOut_payload_0_14468;
  reg        [7:0]    _zz_dataOut_payload_0_14469;
  reg        [7:0]    _zz_dataOut_payload_0_14470;
  reg        [7:0]    _zz_dataOut_payload_0_14471;
  reg        [7:0]    _zz_dataOut_payload_0_14472;
  reg        [7:0]    _zz_dataOut_payload_0_14473;
  reg        [7:0]    _zz_dataOut_payload_0_14474;
  reg        [7:0]    _zz_dataOut_payload_0_14475;
  reg        [7:0]    _zz_dataOut_payload_0_14476;
  reg        [7:0]    _zz_dataOut_payload_0_14477;
  reg        [7:0]    _zz_dataOut_payload_0_14478;
  reg        [7:0]    _zz_dataOut_payload_0_14479;
  reg        [7:0]    _zz_dataOut_payload_0_14480;
  reg        [7:0]    _zz_dataOut_payload_0_14481;
  reg        [7:0]    _zz_dataOut_payload_0_14482;
  reg        [7:0]    _zz_dataOut_payload_0_14483;
  reg        [7:0]    _zz_dataOut_payload_0_14484;
  reg        [7:0]    _zz_dataOut_payload_0_14485;
  reg        [7:0]    _zz_dataOut_payload_0_14486;
  reg        [7:0]    _zz_dataOut_payload_0_14487;
  reg        [7:0]    _zz_dataOut_payload_0_14488;
  reg        [7:0]    _zz_dataOut_payload_0_14489;
  reg        [7:0]    _zz_dataOut_payload_0_14490;
  reg        [7:0]    _zz_dataOut_payload_0_14491;
  reg        [7:0]    _zz_dataOut_payload_0_14492;
  reg        [7:0]    _zz_dataOut_payload_0_14493;
  reg        [7:0]    _zz_dataOut_payload_0_14494;
  reg        [7:0]    _zz_dataOut_payload_0_14495;
  reg        [7:0]    _zz_dataOut_payload_0_14496;
  reg        [7:0]    _zz_dataOut_payload_0_14497;
  reg        [7:0]    _zz_dataOut_payload_0_14498;
  reg        [7:0]    _zz_dataOut_payload_0_14499;
  reg        [7:0]    _zz_dataOut_payload_0_14500;
  reg        [7:0]    _zz_dataOut_payload_0_14501;
  reg        [7:0]    _zz_dataOut_payload_0_14502;
  reg        [7:0]    _zz_dataOut_payload_0_14503;
  reg        [7:0]    _zz_dataOut_payload_0_14504;
  reg        [7:0]    _zz_dataOut_payload_0_14505;
  reg        [7:0]    _zz_dataOut_payload_0_14506;
  reg        [7:0]    _zz_dataOut_payload_0_14507;
  reg        [7:0]    _zz_dataOut_payload_0_14508;
  reg        [7:0]    _zz_dataOut_payload_0_14509;
  reg        [7:0]    _zz_dataOut_payload_0_14510;
  reg        [7:0]    _zz_dataOut_payload_0_14511;
  wire                _zz_dataOut_payload_0_14512;
  wire       [7:0]    _zz_dataOut_payload_0_14513;
  wire       [7:0]    _zz_dataOut_payload_0_14514;
  wire                _zz_dataOut_payload_0_14515;
  wire       [7:0]    _zz_dataOut_payload_0_14516;
  wire       [7:0]    _zz_dataOut_payload_0_14517;
  wire                _zz_dataOut_payload_0_14518;
  wire       [7:0]    _zz_dataOut_payload_0_14519;
  wire       [7:0]    _zz_dataOut_payload_0_14520;
  wire                _zz_dataOut_payload_0_14521;
  wire       [7:0]    _zz_dataOut_payload_0_14522;
  wire       [7:0]    _zz_dataOut_payload_0_14523;
  wire                _zz_dataOut_payload_0_14524;
  wire       [7:0]    _zz_dataOut_payload_0_14525;
  wire       [7:0]    _zz_dataOut_payload_0_14526;
  wire                _zz_dataOut_payload_0_14527;
  wire       [7:0]    _zz_dataOut_payload_0_14528;
  wire       [7:0]    _zz_dataOut_payload_0_14529;
  wire                _zz_dataOut_payload_0_14530;
  wire       [7:0]    _zz_dataOut_payload_0_14531;
  wire       [7:0]    _zz_dataOut_payload_0_14532;
  wire                _zz_dataOut_payload_0_14533;
  wire       [7:0]    _zz_dataOut_payload_0_14534;
  wire       [7:0]    _zz_dataOut_payload_0_14535;
  wire                _zz_dataOut_payload_0_14536;
  wire       [7:0]    _zz_dataOut_payload_0_14537;
  wire       [7:0]    _zz_dataOut_payload_0_14538;
  wire                _zz_dataOut_payload_0_14539;
  wire       [7:0]    _zz_dataOut_payload_0_14540;
  wire       [7:0]    _zz_dataOut_payload_0_14541;
  wire                _zz_dataOut_payload_0_14542;
  wire       [7:0]    _zz_dataOut_payload_0_14543;
  wire       [7:0]    _zz_dataOut_payload_0_14544;
  wire                _zz_dataOut_payload_0_14545;
  wire       [7:0]    _zz_dataOut_payload_0_14546;
  wire       [7:0]    _zz_dataOut_payload_0_14547;
  wire                _zz_dataOut_payload_0_14548;
  wire       [7:0]    _zz_dataOut_payload_0_14549;
  wire       [7:0]    _zz_dataOut_payload_0_14550;
  wire                _zz_dataOut_payload_0_14551;
  wire       [7:0]    _zz_dataOut_payload_0_14552;
  wire       [7:0]    _zz_dataOut_payload_0_14553;
  wire                _zz_dataOut_payload_0_14554;
  wire       [7:0]    _zz_dataOut_payload_0_14555;
  wire       [7:0]    _zz_dataOut_payload_0_14556;
  wire                _zz_dataOut_payload_0_14557;
  wire       [7:0]    _zz_dataOut_payload_0_14558;
  wire       [7:0]    _zz_dataOut_payload_0_14559;
  wire                _zz_dataOut_payload_0_14560;
  wire       [7:0]    _zz_dataOut_payload_0_14561;
  wire       [7:0]    _zz_dataOut_payload_0_14562;
  wire                _zz_dataOut_payload_0_14563;
  wire       [7:0]    _zz_dataOut_payload_0_14564;
  wire       [7:0]    _zz_dataOut_payload_0_14565;
  wire                _zz_dataOut_payload_0_14566;
  wire       [7:0]    _zz_dataOut_payload_0_14567;
  wire       [7:0]    _zz_dataOut_payload_0_14568;
  wire                _zz_dataOut_payload_0_14569;
  wire       [7:0]    _zz_dataOut_payload_0_14570;
  wire       [7:0]    _zz_dataOut_payload_0_14571;
  wire                _zz_dataOut_payload_0_14572;
  wire       [7:0]    _zz_dataOut_payload_0_14573;
  wire       [7:0]    _zz_dataOut_payload_0_14574;
  wire                _zz_dataOut_payload_0_14575;
  wire       [7:0]    _zz_dataOut_payload_0_14576;
  wire       [7:0]    _zz_dataOut_payload_0_14577;
  wire                _zz_dataOut_payload_0_14578;
  wire       [7:0]    _zz_dataOut_payload_0_14579;
  wire       [7:0]    _zz_dataOut_payload_0_14580;
  wire                _zz_dataOut_payload_0_14581;
  wire       [7:0]    _zz_dataOut_payload_0_14582;
  wire       [7:0]    _zz_dataOut_payload_0_14583;
  wire                _zz_dataOut_payload_0_14584;
  wire       [7:0]    _zz_dataOut_payload_0_14585;
  wire       [7:0]    _zz_dataOut_payload_0_14586;
  wire                _zz_dataOut_payload_0_14587;
  wire       [7:0]    _zz_dataOut_payload_0_14588;
  wire       [7:0]    _zz_dataOut_payload_0_14589;
  wire                _zz_dataOut_payload_0_14590;
  wire       [7:0]    _zz_dataOut_payload_0_14591;
  wire       [7:0]    _zz_dataOut_payload_0_14592;
  wire                _zz_dataOut_payload_0_14593;
  wire       [7:0]    _zz_dataOut_payload_0_14594;
  wire       [7:0]    _zz_dataOut_payload_0_14595;
  wire                _zz_dataOut_payload_0_14596;
  wire       [7:0]    _zz_dataOut_payload_0_14597;
  wire       [7:0]    _zz_dataOut_payload_0_14598;
  wire                _zz_dataOut_payload_0_14599;
  wire       [7:0]    _zz_dataOut_payload_0_14600;
  wire       [7:0]    _zz_dataOut_payload_0_14601;
  wire                _zz_dataOut_payload_0_14602;
  wire                _zz_dataOut_payload_0_14603;
  reg        [7:0]    _zz_dataOut_payload_0_14604;
  reg        [7:0]    _zz_dataOut_payload_0_14605;
  reg        [7:0]    _zz_dataOut_payload_0_14606;
  reg        [7:0]    _zz_dataOut_payload_0_14607;
  wire                _zz_dataOut_payload_0_14608;
  wire       [7:0]    _zz_dataOut_payload_0_14609;
  wire       [7:0]    _zz_dataOut_payload_0_14610;
  wire                _zz_dataOut_payload_0_14611;
  wire       [7:0]    _zz_dataOut_payload_0_14612;
  wire       [7:0]    _zz_dataOut_payload_0_14613;
  wire                _zz_dataOut_payload_0_14614;
  wire                _zz_dataOut_payload_0_14615;
  reg        [7:0]    _zz_dataOut_payload_0_14616;
  reg        [7:0]    _zz_dataOut_payload_0_14617;
  reg        [7:0]    _zz_dataOut_payload_0_14618;
  reg        [7:0]    _zz_dataOut_payload_0_14619;
  reg        [7:0]    _zz_dataOut_payload_0_14620;
  reg        [7:0]    _zz_dataOut_payload_0_14621;
  reg        [7:0]    _zz_dataOut_payload_0_14622;
  reg        [7:0]    _zz_dataOut_payload_0_14623;
  reg        [7:0]    _zz_dataOut_payload_0_14624;
  reg        [7:0]    _zz_dataOut_payload_0_14625;
  reg        [7:0]    _zz_dataOut_payload_0_14626;
  reg        [7:0]    _zz_dataOut_payload_0_14627;
  wire                _zz_dataOut_payload_0_14628;
  wire       [7:0]    _zz_dataOut_payload_0_14629;
  wire       [7:0]    _zz_dataOut_payload_0_14630;
  wire                _zz_dataOut_payload_0_14631;
  wire       [7:0]    _zz_dataOut_payload_0_14632;
  wire       [7:0]    _zz_dataOut_payload_0_14633;
  wire                _zz_dataOut_payload_0_14634;
  wire       [7:0]    _zz_dataOut_payload_0_14635;
  wire       [7:0]    _zz_dataOut_payload_0_14636;
  wire                _zz_dataOut_payload_0_14637;
  wire       [7:0]    _zz_dataOut_payload_0_14638;
  wire       [7:0]    _zz_dataOut_payload_0_14639;
  wire                _zz_dataOut_payload_0_14640;
  wire       [7:0]    _zz_dataOut_payload_0_14641;
  wire       [7:0]    _zz_dataOut_payload_0_14642;
  wire                _zz_dataOut_payload_0_14643;
  wire       [7:0]    _zz_dataOut_payload_0_14644;
  wire       [7:0]    _zz_dataOut_payload_0_14645;
  wire                _zz_dataOut_payload_0_14646;
  wire                _zz_dataOut_payload_0_14647;
  reg        [7:0]    _zz_dataOut_payload_0_14648;
  reg        [7:0]    _zz_dataOut_payload_0_14649;
  reg        [7:0]    _zz_dataOut_payload_0_14650;
  reg        [7:0]    _zz_dataOut_payload_0_14651;
  wire                _zz_dataOut_payload_0_14652;
  wire       [7:0]    _zz_dataOut_payload_0_14653;
  wire       [7:0]    _zz_dataOut_payload_0_14654;
  wire                _zz_dataOut_payload_0_14655;
  wire       [7:0]    _zz_dataOut_payload_0_14656;
  wire       [7:0]    _zz_dataOut_payload_0_14657;
  wire                _zz_dataOut_payload_0_14658;
  wire                _zz_dataOut_payload_0_14659;
  reg        [7:0]    _zz_dataOut_payload_0_14660;
  reg        [7:0]    _zz_dataOut_payload_0_14661;
  reg        [7:0]    _zz_dataOut_payload_0_14662;
  reg        [7:0]    _zz_dataOut_payload_0_14663;
  reg        [7:0]    _zz_dataOut_payload_0_14664;
  reg        [7:0]    _zz_dataOut_payload_0_14665;
  reg        [7:0]    _zz_dataOut_payload_0_14666;
  reg        [7:0]    _zz_dataOut_payload_0_14667;
  reg        [7:0]    _zz_dataOut_payload_0_14668;
  reg        [7:0]    _zz_dataOut_payload_0_14669;
  reg        [7:0]    _zz_dataOut_payload_0_14670;
  reg        [7:0]    _zz_dataOut_payload_0_14671;
  reg        [7:0]    _zz_dataOut_payload_0_14672;
  reg        [7:0]    _zz_dataOut_payload_0_14673;
  reg        [7:0]    _zz_dataOut_payload_0_14674;
  reg        [7:0]    _zz_dataOut_payload_0_14675;
  reg        [7:0]    _zz_dataOut_payload_0_14676;
  reg        [7:0]    _zz_dataOut_payload_0_14677;
  reg        [7:0]    _zz_dataOut_payload_0_14678;
  reg        [7:0]    _zz_dataOut_payload_0_14679;
  reg        [7:0]    _zz_dataOut_payload_0_14680;
  reg        [7:0]    _zz_dataOut_payload_0_14681;
  reg        [7:0]    _zz_dataOut_payload_0_14682;
  reg        [7:0]    _zz_dataOut_payload_0_14683;
  reg        [7:0]    _zz_dataOut_payload_0_14684;
  reg        [7:0]    _zz_dataOut_payload_0_14685;
  reg        [7:0]    _zz_dataOut_payload_0_14686;
  reg        [7:0]    _zz_dataOut_payload_0_14687;
  wire                _zz_dataOut_payload_0_14688;
  wire       [7:0]    _zz_dataOut_payload_0_14689;
  wire       [7:0]    _zz_dataOut_payload_0_14690;
  wire                _zz_dataOut_payload_0_14691;
  wire       [7:0]    _zz_dataOut_payload_0_14692;
  wire       [7:0]    _zz_dataOut_payload_0_14693;
  wire                _zz_dataOut_payload_0_14694;
  wire       [7:0]    _zz_dataOut_payload_0_14695;
  wire       [7:0]    _zz_dataOut_payload_0_14696;
  wire                _zz_dataOut_payload_0_14697;
  wire       [7:0]    _zz_dataOut_payload_0_14698;
  wire       [7:0]    _zz_dataOut_payload_0_14699;
  wire                _zz_dataOut_payload_0_14700;
  wire       [7:0]    _zz_dataOut_payload_0_14701;
  wire       [7:0]    _zz_dataOut_payload_0_14702;
  wire                _zz_dataOut_payload_0_14703;
  wire       [7:0]    _zz_dataOut_payload_0_14704;
  wire       [7:0]    _zz_dataOut_payload_0_14705;
  wire                _zz_dataOut_payload_0_14706;
  wire       [7:0]    _zz_dataOut_payload_0_14707;
  wire       [7:0]    _zz_dataOut_payload_0_14708;
  wire                _zz_dataOut_payload_0_14709;
  wire       [7:0]    _zz_dataOut_payload_0_14710;
  wire       [7:0]    _zz_dataOut_payload_0_14711;
  wire                _zz_dataOut_payload_0_14712;
  wire       [7:0]    _zz_dataOut_payload_0_14713;
  wire       [7:0]    _zz_dataOut_payload_0_14714;
  wire                _zz_dataOut_payload_0_14715;
  wire       [7:0]    _zz_dataOut_payload_0_14716;
  wire       [7:0]    _zz_dataOut_payload_0_14717;
  wire                _zz_dataOut_payload_0_14718;
  wire       [7:0]    _zz_dataOut_payload_0_14719;
  wire       [7:0]    _zz_dataOut_payload_0_14720;
  wire                _zz_dataOut_payload_0_14721;
  wire       [7:0]    _zz_dataOut_payload_0_14722;
  wire       [7:0]    _zz_dataOut_payload_0_14723;
  wire                _zz_dataOut_payload_0_14724;
  wire       [7:0]    _zz_dataOut_payload_0_14725;
  wire       [7:0]    _zz_dataOut_payload_0_14726;
  wire                _zz_dataOut_payload_0_14727;
  wire       [7:0]    _zz_dataOut_payload_0_14728;
  wire       [7:0]    _zz_dataOut_payload_0_14729;
  wire                _zz_dataOut_payload_0_14730;
  wire                _zz_dataOut_payload_0_14731;
  reg        [7:0]    _zz_dataOut_payload_0_14732;
  reg        [7:0]    _zz_dataOut_payload_0_14733;
  reg        [7:0]    _zz_dataOut_payload_0_14734;
  reg        [7:0]    _zz_dataOut_payload_0_14735;
  wire                _zz_dataOut_payload_0_14736;
  wire       [7:0]    _zz_dataOut_payload_0_14737;
  wire       [7:0]    _zz_dataOut_payload_0_14738;
  wire                _zz_dataOut_payload_0_14739;
  wire       [7:0]    _zz_dataOut_payload_0_14740;
  wire       [7:0]    _zz_dataOut_payload_0_14741;
  wire                _zz_dataOut_payload_0_14742;
  wire                _zz_dataOut_payload_0_14743;
  reg        [7:0]    _zz_dataOut_payload_0_14744;
  reg        [7:0]    _zz_dataOut_payload_0_14745;
  reg        [7:0]    _zz_dataOut_payload_0_14746;
  reg        [7:0]    _zz_dataOut_payload_0_14747;
  reg        [7:0]    _zz_dataOut_payload_0_14748;
  reg        [7:0]    _zz_dataOut_payload_0_14749;
  reg        [7:0]    _zz_dataOut_payload_0_14750;
  reg        [7:0]    _zz_dataOut_payload_0_14751;
  reg        [7:0]    _zz_dataOut_payload_0_14752;
  reg        [7:0]    _zz_dataOut_payload_0_14753;
  reg        [7:0]    _zz_dataOut_payload_0_14754;
  reg        [7:0]    _zz_dataOut_payload_0_14755;
  wire                _zz_dataOut_payload_0_14756;
  wire       [7:0]    _zz_dataOut_payload_0_14757;
  wire       [7:0]    _zz_dataOut_payload_0_14758;
  wire                _zz_dataOut_payload_0_14759;
  wire       [7:0]    _zz_dataOut_payload_0_14760;
  wire       [7:0]    _zz_dataOut_payload_0_14761;
  wire                _zz_dataOut_payload_0_14762;
  wire       [7:0]    _zz_dataOut_payload_0_14763;
  wire       [7:0]    _zz_dataOut_payload_0_14764;
  wire                _zz_dataOut_payload_0_14765;
  wire       [7:0]    _zz_dataOut_payload_0_14766;
  wire       [7:0]    _zz_dataOut_payload_0_14767;
  wire                _zz_dataOut_payload_0_14768;
  wire       [7:0]    _zz_dataOut_payload_0_14769;
  wire       [7:0]    _zz_dataOut_payload_0_14770;
  wire                _zz_dataOut_payload_0_14771;
  wire       [7:0]    _zz_dataOut_payload_0_14772;
  wire       [7:0]    _zz_dataOut_payload_0_14773;
  wire                _zz_dataOut_payload_0_14774;
  wire                _zz_dataOut_payload_0_14775;
  reg        [7:0]    _zz_dataOut_payload_0_14776;
  reg        [7:0]    _zz_dataOut_payload_0_14777;
  reg        [7:0]    _zz_dataOut_payload_0_14778;
  reg        [7:0]    _zz_dataOut_payload_0_14779;
  wire                _zz_dataOut_payload_0_14780;
  wire       [7:0]    _zz_dataOut_payload_0_14781;
  wire       [7:0]    _zz_dataOut_payload_0_14782;
  wire                _zz_dataOut_payload_0_14783;
  wire       [7:0]    _zz_dataOut_payload_0_14784;
  wire       [7:0]    _zz_dataOut_payload_0_14785;
  wire                _zz_dataOut_payload_0_14786;
  wire                _zz_dataOut_payload_0_14787;
  reg        [7:0]    _zz_dataOut_payload_0_14788;
  reg        [7:0]    _zz_dataOut_payload_0_14789;
  reg        [7:0]    _zz_dataOut_payload_0_14790;
  reg        [7:0]    _zz_dataOut_payload_0_14791;
  reg        [7:0]    _zz_dataOut_payload_0_14792;
  reg        [7:0]    _zz_dataOut_payload_0_14793;
  reg        [7:0]    _zz_dataOut_payload_0_14794;
  reg        [7:0]    _zz_dataOut_payload_0_14795;
  reg        [7:0]    _zz_dataOut_payload_0_14796;
  reg        [7:0]    _zz_dataOut_payload_0_14797;
  reg        [7:0]    _zz_dataOut_payload_0_14798;
  reg        [7:0]    _zz_dataOut_payload_0_14799;
  reg        [7:0]    _zz_dataOut_payload_0_14800;
  reg        [7:0]    _zz_dataOut_payload_0_14801;
  reg        [7:0]    _zz_dataOut_payload_0_14802;
  reg        [7:0]    _zz_dataOut_payload_0_14803;
  reg        [7:0]    _zz_dataOut_payload_0_14804;
  reg        [7:0]    _zz_dataOut_payload_0_14805;
  reg        [7:0]    _zz_dataOut_payload_0_14806;
  reg        [7:0]    _zz_dataOut_payload_0_14807;
  reg        [7:0]    _zz_dataOut_payload_0_14808;
  reg        [7:0]    _zz_dataOut_payload_0_14809;
  reg        [7:0]    _zz_dataOut_payload_0_14810;
  reg        [7:0]    _zz_dataOut_payload_0_14811;
  reg        [7:0]    _zz_dataOut_payload_0_14812;
  reg        [7:0]    _zz_dataOut_payload_0_14813;
  reg        [7:0]    _zz_dataOut_payload_0_14814;
  reg        [7:0]    _zz_dataOut_payload_0_14815;
  reg        [7:0]    _zz_dataOut_payload_0_14816;
  reg        [7:0]    _zz_dataOut_payload_0_14817;
  reg        [7:0]    _zz_dataOut_payload_0_14818;
  reg        [7:0]    _zz_dataOut_payload_0_14819;
  reg        [7:0]    _zz_dataOut_payload_0_14820;
  reg        [7:0]    _zz_dataOut_payload_0_14821;
  reg        [7:0]    _zz_dataOut_payload_0_14822;
  reg        [7:0]    _zz_dataOut_payload_0_14823;
  reg        [7:0]    _zz_dataOut_payload_0_14824;
  reg        [7:0]    _zz_dataOut_payload_0_14825;
  reg        [7:0]    _zz_dataOut_payload_0_14826;
  reg        [7:0]    _zz_dataOut_payload_0_14827;
  reg        [7:0]    _zz_dataOut_payload_0_14828;
  reg        [7:0]    _zz_dataOut_payload_0_14829;
  reg        [7:0]    _zz_dataOut_payload_0_14830;
  reg        [7:0]    _zz_dataOut_payload_0_14831;
  reg        [7:0]    _zz_dataOut_payload_0_14832;
  reg        [7:0]    _zz_dataOut_payload_0_14833;
  reg        [7:0]    _zz_dataOut_payload_0_14834;
  reg        [7:0]    _zz_dataOut_payload_0_14835;
  reg        [7:0]    _zz_dataOut_payload_0_14836;
  reg        [7:0]    _zz_dataOut_payload_0_14837;
  reg        [7:0]    _zz_dataOut_payload_0_14838;
  reg        [7:0]    _zz_dataOut_payload_0_14839;
  reg        [7:0]    _zz_dataOut_payload_0_14840;
  reg        [7:0]    _zz_dataOut_payload_0_14841;
  reg        [7:0]    _zz_dataOut_payload_0_14842;
  reg        [7:0]    _zz_dataOut_payload_0_14843;
  reg        [7:0]    _zz_dataOut_payload_0_14844;
  reg        [7:0]    _zz_dataOut_payload_0_14845;
  reg        [7:0]    _zz_dataOut_payload_0_14846;
  reg        [7:0]    _zz_dataOut_payload_0_14847;
  reg        [7:0]    _zz_dataOut_payload_0_14848;
  reg        [7:0]    _zz_dataOut_payload_0_14849;
  reg        [7:0]    _zz_dataOut_payload_0_14850;
  reg        [7:0]    _zz_dataOut_payload_0_14851;
  reg        [7:0]    _zz_dataOut_payload_0_14852;
  reg        [7:0]    _zz_dataOut_payload_0_14853;
  reg        [7:0]    _zz_dataOut_payload_0_14854;
  reg        [7:0]    _zz_dataOut_payload_0_14855;
  reg        [7:0]    _zz_dataOut_payload_0_14856;
  reg        [7:0]    _zz_dataOut_payload_0_14857;
  reg        [7:0]    _zz_dataOut_payload_0_14858;
  reg        [7:0]    _zz_dataOut_payload_0_14859;
  reg        [7:0]    _zz_dataOut_payload_0_14860;
  reg        [7:0]    _zz_dataOut_payload_0_14861;
  reg        [7:0]    _zz_dataOut_payload_0_14862;
  reg        [7:0]    _zz_dataOut_payload_0_14863;
  reg        [7:0]    _zz_dataOut_payload_0_14864;
  reg        [7:0]    _zz_dataOut_payload_0_14865;
  reg        [7:0]    _zz_dataOut_payload_0_14866;
  reg        [7:0]    _zz_dataOut_payload_0_14867;
  reg        [7:0]    _zz_dataOut_payload_0_14868;
  reg        [7:0]    _zz_dataOut_payload_0_14869;
  reg        [7:0]    _zz_dataOut_payload_0_14870;
  reg        [7:0]    _zz_dataOut_payload_0_14871;
  reg        [7:0]    _zz_dataOut_payload_0_14872;
  reg        [7:0]    _zz_dataOut_payload_0_14873;
  reg        [7:0]    _zz_dataOut_payload_0_14874;
  reg        [7:0]    _zz_dataOut_payload_0_14875;
  reg        [7:0]    _zz_dataOut_payload_0_14876;
  reg        [7:0]    _zz_dataOut_payload_0_14877;
  reg        [7:0]    _zz_dataOut_payload_0_14878;
  reg        [7:0]    _zz_dataOut_payload_0_14879;
  reg        [7:0]    _zz_dataOut_payload_0_14880;
  reg        [7:0]    _zz_dataOut_payload_0_14881;
  reg        [7:0]    _zz_dataOut_payload_0_14882;
  reg        [7:0]    _zz_dataOut_payload_0_14883;
  reg        [7:0]    _zz_dataOut_payload_0_14884;
  reg        [7:0]    _zz_dataOut_payload_0_14885;
  reg        [7:0]    _zz_dataOut_payload_0_14886;
  reg        [7:0]    _zz_dataOut_payload_0_14887;
  reg        [7:0]    _zz_dataOut_payload_0_14888;
  reg        [7:0]    _zz_dataOut_payload_0_14889;
  reg        [7:0]    _zz_dataOut_payload_0_14890;
  reg        [7:0]    _zz_dataOut_payload_0_14891;
  reg        [7:0]    _zz_dataOut_payload_0_14892;
  reg        [7:0]    _zz_dataOut_payload_0_14893;
  reg        [7:0]    _zz_dataOut_payload_0_14894;
  reg        [7:0]    _zz_dataOut_payload_0_14895;
  reg        [7:0]    _zz_dataOut_payload_0_14896;
  reg        [7:0]    _zz_dataOut_payload_0_14897;
  reg        [7:0]    _zz_dataOut_payload_0_14898;
  reg        [7:0]    _zz_dataOut_payload_0_14899;
  reg        [7:0]    _zz_dataOut_payload_0_14900;
  reg        [7:0]    _zz_dataOut_payload_0_14901;
  reg        [7:0]    _zz_dataOut_payload_0_14902;
  reg        [7:0]    _zz_dataOut_payload_0_14903;
  reg        [7:0]    _zz_dataOut_payload_0_14904;
  reg        [7:0]    _zz_dataOut_payload_0_14905;
  reg        [7:0]    _zz_dataOut_payload_0_14906;
  reg        [7:0]    _zz_dataOut_payload_0_14907;
  reg        [7:0]    _zz_dataOut_payload_0_14908;
  reg        [7:0]    _zz_dataOut_payload_0_14909;
  reg        [7:0]    _zz_dataOut_payload_0_14910;
  reg        [7:0]    _zz_dataOut_payload_0_14911;
  wire                _zz_dataOut_payload_0_14912;
  wire       [7:0]    _zz_dataOut_payload_0_14913;
  wire       [7:0]    _zz_dataOut_payload_0_14914;
  wire                _zz_dataOut_payload_0_14915;
  wire       [7:0]    _zz_dataOut_payload_0_14916;
  wire       [7:0]    _zz_dataOut_payload_0_14917;
  wire                _zz_dataOut_payload_0_14918;
  wire       [7:0]    _zz_dataOut_payload_0_14919;
  wire       [7:0]    _zz_dataOut_payload_0_14920;
  wire                _zz_dataOut_payload_0_14921;
  wire       [7:0]    _zz_dataOut_payload_0_14922;
  wire       [7:0]    _zz_dataOut_payload_0_14923;
  wire                _zz_dataOut_payload_0_14924;
  wire       [7:0]    _zz_dataOut_payload_0_14925;
  wire       [7:0]    _zz_dataOut_payload_0_14926;
  wire                _zz_dataOut_payload_0_14927;
  wire       [7:0]    _zz_dataOut_payload_0_14928;
  wire       [7:0]    _zz_dataOut_payload_0_14929;
  wire                _zz_dataOut_payload_0_14930;
  wire       [7:0]    _zz_dataOut_payload_0_14931;
  wire       [7:0]    _zz_dataOut_payload_0_14932;
  wire                _zz_dataOut_payload_0_14933;
  wire       [7:0]    _zz_dataOut_payload_0_14934;
  wire       [7:0]    _zz_dataOut_payload_0_14935;
  wire                _zz_dataOut_payload_0_14936;
  wire       [7:0]    _zz_dataOut_payload_0_14937;
  wire       [7:0]    _zz_dataOut_payload_0_14938;
  wire                _zz_dataOut_payload_0_14939;
  wire       [7:0]    _zz_dataOut_payload_0_14940;
  wire       [7:0]    _zz_dataOut_payload_0_14941;
  wire                _zz_dataOut_payload_0_14942;
  wire       [7:0]    _zz_dataOut_payload_0_14943;
  wire       [7:0]    _zz_dataOut_payload_0_14944;
  wire                _zz_dataOut_payload_0_14945;
  wire       [7:0]    _zz_dataOut_payload_0_14946;
  wire       [7:0]    _zz_dataOut_payload_0_14947;
  wire                _zz_dataOut_payload_0_14948;
  wire       [7:0]    _zz_dataOut_payload_0_14949;
  wire       [7:0]    _zz_dataOut_payload_0_14950;
  wire                _zz_dataOut_payload_0_14951;
  wire       [7:0]    _zz_dataOut_payload_0_14952;
  wire       [7:0]    _zz_dataOut_payload_0_14953;
  wire                _zz_dataOut_payload_0_14954;
  wire       [7:0]    _zz_dataOut_payload_0_14955;
  wire       [7:0]    _zz_dataOut_payload_0_14956;
  wire                _zz_dataOut_payload_0_14957;
  wire       [7:0]    _zz_dataOut_payload_0_14958;
  wire       [7:0]    _zz_dataOut_payload_0_14959;
  wire                _zz_dataOut_payload_0_14960;
  wire       [7:0]    _zz_dataOut_payload_0_14961;
  wire       [7:0]    _zz_dataOut_payload_0_14962;
  wire                _zz_dataOut_payload_0_14963;
  wire       [7:0]    _zz_dataOut_payload_0_14964;
  wire       [7:0]    _zz_dataOut_payload_0_14965;
  wire                _zz_dataOut_payload_0_14966;
  wire       [7:0]    _zz_dataOut_payload_0_14967;
  wire       [7:0]    _zz_dataOut_payload_0_14968;
  wire                _zz_dataOut_payload_0_14969;
  wire       [7:0]    _zz_dataOut_payload_0_14970;
  wire       [7:0]    _zz_dataOut_payload_0_14971;
  wire                _zz_dataOut_payload_0_14972;
  wire       [7:0]    _zz_dataOut_payload_0_14973;
  wire       [7:0]    _zz_dataOut_payload_0_14974;
  wire                _zz_dataOut_payload_0_14975;
  wire       [7:0]    _zz_dataOut_payload_0_14976;
  wire       [7:0]    _zz_dataOut_payload_0_14977;
  wire                _zz_dataOut_payload_0_14978;
  wire       [7:0]    _zz_dataOut_payload_0_14979;
  wire       [7:0]    _zz_dataOut_payload_0_14980;
  wire                _zz_dataOut_payload_0_14981;
  wire       [7:0]    _zz_dataOut_payload_0_14982;
  wire       [7:0]    _zz_dataOut_payload_0_14983;
  wire                _zz_dataOut_payload_0_14984;
  wire       [7:0]    _zz_dataOut_payload_0_14985;
  wire       [7:0]    _zz_dataOut_payload_0_14986;
  wire                _zz_dataOut_payload_0_14987;
  wire       [7:0]    _zz_dataOut_payload_0_14988;
  wire       [7:0]    _zz_dataOut_payload_0_14989;
  wire                _zz_dataOut_payload_0_14990;
  wire       [7:0]    _zz_dataOut_payload_0_14991;
  wire       [7:0]    _zz_dataOut_payload_0_14992;
  wire                _zz_dataOut_payload_0_14993;
  wire       [7:0]    _zz_dataOut_payload_0_14994;
  wire       [7:0]    _zz_dataOut_payload_0_14995;
  wire                _zz_dataOut_payload_0_14996;
  wire       [7:0]    _zz_dataOut_payload_0_14997;
  wire       [7:0]    _zz_dataOut_payload_0_14998;
  wire                _zz_dataOut_payload_0_14999;
  wire       [7:0]    _zz_dataOut_payload_0_15000;
  wire       [7:0]    _zz_dataOut_payload_0_15001;
  wire                _zz_dataOut_payload_0_15002;
  wire       [7:0]    _zz_dataOut_payload_0_15003;
  wire       [7:0]    _zz_dataOut_payload_0_15004;
  wire                _zz_dataOut_payload_0_15005;
  wire       [7:0]    _zz_dataOut_payload_0_15006;
  wire       [7:0]    _zz_dataOut_payload_0_15007;
  wire                _zz_dataOut_payload_0_15008;
  wire       [7:0]    _zz_dataOut_payload_0_15009;
  wire       [7:0]    _zz_dataOut_payload_0_15010;
  wire                _zz_dataOut_payload_0_15011;
  wire       [7:0]    _zz_dataOut_payload_0_15012;
  wire       [7:0]    _zz_dataOut_payload_0_15013;
  wire                _zz_dataOut_payload_0_15014;
  wire       [7:0]    _zz_dataOut_payload_0_15015;
  wire       [7:0]    _zz_dataOut_payload_0_15016;
  wire                _zz_dataOut_payload_0_15017;
  wire       [7:0]    _zz_dataOut_payload_0_15018;
  wire       [7:0]    _zz_dataOut_payload_0_15019;
  wire                _zz_dataOut_payload_0_15020;
  wire       [7:0]    _zz_dataOut_payload_0_15021;
  wire       [7:0]    _zz_dataOut_payload_0_15022;
  wire                _zz_dataOut_payload_0_15023;
  wire       [7:0]    _zz_dataOut_payload_0_15024;
  wire       [7:0]    _zz_dataOut_payload_0_15025;
  wire                _zz_dataOut_payload_0_15026;
  wire       [7:0]    _zz_dataOut_payload_0_15027;
  wire       [7:0]    _zz_dataOut_payload_0_15028;
  wire                _zz_dataOut_payload_0_15029;
  wire       [7:0]    _zz_dataOut_payload_0_15030;
  wire       [7:0]    _zz_dataOut_payload_0_15031;
  wire                _zz_dataOut_payload_0_15032;
  wire       [7:0]    _zz_dataOut_payload_0_15033;
  wire       [7:0]    _zz_dataOut_payload_0_15034;
  wire                _zz_dataOut_payload_0_15035;
  wire       [7:0]    _zz_dataOut_payload_0_15036;
  wire       [7:0]    _zz_dataOut_payload_0_15037;
  wire                _zz_dataOut_payload_0_15038;
  wire       [7:0]    _zz_dataOut_payload_0_15039;
  wire       [7:0]    _zz_dataOut_payload_0_15040;
  wire                _zz_dataOut_payload_0_15041;
  wire       [7:0]    _zz_dataOut_payload_0_15042;
  wire       [7:0]    _zz_dataOut_payload_0_15043;
  wire                _zz_dataOut_payload_0_15044;
  wire       [7:0]    _zz_dataOut_payload_0_15045;
  wire       [7:0]    _zz_dataOut_payload_0_15046;
  wire                _zz_dataOut_payload_0_15047;
  wire       [7:0]    _zz_dataOut_payload_0_15048;
  wire       [7:0]    _zz_dataOut_payload_0_15049;
  wire                _zz_dataOut_payload_0_15050;
  wire       [7:0]    _zz_dataOut_payload_0_15051;
  wire       [7:0]    _zz_dataOut_payload_0_15052;
  wire                _zz_dataOut_payload_0_15053;
  wire       [7:0]    _zz_dataOut_payload_0_15054;
  wire       [7:0]    _zz_dataOut_payload_0_15055;
  wire                _zz_dataOut_payload_0_15056;
  wire       [7:0]    _zz_dataOut_payload_0_15057;
  wire       [7:0]    _zz_dataOut_payload_0_15058;
  wire                _zz_dataOut_payload_0_15059;
  wire       [7:0]    _zz_dataOut_payload_0_15060;
  wire       [7:0]    _zz_dataOut_payload_0_15061;
  wire                _zz_dataOut_payload_0_15062;
  wire       [7:0]    _zz_dataOut_payload_0_15063;
  wire       [7:0]    _zz_dataOut_payload_0_15064;
  wire                _zz_dataOut_payload_0_15065;
  wire       [7:0]    _zz_dataOut_payload_0_15066;
  wire       [7:0]    _zz_dataOut_payload_0_15067;
  wire                _zz_dataOut_payload_0_15068;
  wire       [7:0]    _zz_dataOut_payload_0_15069;
  wire       [7:0]    _zz_dataOut_payload_0_15070;
  wire                _zz_dataOut_payload_0_15071;
  wire       [7:0]    _zz_dataOut_payload_0_15072;
  wire       [7:0]    _zz_dataOut_payload_0_15073;
  wire                _zz_dataOut_payload_0_15074;
  wire       [7:0]    _zz_dataOut_payload_0_15075;
  wire       [7:0]    _zz_dataOut_payload_0_15076;
  wire                _zz_dataOut_payload_0_15077;
  wire       [7:0]    _zz_dataOut_payload_0_15078;
  wire       [7:0]    _zz_dataOut_payload_0_15079;
  wire                _zz_dataOut_payload_0_15080;
  wire       [7:0]    _zz_dataOut_payload_0_15081;
  wire       [7:0]    _zz_dataOut_payload_0_15082;
  wire                _zz_dataOut_payload_0_15083;
  wire       [7:0]    _zz_dataOut_payload_0_15084;
  wire       [7:0]    _zz_dataOut_payload_0_15085;
  wire                _zz_dataOut_payload_0_15086;
  wire       [7:0]    _zz_dataOut_payload_0_15087;
  wire       [7:0]    _zz_dataOut_payload_0_15088;
  wire                _zz_dataOut_payload_0_15089;
  wire       [7:0]    _zz_dataOut_payload_0_15090;
  wire       [7:0]    _zz_dataOut_payload_0_15091;
  wire                _zz_dataOut_payload_0_15092;
  wire       [7:0]    _zz_dataOut_payload_0_15093;
  wire       [7:0]    _zz_dataOut_payload_0_15094;
  wire                _zz_dataOut_payload_0_15095;
  wire       [7:0]    _zz_dataOut_payload_0_15096;
  wire       [7:0]    _zz_dataOut_payload_0_15097;
  wire                _zz_dataOut_payload_0_15098;
  wire                _zz_dataOut_payload_0_15099;
  reg        [7:0]    _zz_dataOut_payload_0_15100;
  reg        [7:0]    _zz_dataOut_payload_0_15101;
  reg        [7:0]    _zz_dataOut_payload_0_15102;
  reg        [7:0]    _zz_dataOut_payload_0_15103;
  wire                _zz_dataOut_payload_0_15104;
  wire       [7:0]    _zz_dataOut_payload_0_15105;
  wire       [7:0]    _zz_dataOut_payload_0_15106;
  wire                _zz_dataOut_payload_0_15107;
  wire       [7:0]    _zz_dataOut_payload_0_15108;
  wire       [7:0]    _zz_dataOut_payload_0_15109;
  wire                _zz_dataOut_payload_0_15110;
  wire                _zz_dataOut_payload_0_15111;
  reg        [7:0]    _zz_dataOut_payload_0_15112;
  reg        [7:0]    _zz_dataOut_payload_0_15113;
  reg        [7:0]    _zz_dataOut_payload_0_15114;
  reg        [7:0]    _zz_dataOut_payload_0_15115;
  reg        [7:0]    _zz_dataOut_payload_0_15116;
  reg        [7:0]    _zz_dataOut_payload_0_15117;
  reg        [7:0]    _zz_dataOut_payload_0_15118;
  reg        [7:0]    _zz_dataOut_payload_0_15119;
  reg        [7:0]    _zz_dataOut_payload_0_15120;
  reg        [7:0]    _zz_dataOut_payload_0_15121;
  reg        [7:0]    _zz_dataOut_payload_0_15122;
  reg        [7:0]    _zz_dataOut_payload_0_15123;
  wire                _zz_dataOut_payload_0_15124;
  wire       [7:0]    _zz_dataOut_payload_0_15125;
  wire       [7:0]    _zz_dataOut_payload_0_15126;
  wire                _zz_dataOut_payload_0_15127;
  wire       [7:0]    _zz_dataOut_payload_0_15128;
  wire       [7:0]    _zz_dataOut_payload_0_15129;
  wire                _zz_dataOut_payload_0_15130;
  wire       [7:0]    _zz_dataOut_payload_0_15131;
  wire       [7:0]    _zz_dataOut_payload_0_15132;
  wire                _zz_dataOut_payload_0_15133;
  wire       [7:0]    _zz_dataOut_payload_0_15134;
  wire       [7:0]    _zz_dataOut_payload_0_15135;
  wire                _zz_dataOut_payload_0_15136;
  wire       [7:0]    _zz_dataOut_payload_0_15137;
  wire       [7:0]    _zz_dataOut_payload_0_15138;
  wire                _zz_dataOut_payload_0_15139;
  wire       [7:0]    _zz_dataOut_payload_0_15140;
  wire       [7:0]    _zz_dataOut_payload_0_15141;
  wire                _zz_dataOut_payload_0_15142;
  wire                _zz_dataOut_payload_0_15143;
  reg        [7:0]    _zz_dataOut_payload_0_15144;
  reg        [7:0]    _zz_dataOut_payload_0_15145;
  reg        [7:0]    _zz_dataOut_payload_0_15146;
  reg        [7:0]    _zz_dataOut_payload_0_15147;
  wire                _zz_dataOut_payload_0_15148;
  wire       [7:0]    _zz_dataOut_payload_0_15149;
  wire       [7:0]    _zz_dataOut_payload_0_15150;
  wire                _zz_dataOut_payload_0_15151;
  wire       [7:0]    _zz_dataOut_payload_0_15152;
  wire       [7:0]    _zz_dataOut_payload_0_15153;
  wire                _zz_dataOut_payload_0_15154;
  wire                _zz_dataOut_payload_0_15155;
  reg        [7:0]    _zz_dataOut_payload_0_15156;
  reg        [7:0]    _zz_dataOut_payload_0_15157;
  reg        [7:0]    _zz_dataOut_payload_0_15158;
  reg        [7:0]    _zz_dataOut_payload_0_15159;
  reg        [7:0]    _zz_dataOut_payload_0_15160;
  reg        [7:0]    _zz_dataOut_payload_0_15161;
  reg        [7:0]    _zz_dataOut_payload_0_15162;
  reg        [7:0]    _zz_dataOut_payload_0_15163;
  reg        [7:0]    _zz_dataOut_payload_0_15164;
  reg        [7:0]    _zz_dataOut_payload_0_15165;
  reg        [7:0]    _zz_dataOut_payload_0_15166;
  reg        [7:0]    _zz_dataOut_payload_0_15167;
  reg        [7:0]    _zz_dataOut_payload_0_15168;
  reg        [7:0]    _zz_dataOut_payload_0_15169;
  reg        [7:0]    _zz_dataOut_payload_0_15170;
  reg        [7:0]    _zz_dataOut_payload_0_15171;
  reg        [7:0]    _zz_dataOut_payload_0_15172;
  reg        [7:0]    _zz_dataOut_payload_0_15173;
  reg        [7:0]    _zz_dataOut_payload_0_15174;
  reg        [7:0]    _zz_dataOut_payload_0_15175;
  reg        [7:0]    _zz_dataOut_payload_0_15176;
  reg        [7:0]    _zz_dataOut_payload_0_15177;
  reg        [7:0]    _zz_dataOut_payload_0_15178;
  reg        [7:0]    _zz_dataOut_payload_0_15179;
  reg        [7:0]    _zz_dataOut_payload_0_15180;
  reg        [7:0]    _zz_dataOut_payload_0_15181;
  reg        [7:0]    _zz_dataOut_payload_0_15182;
  reg        [7:0]    _zz_dataOut_payload_0_15183;
  wire                _zz_dataOut_payload_0_15184;
  wire       [7:0]    _zz_dataOut_payload_0_15185;
  wire       [7:0]    _zz_dataOut_payload_0_15186;
  wire                _zz_dataOut_payload_0_15187;
  wire       [7:0]    _zz_dataOut_payload_0_15188;
  wire       [7:0]    _zz_dataOut_payload_0_15189;
  wire                _zz_dataOut_payload_0_15190;
  wire       [7:0]    _zz_dataOut_payload_0_15191;
  wire       [7:0]    _zz_dataOut_payload_0_15192;
  wire                _zz_dataOut_payload_0_15193;
  wire       [7:0]    _zz_dataOut_payload_0_15194;
  wire       [7:0]    _zz_dataOut_payload_0_15195;
  wire                _zz_dataOut_payload_0_15196;
  wire       [7:0]    _zz_dataOut_payload_0_15197;
  wire       [7:0]    _zz_dataOut_payload_0_15198;
  wire                _zz_dataOut_payload_0_15199;
  wire       [7:0]    _zz_dataOut_payload_0_15200;
  wire       [7:0]    _zz_dataOut_payload_0_15201;
  wire                _zz_dataOut_payload_0_15202;
  wire       [7:0]    _zz_dataOut_payload_0_15203;
  wire       [7:0]    _zz_dataOut_payload_0_15204;
  wire                _zz_dataOut_payload_0_15205;
  wire       [7:0]    _zz_dataOut_payload_0_15206;
  wire       [7:0]    _zz_dataOut_payload_0_15207;
  wire                _zz_dataOut_payload_0_15208;
  wire       [7:0]    _zz_dataOut_payload_0_15209;
  wire       [7:0]    _zz_dataOut_payload_0_15210;
  wire                _zz_dataOut_payload_0_15211;
  wire       [7:0]    _zz_dataOut_payload_0_15212;
  wire       [7:0]    _zz_dataOut_payload_0_15213;
  wire                _zz_dataOut_payload_0_15214;
  wire       [7:0]    _zz_dataOut_payload_0_15215;
  wire       [7:0]    _zz_dataOut_payload_0_15216;
  wire                _zz_dataOut_payload_0_15217;
  wire       [7:0]    _zz_dataOut_payload_0_15218;
  wire       [7:0]    _zz_dataOut_payload_0_15219;
  wire                _zz_dataOut_payload_0_15220;
  wire       [7:0]    _zz_dataOut_payload_0_15221;
  wire       [7:0]    _zz_dataOut_payload_0_15222;
  wire                _zz_dataOut_payload_0_15223;
  wire       [7:0]    _zz_dataOut_payload_0_15224;
  wire       [7:0]    _zz_dataOut_payload_0_15225;
  wire                _zz_dataOut_payload_0_15226;
  wire                _zz_dataOut_payload_0_15227;
  reg        [7:0]    _zz_dataOut_payload_0_15228;
  reg        [7:0]    _zz_dataOut_payload_0_15229;
  reg        [7:0]    _zz_dataOut_payload_0_15230;
  reg        [7:0]    _zz_dataOut_payload_0_15231;
  wire                _zz_dataOut_payload_0_15232;
  wire       [7:0]    _zz_dataOut_payload_0_15233;
  wire       [7:0]    _zz_dataOut_payload_0_15234;
  wire                _zz_dataOut_payload_0_15235;
  wire       [7:0]    _zz_dataOut_payload_0_15236;
  wire       [7:0]    _zz_dataOut_payload_0_15237;
  wire                _zz_dataOut_payload_0_15238;
  wire                _zz_dataOut_payload_0_15239;
  reg        [7:0]    _zz_dataOut_payload_0_15240;
  reg        [7:0]    _zz_dataOut_payload_0_15241;
  reg        [7:0]    _zz_dataOut_payload_0_15242;
  reg        [7:0]    _zz_dataOut_payload_0_15243;
  reg        [7:0]    _zz_dataOut_payload_0_15244;
  reg        [7:0]    _zz_dataOut_payload_0_15245;
  reg        [7:0]    _zz_dataOut_payload_0_15246;
  reg        [7:0]    _zz_dataOut_payload_0_15247;
  reg        [7:0]    _zz_dataOut_payload_0_15248;
  reg        [7:0]    _zz_dataOut_payload_0_15249;
  reg        [7:0]    _zz_dataOut_payload_0_15250;
  reg        [7:0]    _zz_dataOut_payload_0_15251;
  wire                _zz_dataOut_payload_0_15252;
  wire       [7:0]    _zz_dataOut_payload_0_15253;
  wire       [7:0]    _zz_dataOut_payload_0_15254;
  wire                _zz_dataOut_payload_0_15255;
  wire       [7:0]    _zz_dataOut_payload_0_15256;
  wire       [7:0]    _zz_dataOut_payload_0_15257;
  wire                _zz_dataOut_payload_0_15258;
  wire       [7:0]    _zz_dataOut_payload_0_15259;
  wire       [7:0]    _zz_dataOut_payload_0_15260;
  wire                _zz_dataOut_payload_0_15261;
  wire       [7:0]    _zz_dataOut_payload_0_15262;
  wire       [7:0]    _zz_dataOut_payload_0_15263;
  wire                _zz_dataOut_payload_0_15264;
  wire       [7:0]    _zz_dataOut_payload_0_15265;
  wire       [7:0]    _zz_dataOut_payload_0_15266;
  wire                _zz_dataOut_payload_0_15267;
  wire       [7:0]    _zz_dataOut_payload_0_15268;
  wire       [7:0]    _zz_dataOut_payload_0_15269;
  wire                _zz_dataOut_payload_0_15270;
  wire                _zz_dataOut_payload_0_15271;
  reg        [7:0]    _zz_dataOut_payload_0_15272;
  reg        [7:0]    _zz_dataOut_payload_0_15273;
  reg        [7:0]    _zz_dataOut_payload_0_15274;
  reg        [7:0]    _zz_dataOut_payload_0_15275;
  wire                _zz_dataOut_payload_0_15276;
  wire       [7:0]    _zz_dataOut_payload_0_15277;
  wire       [7:0]    _zz_dataOut_payload_0_15278;
  wire                _zz_dataOut_payload_0_15279;
  wire       [7:0]    _zz_dataOut_payload_0_15280;
  wire       [7:0]    _zz_dataOut_payload_0_15281;
  wire                _zz_dataOut_payload_0_15282;
  wire                _zz_dataOut_payload_0_15283;
  reg        [7:0]    _zz_dataOut_payload_0_15284;
  reg        [7:0]    _zz_dataOut_payload_0_15285;
  reg        [7:0]    _zz_dataOut_payload_0_15286;
  reg        [7:0]    _zz_dataOut_payload_0_15287;
  reg        [7:0]    _zz_dataOut_payload_0_15288;
  reg        [7:0]    _zz_dataOut_payload_0_15289;
  reg        [7:0]    _zz_dataOut_payload_0_15290;
  reg        [7:0]    _zz_dataOut_payload_0_15291;
  reg        [7:0]    _zz_dataOut_payload_0_15292;
  reg        [7:0]    _zz_dataOut_payload_0_15293;
  reg        [7:0]    _zz_dataOut_payload_0_15294;
  reg        [7:0]    _zz_dataOut_payload_0_15295;
  reg        [7:0]    _zz_dataOut_payload_0_15296;
  reg        [7:0]    _zz_dataOut_payload_0_15297;
  reg        [7:0]    _zz_dataOut_payload_0_15298;
  reg        [7:0]    _zz_dataOut_payload_0_15299;
  reg        [7:0]    _zz_dataOut_payload_0_15300;
  reg        [7:0]    _zz_dataOut_payload_0_15301;
  reg        [7:0]    _zz_dataOut_payload_0_15302;
  reg        [7:0]    _zz_dataOut_payload_0_15303;
  reg        [7:0]    _zz_dataOut_payload_0_15304;
  reg        [7:0]    _zz_dataOut_payload_0_15305;
  reg        [7:0]    _zz_dataOut_payload_0_15306;
  reg        [7:0]    _zz_dataOut_payload_0_15307;
  reg        [7:0]    _zz_dataOut_payload_0_15308;
  reg        [7:0]    _zz_dataOut_payload_0_15309;
  reg        [7:0]    _zz_dataOut_payload_0_15310;
  reg        [7:0]    _zz_dataOut_payload_0_15311;
  reg        [7:0]    _zz_dataOut_payload_0_15312;
  reg        [7:0]    _zz_dataOut_payload_0_15313;
  reg        [7:0]    _zz_dataOut_payload_0_15314;
  reg        [7:0]    _zz_dataOut_payload_0_15315;
  reg        [7:0]    _zz_dataOut_payload_0_15316;
  reg        [7:0]    _zz_dataOut_payload_0_15317;
  reg        [7:0]    _zz_dataOut_payload_0_15318;
  reg        [7:0]    _zz_dataOut_payload_0_15319;
  reg        [7:0]    _zz_dataOut_payload_0_15320;
  reg        [7:0]    _zz_dataOut_payload_0_15321;
  reg        [7:0]    _zz_dataOut_payload_0_15322;
  reg        [7:0]    _zz_dataOut_payload_0_15323;
  reg        [7:0]    _zz_dataOut_payload_0_15324;
  reg        [7:0]    _zz_dataOut_payload_0_15325;
  reg        [7:0]    _zz_dataOut_payload_0_15326;
  reg        [7:0]    _zz_dataOut_payload_0_15327;
  reg        [7:0]    _zz_dataOut_payload_0_15328;
  reg        [7:0]    _zz_dataOut_payload_0_15329;
  reg        [7:0]    _zz_dataOut_payload_0_15330;
  reg        [7:0]    _zz_dataOut_payload_0_15331;
  reg        [7:0]    _zz_dataOut_payload_0_15332;
  reg        [7:0]    _zz_dataOut_payload_0_15333;
  reg        [7:0]    _zz_dataOut_payload_0_15334;
  reg        [7:0]    _zz_dataOut_payload_0_15335;
  reg        [7:0]    _zz_dataOut_payload_0_15336;
  reg        [7:0]    _zz_dataOut_payload_0_15337;
  reg        [7:0]    _zz_dataOut_payload_0_15338;
  reg        [7:0]    _zz_dataOut_payload_0_15339;
  reg        [7:0]    _zz_dataOut_payload_0_15340;
  reg        [7:0]    _zz_dataOut_payload_0_15341;
  reg        [7:0]    _zz_dataOut_payload_0_15342;
  reg        [7:0]    _zz_dataOut_payload_0_15343;
  wire                _zz_dataOut_payload_0_15344;
  wire       [7:0]    _zz_dataOut_payload_0_15345;
  wire       [7:0]    _zz_dataOut_payload_0_15346;
  wire                _zz_dataOut_payload_0_15347;
  wire       [7:0]    _zz_dataOut_payload_0_15348;
  wire       [7:0]    _zz_dataOut_payload_0_15349;
  wire                _zz_dataOut_payload_0_15350;
  wire       [7:0]    _zz_dataOut_payload_0_15351;
  wire       [7:0]    _zz_dataOut_payload_0_15352;
  wire                _zz_dataOut_payload_0_15353;
  wire       [7:0]    _zz_dataOut_payload_0_15354;
  wire       [7:0]    _zz_dataOut_payload_0_15355;
  wire                _zz_dataOut_payload_0_15356;
  wire       [7:0]    _zz_dataOut_payload_0_15357;
  wire       [7:0]    _zz_dataOut_payload_0_15358;
  wire                _zz_dataOut_payload_0_15359;
  wire       [7:0]    _zz_dataOut_payload_0_15360;
  wire       [7:0]    _zz_dataOut_payload_0_15361;
  wire                _zz_dataOut_payload_0_15362;
  wire       [7:0]    _zz_dataOut_payload_0_15363;
  wire       [7:0]    _zz_dataOut_payload_0_15364;
  wire                _zz_dataOut_payload_0_15365;
  wire       [7:0]    _zz_dataOut_payload_0_15366;
  wire       [7:0]    _zz_dataOut_payload_0_15367;
  wire                _zz_dataOut_payload_0_15368;
  wire       [7:0]    _zz_dataOut_payload_0_15369;
  wire       [7:0]    _zz_dataOut_payload_0_15370;
  wire                _zz_dataOut_payload_0_15371;
  wire       [7:0]    _zz_dataOut_payload_0_15372;
  wire       [7:0]    _zz_dataOut_payload_0_15373;
  wire                _zz_dataOut_payload_0_15374;
  wire       [7:0]    _zz_dataOut_payload_0_15375;
  wire       [7:0]    _zz_dataOut_payload_0_15376;
  wire                _zz_dataOut_payload_0_15377;
  wire       [7:0]    _zz_dataOut_payload_0_15378;
  wire       [7:0]    _zz_dataOut_payload_0_15379;
  wire                _zz_dataOut_payload_0_15380;
  wire       [7:0]    _zz_dataOut_payload_0_15381;
  wire       [7:0]    _zz_dataOut_payload_0_15382;
  wire                _zz_dataOut_payload_0_15383;
  wire       [7:0]    _zz_dataOut_payload_0_15384;
  wire       [7:0]    _zz_dataOut_payload_0_15385;
  wire                _zz_dataOut_payload_0_15386;
  wire       [7:0]    _zz_dataOut_payload_0_15387;
  wire       [7:0]    _zz_dataOut_payload_0_15388;
  wire                _zz_dataOut_payload_0_15389;
  wire       [7:0]    _zz_dataOut_payload_0_15390;
  wire       [7:0]    _zz_dataOut_payload_0_15391;
  wire                _zz_dataOut_payload_0_15392;
  wire       [7:0]    _zz_dataOut_payload_0_15393;
  wire       [7:0]    _zz_dataOut_payload_0_15394;
  wire                _zz_dataOut_payload_0_15395;
  wire       [7:0]    _zz_dataOut_payload_0_15396;
  wire       [7:0]    _zz_dataOut_payload_0_15397;
  wire                _zz_dataOut_payload_0_15398;
  wire       [7:0]    _zz_dataOut_payload_0_15399;
  wire       [7:0]    _zz_dataOut_payload_0_15400;
  wire                _zz_dataOut_payload_0_15401;
  wire       [7:0]    _zz_dataOut_payload_0_15402;
  wire       [7:0]    _zz_dataOut_payload_0_15403;
  wire                _zz_dataOut_payload_0_15404;
  wire       [7:0]    _zz_dataOut_payload_0_15405;
  wire       [7:0]    _zz_dataOut_payload_0_15406;
  wire                _zz_dataOut_payload_0_15407;
  wire       [7:0]    _zz_dataOut_payload_0_15408;
  wire       [7:0]    _zz_dataOut_payload_0_15409;
  wire                _zz_dataOut_payload_0_15410;
  wire       [7:0]    _zz_dataOut_payload_0_15411;
  wire       [7:0]    _zz_dataOut_payload_0_15412;
  wire                _zz_dataOut_payload_0_15413;
  wire       [7:0]    _zz_dataOut_payload_0_15414;
  wire       [7:0]    _zz_dataOut_payload_0_15415;
  wire                _zz_dataOut_payload_0_15416;
  wire       [7:0]    _zz_dataOut_payload_0_15417;
  wire       [7:0]    _zz_dataOut_payload_0_15418;
  wire                _zz_dataOut_payload_0_15419;
  wire       [7:0]    _zz_dataOut_payload_0_15420;
  wire       [7:0]    _zz_dataOut_payload_0_15421;
  wire                _zz_dataOut_payload_0_15422;
  wire       [7:0]    _zz_dataOut_payload_0_15423;
  wire       [7:0]    _zz_dataOut_payload_0_15424;
  wire                _zz_dataOut_payload_0_15425;
  wire       [7:0]    _zz_dataOut_payload_0_15426;
  wire       [7:0]    _zz_dataOut_payload_0_15427;
  wire                _zz_dataOut_payload_0_15428;
  wire       [7:0]    _zz_dataOut_payload_0_15429;
  wire       [7:0]    _zz_dataOut_payload_0_15430;
  wire                _zz_dataOut_payload_0_15431;
  wire       [7:0]    _zz_dataOut_payload_0_15432;
  wire       [7:0]    _zz_dataOut_payload_0_15433;
  wire                _zz_dataOut_payload_0_15434;
  wire                _zz_dataOut_payload_0_15435;
  reg        [7:0]    _zz_dataOut_payload_0_15436;
  reg        [7:0]    _zz_dataOut_payload_0_15437;
  reg        [7:0]    _zz_dataOut_payload_0_15438;
  reg        [7:0]    _zz_dataOut_payload_0_15439;
  wire                _zz_dataOut_payload_0_15440;
  wire       [7:0]    _zz_dataOut_payload_0_15441;
  wire       [7:0]    _zz_dataOut_payload_0_15442;
  wire                _zz_dataOut_payload_0_15443;
  wire       [7:0]    _zz_dataOut_payload_0_15444;
  wire       [7:0]    _zz_dataOut_payload_0_15445;
  wire                _zz_dataOut_payload_0_15446;
  wire                _zz_dataOut_payload_0_15447;
  reg        [7:0]    _zz_dataOut_payload_0_15448;
  reg        [7:0]    _zz_dataOut_payload_0_15449;
  reg        [7:0]    _zz_dataOut_payload_0_15450;
  reg        [7:0]    _zz_dataOut_payload_0_15451;
  reg        [7:0]    _zz_dataOut_payload_0_15452;
  reg        [7:0]    _zz_dataOut_payload_0_15453;
  reg        [7:0]    _zz_dataOut_payload_0_15454;
  reg        [7:0]    _zz_dataOut_payload_0_15455;
  reg        [7:0]    _zz_dataOut_payload_0_15456;
  reg        [7:0]    _zz_dataOut_payload_0_15457;
  reg        [7:0]    _zz_dataOut_payload_0_15458;
  reg        [7:0]    _zz_dataOut_payload_0_15459;
  wire                _zz_dataOut_payload_0_15460;
  wire       [7:0]    _zz_dataOut_payload_0_15461;
  wire       [7:0]    _zz_dataOut_payload_0_15462;
  wire                _zz_dataOut_payload_0_15463;
  wire       [7:0]    _zz_dataOut_payload_0_15464;
  wire       [7:0]    _zz_dataOut_payload_0_15465;
  wire                _zz_dataOut_payload_0_15466;
  wire       [7:0]    _zz_dataOut_payload_0_15467;
  wire       [7:0]    _zz_dataOut_payload_0_15468;
  wire                _zz_dataOut_payload_0_15469;
  wire       [7:0]    _zz_dataOut_payload_0_15470;
  wire       [7:0]    _zz_dataOut_payload_0_15471;
  wire                _zz_dataOut_payload_0_15472;
  wire       [7:0]    _zz_dataOut_payload_0_15473;
  wire       [7:0]    _zz_dataOut_payload_0_15474;
  wire                _zz_dataOut_payload_0_15475;
  wire       [7:0]    _zz_dataOut_payload_0_15476;
  wire       [7:0]    _zz_dataOut_payload_0_15477;
  wire                _zz_dataOut_payload_0_15478;
  wire                _zz_dataOut_payload_0_15479;
  reg        [7:0]    _zz_dataOut_payload_0_15480;
  reg        [7:0]    _zz_dataOut_payload_0_15481;
  reg        [7:0]    _zz_dataOut_payload_0_15482;
  reg        [7:0]    _zz_dataOut_payload_0_15483;
  wire                _zz_dataOut_payload_0_15484;
  wire       [7:0]    _zz_dataOut_payload_0_15485;
  wire       [7:0]    _zz_dataOut_payload_0_15486;
  wire                _zz_dataOut_payload_0_15487;
  wire       [7:0]    _zz_dataOut_payload_0_15488;
  wire       [7:0]    _zz_dataOut_payload_0_15489;
  wire                _zz_dataOut_payload_0_15490;
  wire                _zz_dataOut_payload_0_15491;
  reg        [7:0]    _zz_dataOut_payload_0_15492;
  reg        [7:0]    _zz_dataOut_payload_0_15493;
  reg        [7:0]    _zz_dataOut_payload_0_15494;
  reg        [7:0]    _zz_dataOut_payload_0_15495;
  reg        [7:0]    _zz_dataOut_payload_0_15496;
  reg        [7:0]    _zz_dataOut_payload_0_15497;
  reg        [7:0]    _zz_dataOut_payload_0_15498;
  reg        [7:0]    _zz_dataOut_payload_0_15499;
  reg        [7:0]    _zz_dataOut_payload_0_15500;
  reg        [7:0]    _zz_dataOut_payload_0_15501;
  reg        [7:0]    _zz_dataOut_payload_0_15502;
  reg        [7:0]    _zz_dataOut_payload_0_15503;
  reg        [7:0]    _zz_dataOut_payload_0_15504;
  reg        [7:0]    _zz_dataOut_payload_0_15505;
  reg        [7:0]    _zz_dataOut_payload_0_15506;
  reg        [7:0]    _zz_dataOut_payload_0_15507;
  reg        [7:0]    _zz_dataOut_payload_0_15508;
  reg        [7:0]    _zz_dataOut_payload_0_15509;
  reg        [7:0]    _zz_dataOut_payload_0_15510;
  reg        [7:0]    _zz_dataOut_payload_0_15511;
  reg        [7:0]    _zz_dataOut_payload_0_15512;
  reg        [7:0]    _zz_dataOut_payload_0_15513;
  reg        [7:0]    _zz_dataOut_payload_0_15514;
  reg        [7:0]    _zz_dataOut_payload_0_15515;
  reg        [7:0]    _zz_dataOut_payload_0_15516;
  reg        [7:0]    _zz_dataOut_payload_0_15517;
  reg        [7:0]    _zz_dataOut_payload_0_15518;
  reg        [7:0]    _zz_dataOut_payload_0_15519;
  wire                _zz_dataOut_payload_0_15520;
  wire       [7:0]    _zz_dataOut_payload_0_15521;
  wire       [7:0]    _zz_dataOut_payload_0_15522;
  wire                _zz_dataOut_payload_0_15523;
  wire       [7:0]    _zz_dataOut_payload_0_15524;
  wire       [7:0]    _zz_dataOut_payload_0_15525;
  wire                _zz_dataOut_payload_0_15526;
  wire       [7:0]    _zz_dataOut_payload_0_15527;
  wire       [7:0]    _zz_dataOut_payload_0_15528;
  wire                _zz_dataOut_payload_0_15529;
  wire       [7:0]    _zz_dataOut_payload_0_15530;
  wire       [7:0]    _zz_dataOut_payload_0_15531;
  wire                _zz_dataOut_payload_0_15532;
  wire       [7:0]    _zz_dataOut_payload_0_15533;
  wire       [7:0]    _zz_dataOut_payload_0_15534;
  wire                _zz_dataOut_payload_0_15535;
  wire       [7:0]    _zz_dataOut_payload_0_15536;
  wire       [7:0]    _zz_dataOut_payload_0_15537;
  wire                _zz_dataOut_payload_0_15538;
  wire       [7:0]    _zz_dataOut_payload_0_15539;
  wire       [7:0]    _zz_dataOut_payload_0_15540;
  wire                _zz_dataOut_payload_0_15541;
  wire       [7:0]    _zz_dataOut_payload_0_15542;
  wire       [7:0]    _zz_dataOut_payload_0_15543;
  wire                _zz_dataOut_payload_0_15544;
  wire       [7:0]    _zz_dataOut_payload_0_15545;
  wire       [7:0]    _zz_dataOut_payload_0_15546;
  wire                _zz_dataOut_payload_0_15547;
  wire       [7:0]    _zz_dataOut_payload_0_15548;
  wire       [7:0]    _zz_dataOut_payload_0_15549;
  wire                _zz_dataOut_payload_0_15550;
  wire       [7:0]    _zz_dataOut_payload_0_15551;
  wire       [7:0]    _zz_dataOut_payload_0_15552;
  wire                _zz_dataOut_payload_0_15553;
  wire       [7:0]    _zz_dataOut_payload_0_15554;
  wire       [7:0]    _zz_dataOut_payload_0_15555;
  wire                _zz_dataOut_payload_0_15556;
  wire       [7:0]    _zz_dataOut_payload_0_15557;
  wire       [7:0]    _zz_dataOut_payload_0_15558;
  wire                _zz_dataOut_payload_0_15559;
  wire       [7:0]    _zz_dataOut_payload_0_15560;
  wire       [7:0]    _zz_dataOut_payload_0_15561;
  wire                _zz_dataOut_payload_0_15562;
  wire                _zz_dataOut_payload_0_15563;
  reg        [7:0]    _zz_dataOut_payload_0_15564;
  reg        [7:0]    _zz_dataOut_payload_0_15565;
  reg        [7:0]    _zz_dataOut_payload_0_15566;
  reg        [7:0]    _zz_dataOut_payload_0_15567;
  wire                _zz_dataOut_payload_0_15568;
  wire       [7:0]    _zz_dataOut_payload_0_15569;
  wire       [7:0]    _zz_dataOut_payload_0_15570;
  wire                _zz_dataOut_payload_0_15571;
  wire       [7:0]    _zz_dataOut_payload_0_15572;
  wire       [7:0]    _zz_dataOut_payload_0_15573;
  wire                _zz_dataOut_payload_0_15574;
  wire                _zz_dataOut_payload_0_15575;
  reg        [7:0]    _zz_dataOut_payload_0_15576;
  reg        [7:0]    _zz_dataOut_payload_0_15577;
  reg        [7:0]    _zz_dataOut_payload_0_15578;
  reg        [7:0]    _zz_dataOut_payload_0_15579;
  reg        [7:0]    _zz_dataOut_payload_0_15580;
  reg        [7:0]    _zz_dataOut_payload_0_15581;
  reg        [7:0]    _zz_dataOut_payload_0_15582;
  reg        [7:0]    _zz_dataOut_payload_0_15583;
  reg        [7:0]    _zz_dataOut_payload_0_15584;
  reg        [7:0]    _zz_dataOut_payload_0_15585;
  reg        [7:0]    _zz_dataOut_payload_0_15586;
  reg        [7:0]    _zz_dataOut_payload_0_15587;
  wire                _zz_dataOut_payload_0_15588;
  wire       [7:0]    _zz_dataOut_payload_0_15589;
  wire       [7:0]    _zz_dataOut_payload_0_15590;
  wire                _zz_dataOut_payload_0_15591;
  wire       [7:0]    _zz_dataOut_payload_0_15592;
  wire       [7:0]    _zz_dataOut_payload_0_15593;
  wire                _zz_dataOut_payload_0_15594;
  wire       [7:0]    _zz_dataOut_payload_0_15595;
  wire       [7:0]    _zz_dataOut_payload_0_15596;
  wire                _zz_dataOut_payload_0_15597;
  wire       [7:0]    _zz_dataOut_payload_0_15598;
  wire       [7:0]    _zz_dataOut_payload_0_15599;
  wire                _zz_dataOut_payload_0_15600;
  wire       [7:0]    _zz_dataOut_payload_0_15601;
  wire       [7:0]    _zz_dataOut_payload_0_15602;
  wire                _zz_dataOut_payload_0_15603;
  wire       [7:0]    _zz_dataOut_payload_0_15604;
  wire       [7:0]    _zz_dataOut_payload_0_15605;
  wire                _zz_dataOut_payload_0_15606;
  wire                _zz_dataOut_payload_0_15607;
  reg        [7:0]    _zz_dataOut_payload_0_15608;
  reg        [7:0]    _zz_dataOut_payload_0_15609;
  reg        [7:0]    _zz_dataOut_payload_0_15610;
  reg        [7:0]    _zz_dataOut_payload_0_15611;
  wire                _zz_dataOut_payload_0_15612;
  wire       [7:0]    _zz_dataOut_payload_0_15613;
  wire       [7:0]    _zz_dataOut_payload_0_15614;
  wire                _zz_dataOut_payload_0_15615;
  wire       [7:0]    _zz_dataOut_payload_0_15616;
  wire       [7:0]    _zz_dataOut_payload_0_15617;
  wire                _zz_dataOut_payload_0_15618;
  wire                _zz_dataOut_payload_0_15619;
  reg        [7:0]    _zz_dataOut_payload_0_15620;
  reg        [7:0]    _zz_dataOut_payload_0_15621;
  reg        [7:0]    _zz_dataOut_payload_0_15622;
  reg        [7:0]    _zz_dataOut_payload_0_15623;
  reg        [7:0]    _zz_dataOut_payload_0_15624;
  reg        [7:0]    _zz_dataOut_payload_0_15625;
  reg        [7:0]    _zz_dataOut_payload_0_15626;
  reg        [7:0]    _zz_dataOut_payload_0_15627;
  reg        [7:0]    _zz_dataOut_payload_0_15628;
  reg        [7:0]    _zz_dataOut_payload_0_15629;
  reg        [7:0]    _zz_dataOut_payload_0_15630;
  reg        [7:0]    _zz_dataOut_payload_0_15631;
  reg        [7:0]    _zz_dataOut_payload_0_15632;
  reg        [7:0]    _zz_dataOut_payload_0_15633;
  reg        [7:0]    _zz_dataOut_payload_0_15634;
  reg        [7:0]    _zz_dataOut_payload_0_15635;
  reg        [7:0]    _zz_dataOut_payload_0_15636;
  reg        [7:0]    _zz_dataOut_payload_0_15637;
  reg        [7:0]    _zz_dataOut_payload_0_15638;
  reg        [7:0]    _zz_dataOut_payload_0_15639;
  reg        [7:0]    _zz_dataOut_payload_0_15640;
  reg        [7:0]    _zz_dataOut_payload_0_15641;
  reg        [7:0]    _zz_dataOut_payload_0_15642;
  reg        [7:0]    _zz_dataOut_payload_0_15643;
  reg        [7:0]    _zz_dataOut_payload_0_15644;
  reg        [7:0]    _zz_dataOut_payload_0_15645;
  reg        [7:0]    _zz_dataOut_payload_0_15646;
  reg        [7:0]    _zz_dataOut_payload_0_15647;
  reg        [7:0]    _zz_dataOut_payload_0_15648;
  reg        [7:0]    _zz_dataOut_payload_0_15649;
  reg        [7:0]    _zz_dataOut_payload_0_15650;
  reg        [7:0]    _zz_dataOut_payload_0_15651;
  reg        [7:0]    _zz_dataOut_payload_0_15652;
  reg        [7:0]    _zz_dataOut_payload_0_15653;
  reg        [7:0]    _zz_dataOut_payload_0_15654;
  reg        [7:0]    _zz_dataOut_payload_0_15655;
  reg        [7:0]    _zz_dataOut_payload_0_15656;
  reg        [7:0]    _zz_dataOut_payload_0_15657;
  reg        [7:0]    _zz_dataOut_payload_0_15658;
  reg        [7:0]    _zz_dataOut_payload_0_15659;
  reg        [7:0]    _zz_dataOut_payload_0_15660;
  reg        [7:0]    _zz_dataOut_payload_0_15661;
  reg        [7:0]    _zz_dataOut_payload_0_15662;
  reg        [7:0]    _zz_dataOut_payload_0_15663;
  reg        [7:0]    _zz_dataOut_payload_0_15664;
  reg        [7:0]    _zz_dataOut_payload_0_15665;
  reg        [7:0]    _zz_dataOut_payload_0_15666;
  reg        [7:0]    _zz_dataOut_payload_0_15667;
  reg        [7:0]    _zz_dataOut_payload_0_15668;
  reg        [7:0]    _zz_dataOut_payload_0_15669;
  reg        [7:0]    _zz_dataOut_payload_0_15670;
  reg        [7:0]    _zz_dataOut_payload_0_15671;
  reg        [7:0]    _zz_dataOut_payload_0_15672;
  reg        [7:0]    _zz_dataOut_payload_0_15673;
  reg        [7:0]    _zz_dataOut_payload_0_15674;
  reg        [7:0]    _zz_dataOut_payload_0_15675;
  reg        [7:0]    _zz_dataOut_payload_0_15676;
  reg        [7:0]    _zz_dataOut_payload_0_15677;
  reg        [7:0]    _zz_dataOut_payload_0_15678;
  reg        [7:0]    _zz_dataOut_payload_0_15679;
  reg        [7:0]    _zz_dataOut_payload_0_15680;
  reg        [7:0]    _zz_dataOut_payload_0_15681;
  reg        [7:0]    _zz_dataOut_payload_0_15682;
  reg        [7:0]    _zz_dataOut_payload_0_15683;
  reg        [7:0]    _zz_dataOut_payload_0_15684;
  reg        [7:0]    _zz_dataOut_payload_0_15685;
  reg        [7:0]    _zz_dataOut_payload_0_15686;
  reg        [7:0]    _zz_dataOut_payload_0_15687;
  reg        [7:0]    _zz_dataOut_payload_0_15688;
  reg        [7:0]    _zz_dataOut_payload_0_15689;
  reg        [7:0]    _zz_dataOut_payload_0_15690;
  reg        [7:0]    _zz_dataOut_payload_0_15691;
  reg        [7:0]    _zz_dataOut_payload_0_15692;
  reg        [7:0]    _zz_dataOut_payload_0_15693;
  reg        [7:0]    _zz_dataOut_payload_0_15694;
  reg        [7:0]    _zz_dataOut_payload_0_15695;
  reg        [7:0]    _zz_dataOut_payload_0_15696;
  reg        [7:0]    _zz_dataOut_payload_0_15697;
  reg        [7:0]    _zz_dataOut_payload_0_15698;
  reg        [7:0]    _zz_dataOut_payload_0_15699;
  reg        [7:0]    _zz_dataOut_payload_0_15700;
  reg        [7:0]    _zz_dataOut_payload_0_15701;
  reg        [7:0]    _zz_dataOut_payload_0_15702;
  reg        [7:0]    _zz_dataOut_payload_0_15703;
  reg        [7:0]    _zz_dataOut_payload_0_15704;
  reg        [7:0]    _zz_dataOut_payload_0_15705;
  reg        [7:0]    _zz_dataOut_payload_0_15706;
  reg        [7:0]    _zz_dataOut_payload_0_15707;
  reg        [7:0]    _zz_dataOut_payload_0_15708;
  reg        [7:0]    _zz_dataOut_payload_0_15709;
  reg        [7:0]    _zz_dataOut_payload_0_15710;
  reg        [7:0]    _zz_dataOut_payload_0_15711;
  reg        [7:0]    _zz_dataOut_payload_0_15712;
  reg        [7:0]    _zz_dataOut_payload_0_15713;
  reg        [7:0]    _zz_dataOut_payload_0_15714;
  reg        [7:0]    _zz_dataOut_payload_0_15715;
  reg        [7:0]    _zz_dataOut_payload_0_15716;
  reg        [7:0]    _zz_dataOut_payload_0_15717;
  reg        [7:0]    _zz_dataOut_payload_0_15718;
  reg        [7:0]    _zz_dataOut_payload_0_15719;
  reg        [7:0]    _zz_dataOut_payload_0_15720;
  reg        [7:0]    _zz_dataOut_payload_0_15721;
  reg        [7:0]    _zz_dataOut_payload_0_15722;
  reg        [7:0]    _zz_dataOut_payload_0_15723;
  reg        [7:0]    _zz_dataOut_payload_0_15724;
  reg        [7:0]    _zz_dataOut_payload_0_15725;
  reg        [7:0]    _zz_dataOut_payload_0_15726;
  reg        [7:0]    _zz_dataOut_payload_0_15727;
  reg        [7:0]    _zz_dataOut_payload_0_15728;
  reg        [7:0]    _zz_dataOut_payload_0_15729;
  reg        [7:0]    _zz_dataOut_payload_0_15730;
  reg        [7:0]    _zz_dataOut_payload_0_15731;
  reg        [7:0]    _zz_dataOut_payload_0_15732;
  reg        [7:0]    _zz_dataOut_payload_0_15733;
  reg        [7:0]    _zz_dataOut_payload_0_15734;
  reg        [7:0]    _zz_dataOut_payload_0_15735;
  reg        [7:0]    _zz_dataOut_payload_0_15736;
  reg        [7:0]    _zz_dataOut_payload_0_15737;
  reg        [7:0]    _zz_dataOut_payload_0_15738;
  reg        [7:0]    _zz_dataOut_payload_0_15739;
  reg        [7:0]    _zz_dataOut_payload_0_15740;
  reg        [7:0]    _zz_dataOut_payload_0_15741;
  reg        [7:0]    _zz_dataOut_payload_0_15742;
  reg        [7:0]    _zz_dataOut_payload_0_15743;
  reg        [7:0]    _zz_dataOut_payload_0_15744;
  reg        [7:0]    _zz_dataOut_payload_0_15745;
  reg        [7:0]    _zz_dataOut_payload_0_15746;
  reg        [7:0]    _zz_dataOut_payload_0_15747;
  reg        [7:0]    _zz_dataOut_payload_0_15748;
  reg        [7:0]    _zz_dataOut_payload_0_15749;
  reg        [7:0]    _zz_dataOut_payload_0_15750;
  reg        [7:0]    _zz_dataOut_payload_0_15751;
  reg        [7:0]    _zz_dataOut_payload_0_15752;
  reg        [7:0]    _zz_dataOut_payload_0_15753;
  reg        [7:0]    _zz_dataOut_payload_0_15754;
  reg        [7:0]    _zz_dataOut_payload_0_15755;
  reg        [7:0]    _zz_dataOut_payload_0_15756;
  reg        [7:0]    _zz_dataOut_payload_0_15757;
  reg        [7:0]    _zz_dataOut_payload_0_15758;
  reg        [7:0]    _zz_dataOut_payload_0_15759;
  reg        [7:0]    _zz_dataOut_payload_0_15760;
  reg        [7:0]    _zz_dataOut_payload_0_15761;
  reg        [7:0]    _zz_dataOut_payload_0_15762;
  reg        [7:0]    _zz_dataOut_payload_0_15763;
  reg        [7:0]    _zz_dataOut_payload_0_15764;
  reg        [7:0]    _zz_dataOut_payload_0_15765;
  reg        [7:0]    _zz_dataOut_payload_0_15766;
  reg        [7:0]    _zz_dataOut_payload_0_15767;
  reg        [7:0]    _zz_dataOut_payload_0_15768;
  reg        [7:0]    _zz_dataOut_payload_0_15769;
  reg        [7:0]    _zz_dataOut_payload_0_15770;
  reg        [7:0]    _zz_dataOut_payload_0_15771;
  reg        [7:0]    _zz_dataOut_payload_0_15772;
  reg        [7:0]    _zz_dataOut_payload_0_15773;
  reg        [7:0]    _zz_dataOut_payload_0_15774;
  reg        [7:0]    _zz_dataOut_payload_0_15775;
  reg        [7:0]    _zz_dataOut_payload_0_15776;
  reg        [7:0]    _zz_dataOut_payload_0_15777;
  reg        [7:0]    _zz_dataOut_payload_0_15778;
  reg        [7:0]    _zz_dataOut_payload_0_15779;
  reg        [7:0]    _zz_dataOut_payload_0_15780;
  reg        [7:0]    _zz_dataOut_payload_0_15781;
  reg        [7:0]    _zz_dataOut_payload_0_15782;
  reg        [7:0]    _zz_dataOut_payload_0_15783;
  reg        [7:0]    _zz_dataOut_payload_0_15784;
  reg        [7:0]    _zz_dataOut_payload_0_15785;
  reg        [7:0]    _zz_dataOut_payload_0_15786;
  reg        [7:0]    _zz_dataOut_payload_0_15787;
  reg        [7:0]    _zz_dataOut_payload_0_15788;
  reg        [7:0]    _zz_dataOut_payload_0_15789;
  reg        [7:0]    _zz_dataOut_payload_0_15790;
  reg        [7:0]    _zz_dataOut_payload_0_15791;
  reg        [7:0]    _zz_dataOut_payload_0_15792;
  reg        [7:0]    _zz_dataOut_payload_0_15793;
  reg        [7:0]    _zz_dataOut_payload_0_15794;
  reg        [7:0]    _zz_dataOut_payload_0_15795;
  reg        [7:0]    _zz_dataOut_payload_0_15796;
  reg        [7:0]    _zz_dataOut_payload_0_15797;
  reg        [7:0]    _zz_dataOut_payload_0_15798;
  reg        [7:0]    _zz_dataOut_payload_0_15799;
  reg        [7:0]    _zz_dataOut_payload_0_15800;
  reg        [7:0]    _zz_dataOut_payload_0_15801;
  reg        [7:0]    _zz_dataOut_payload_0_15802;
  reg        [7:0]    _zz_dataOut_payload_0_15803;
  reg        [7:0]    _zz_dataOut_payload_0_15804;
  reg        [7:0]    _zz_dataOut_payload_0_15805;
  reg        [7:0]    _zz_dataOut_payload_0_15806;
  reg        [7:0]    _zz_dataOut_payload_0_15807;
  reg        [7:0]    _zz_dataOut_payload_0_15808;
  reg        [7:0]    _zz_dataOut_payload_0_15809;
  reg        [7:0]    _zz_dataOut_payload_0_15810;
  reg        [7:0]    _zz_dataOut_payload_0_15811;
  reg        [7:0]    _zz_dataOut_payload_0_15812;
  reg        [7:0]    _zz_dataOut_payload_0_15813;
  reg        [7:0]    _zz_dataOut_payload_0_15814;
  reg        [7:0]    _zz_dataOut_payload_0_15815;
  reg        [7:0]    _zz_dataOut_payload_0_15816;
  reg        [7:0]    _zz_dataOut_payload_0_15817;
  reg        [7:0]    _zz_dataOut_payload_0_15818;
  reg        [7:0]    _zz_dataOut_payload_0_15819;
  reg        [7:0]    _zz_dataOut_payload_0_15820;
  reg        [7:0]    _zz_dataOut_payload_0_15821;
  reg        [7:0]    _zz_dataOut_payload_0_15822;
  reg        [7:0]    _zz_dataOut_payload_0_15823;
  reg        [7:0]    _zz_dataOut_payload_0_15824;
  reg        [7:0]    _zz_dataOut_payload_0_15825;
  reg        [7:0]    _zz_dataOut_payload_0_15826;
  reg        [7:0]    _zz_dataOut_payload_0_15827;
  reg        [7:0]    _zz_dataOut_payload_0_15828;
  reg        [7:0]    _zz_dataOut_payload_0_15829;
  reg        [7:0]    _zz_dataOut_payload_0_15830;
  reg        [7:0]    _zz_dataOut_payload_0_15831;
  reg        [7:0]    _zz_dataOut_payload_0_15832;
  reg        [7:0]    _zz_dataOut_payload_0_15833;
  reg        [7:0]    _zz_dataOut_payload_0_15834;
  reg        [7:0]    _zz_dataOut_payload_0_15835;
  reg        [7:0]    _zz_dataOut_payload_0_15836;
  reg        [7:0]    _zz_dataOut_payload_0_15837;
  reg        [7:0]    _zz_dataOut_payload_0_15838;
  reg        [7:0]    _zz_dataOut_payload_0_15839;
  reg        [7:0]    _zz_dataOut_payload_0_15840;
  reg        [7:0]    _zz_dataOut_payload_0_15841;
  reg        [7:0]    _zz_dataOut_payload_0_15842;
  reg        [7:0]    _zz_dataOut_payload_0_15843;
  reg        [7:0]    _zz_dataOut_payload_0_15844;
  reg        [7:0]    _zz_dataOut_payload_0_15845;
  reg        [7:0]    _zz_dataOut_payload_0_15846;
  reg        [7:0]    _zz_dataOut_payload_0_15847;
  reg        [7:0]    _zz_dataOut_payload_0_15848;
  reg        [7:0]    _zz_dataOut_payload_0_15849;
  reg        [7:0]    _zz_dataOut_payload_0_15850;
  reg        [7:0]    _zz_dataOut_payload_0_15851;
  reg        [7:0]    _zz_dataOut_payload_0_15852;
  reg        [7:0]    _zz_dataOut_payload_0_15853;
  reg        [7:0]    _zz_dataOut_payload_0_15854;
  reg        [7:0]    _zz_dataOut_payload_0_15855;
  reg        [7:0]    _zz_dataOut_payload_0_15856;
  reg        [7:0]    _zz_dataOut_payload_0_15857;
  reg        [7:0]    _zz_dataOut_payload_0_15858;
  reg        [7:0]    _zz_dataOut_payload_0_15859;
  reg        [7:0]    _zz_dataOut_payload_0_15860;
  reg        [7:0]    _zz_dataOut_payload_0_15861;
  reg        [7:0]    _zz_dataOut_payload_0_15862;
  reg        [7:0]    _zz_dataOut_payload_0_15863;
  reg        [7:0]    _zz_dataOut_payload_0_15864;
  reg        [7:0]    _zz_dataOut_payload_0_15865;
  reg        [7:0]    _zz_dataOut_payload_0_15866;
  reg        [7:0]    _zz_dataOut_payload_0_15867;
  reg        [7:0]    _zz_dataOut_payload_0_15868;
  reg        [7:0]    _zz_dataOut_payload_0_15869;
  reg        [7:0]    _zz_dataOut_payload_0_15870;
  reg        [7:0]    _zz_dataOut_payload_0_15871;
  reg        [7:0]    _zz_dataOut_payload_0_15872;
  reg        [7:0]    _zz_dataOut_payload_0_15873;
  reg        [7:0]    _zz_dataOut_payload_0_15874;
  reg        [7:0]    _zz_dataOut_payload_0_15875;
  reg        [7:0]    _zz_dataOut_payload_0_15876;
  reg        [7:0]    _zz_dataOut_payload_0_15877;
  reg        [7:0]    _zz_dataOut_payload_0_15878;
  reg        [7:0]    _zz_dataOut_payload_0_15879;
  reg        [7:0]    _zz_dataOut_payload_0_15880;
  reg        [7:0]    _zz_dataOut_payload_0_15881;
  reg        [7:0]    _zz_dataOut_payload_0_15882;
  reg        [7:0]    _zz_dataOut_payload_0_15883;
  reg        [7:0]    _zz_dataOut_payload_0_15884;
  reg        [7:0]    _zz_dataOut_payload_0_15885;
  reg        [7:0]    _zz_dataOut_payload_0_15886;
  reg        [7:0]    _zz_dataOut_payload_0_15887;
  reg        [7:0]    _zz_dataOut_payload_0_15888;
  reg        [7:0]    _zz_dataOut_payload_0_15889;
  reg        [7:0]    _zz_dataOut_payload_0_15890;
  reg        [7:0]    _zz_dataOut_payload_0_15891;
  reg        [7:0]    _zz_dataOut_payload_0_15892;
  reg        [7:0]    _zz_dataOut_payload_0_15893;
  reg        [7:0]    _zz_dataOut_payload_0_15894;
  reg        [7:0]    _zz_dataOut_payload_0_15895;
  reg        [7:0]    _zz_dataOut_payload_0_15896;
  reg        [7:0]    _zz_dataOut_payload_0_15897;
  reg        [7:0]    _zz_dataOut_payload_0_15898;
  reg        [7:0]    _zz_dataOut_payload_0_15899;
  reg        [7:0]    _zz_dataOut_payload_0_15900;
  reg        [7:0]    _zz_dataOut_payload_0_15901;
  reg        [7:0]    _zz_dataOut_payload_0_15902;
  reg        [7:0]    _zz_dataOut_payload_0_15903;
  reg        [7:0]    _zz_dataOut_payload_0_15904;
  reg        [7:0]    _zz_dataOut_payload_0_15905;
  reg        [7:0]    _zz_dataOut_payload_0_15906;
  reg        [7:0]    _zz_dataOut_payload_0_15907;
  reg        [7:0]    _zz_dataOut_payload_0_15908;
  reg        [7:0]    _zz_dataOut_payload_0_15909;
  reg        [7:0]    _zz_dataOut_payload_0_15910;
  reg        [7:0]    _zz_dataOut_payload_0_15911;
  reg        [7:0]    _zz_dataOut_payload_0_15912;
  reg        [7:0]    _zz_dataOut_payload_0_15913;
  reg        [7:0]    _zz_dataOut_payload_0_15914;
  reg        [7:0]    _zz_dataOut_payload_0_15915;
  reg        [7:0]    _zz_dataOut_payload_0_15916;
  reg        [7:0]    _zz_dataOut_payload_0_15917;
  reg        [7:0]    _zz_dataOut_payload_0_15918;
  reg        [7:0]    _zz_dataOut_payload_0_15919;
  reg        [7:0]    _zz_dataOut_payload_0_15920;
  reg        [7:0]    _zz_dataOut_payload_0_15921;
  reg        [7:0]    _zz_dataOut_payload_0_15922;
  reg        [7:0]    _zz_dataOut_payload_0_15923;
  reg        [7:0]    _zz_dataOut_payload_0_15924;
  reg        [7:0]    _zz_dataOut_payload_0_15925;
  reg        [7:0]    _zz_dataOut_payload_0_15926;
  reg        [7:0]    _zz_dataOut_payload_0_15927;
  reg        [7:0]    _zz_dataOut_payload_0_15928;
  reg        [7:0]    _zz_dataOut_payload_0_15929;
  reg        [7:0]    _zz_dataOut_payload_0_15930;
  reg        [7:0]    _zz_dataOut_payload_0_15931;
  reg        [7:0]    _zz_dataOut_payload_0_15932;
  reg        [7:0]    _zz_dataOut_payload_0_15933;
  reg        [7:0]    _zz_dataOut_payload_0_15934;
  reg        [7:0]    _zz_dataOut_payload_0_15935;
  reg        [7:0]    _zz_dataOut_payload_0_15936;
  reg        [7:0]    _zz_dataOut_payload_0_15937;
  reg        [7:0]    _zz_dataOut_payload_0_15938;
  reg        [7:0]    _zz_dataOut_payload_0_15939;
  reg        [7:0]    _zz_dataOut_payload_0_15940;
  reg        [7:0]    _zz_dataOut_payload_0_15941;
  reg        [7:0]    _zz_dataOut_payload_0_15942;
  reg        [7:0]    _zz_dataOut_payload_0_15943;
  reg        [7:0]    _zz_dataOut_payload_0_15944;
  reg        [7:0]    _zz_dataOut_payload_0_15945;
  reg        [7:0]    _zz_dataOut_payload_0_15946;
  reg        [7:0]    _zz_dataOut_payload_0_15947;
  reg        [7:0]    _zz_dataOut_payload_0_15948;
  reg        [7:0]    _zz_dataOut_payload_0_15949;
  reg        [7:0]    _zz_dataOut_payload_0_15950;
  reg        [7:0]    _zz_dataOut_payload_0_15951;
  reg        [7:0]    _zz_dataOut_payload_0_15952;
  reg        [7:0]    _zz_dataOut_payload_0_15953;
  reg        [7:0]    _zz_dataOut_payload_0_15954;
  reg        [7:0]    _zz_dataOut_payload_0_15955;
  reg        [7:0]    _zz_dataOut_payload_0_15956;
  reg        [7:0]    _zz_dataOut_payload_0_15957;
  reg        [7:0]    _zz_dataOut_payload_0_15958;
  reg        [7:0]    _zz_dataOut_payload_0_15959;
  reg        [7:0]    _zz_dataOut_payload_0_15960;
  reg        [7:0]    _zz_dataOut_payload_0_15961;
  reg        [7:0]    _zz_dataOut_payload_0_15962;
  reg        [7:0]    _zz_dataOut_payload_0_15963;
  reg        [7:0]    _zz_dataOut_payload_0_15964;
  reg        [7:0]    _zz_dataOut_payload_0_15965;
  reg        [7:0]    _zz_dataOut_payload_0_15966;
  reg        [7:0]    _zz_dataOut_payload_0_15967;
  reg        [7:0]    _zz_dataOut_payload_0_15968;
  reg        [7:0]    _zz_dataOut_payload_0_15969;
  reg        [7:0]    _zz_dataOut_payload_0_15970;
  reg        [7:0]    _zz_dataOut_payload_0_15971;
  reg        [7:0]    _zz_dataOut_payload_0_15972;
  reg        [7:0]    _zz_dataOut_payload_0_15973;
  reg        [7:0]    _zz_dataOut_payload_0_15974;
  reg        [7:0]    _zz_dataOut_payload_0_15975;
  reg        [7:0]    _zz_dataOut_payload_0_15976;
  reg        [7:0]    _zz_dataOut_payload_0_15977;
  reg        [7:0]    _zz_dataOut_payload_0_15978;
  reg        [7:0]    _zz_dataOut_payload_0_15979;
  reg        [7:0]    _zz_dataOut_payload_0_15980;
  reg        [7:0]    _zz_dataOut_payload_0_15981;
  reg        [7:0]    _zz_dataOut_payload_0_15982;
  reg        [7:0]    _zz_dataOut_payload_0_15983;
  reg        [7:0]    _zz_dataOut_payload_0_15984;
  reg        [7:0]    _zz_dataOut_payload_0_15985;
  reg        [7:0]    _zz_dataOut_payload_0_15986;
  reg        [7:0]    _zz_dataOut_payload_0_15987;
  reg        [7:0]    _zz_dataOut_payload_0_15988;
  reg        [7:0]    _zz_dataOut_payload_0_15989;
  reg        [7:0]    _zz_dataOut_payload_0_15990;
  reg        [7:0]    _zz_dataOut_payload_0_15991;
  reg        [7:0]    _zz_dataOut_payload_0_15992;
  reg        [7:0]    _zz_dataOut_payload_0_15993;
  reg        [7:0]    _zz_dataOut_payload_0_15994;
  reg        [7:0]    _zz_dataOut_payload_0_15995;
  reg        [7:0]    _zz_dataOut_payload_0_15996;
  reg        [7:0]    _zz_dataOut_payload_0_15997;
  reg        [7:0]    _zz_dataOut_payload_0_15998;
  reg        [7:0]    _zz_dataOut_payload_0_15999;
  reg        [7:0]    _zz_dataOut_payload_0_16000;
  reg        [7:0]    _zz_dataOut_payload_0_16001;
  reg        [7:0]    _zz_dataOut_payload_0_16002;
  reg        [7:0]    _zz_dataOut_payload_0_16003;
  reg        [7:0]    _zz_dataOut_payload_0_16004;
  reg        [7:0]    _zz_dataOut_payload_0_16005;
  reg        [7:0]    _zz_dataOut_payload_0_16006;
  reg        [7:0]    _zz_dataOut_payload_0_16007;
  reg        [7:0]    _zz_dataOut_payload_0_16008;
  reg        [7:0]    _zz_dataOut_payload_0_16009;
  reg        [7:0]    _zz_dataOut_payload_0_16010;
  reg        [7:0]    _zz_dataOut_payload_0_16011;
  reg        [7:0]    _zz_dataOut_payload_0_16012;
  reg        [7:0]    _zz_dataOut_payload_0_16013;
  reg        [7:0]    _zz_dataOut_payload_0_16014;
  reg        [7:0]    _zz_dataOut_payload_0_16015;
  reg        [7:0]    _zz_dataOut_payload_0_16016;
  reg        [7:0]    _zz_dataOut_payload_0_16017;
  reg        [7:0]    _zz_dataOut_payload_0_16018;
  reg        [7:0]    _zz_dataOut_payload_0_16019;
  reg        [7:0]    _zz_dataOut_payload_0_16020;
  reg        [7:0]    _zz_dataOut_payload_0_16021;
  reg        [7:0]    _zz_dataOut_payload_0_16022;
  reg        [7:0]    _zz_dataOut_payload_0_16023;
  reg        [7:0]    _zz_dataOut_payload_0_16024;
  reg        [7:0]    _zz_dataOut_payload_0_16025;
  reg        [7:0]    _zz_dataOut_payload_0_16026;
  reg        [7:0]    _zz_dataOut_payload_0_16027;
  reg        [7:0]    _zz_dataOut_payload_0_16028;
  reg        [7:0]    _zz_dataOut_payload_0_16029;
  reg        [7:0]    _zz_dataOut_payload_0_16030;
  reg        [7:0]    _zz_dataOut_payload_0_16031;
  reg        [7:0]    _zz_dataOut_payload_0_16032;
  reg        [7:0]    _zz_dataOut_payload_0_16033;
  reg        [7:0]    _zz_dataOut_payload_0_16034;
  reg        [7:0]    _zz_dataOut_payload_0_16035;
  reg        [7:0]    _zz_dataOut_payload_0_16036;
  reg        [7:0]    _zz_dataOut_payload_0_16037;
  reg        [7:0]    _zz_dataOut_payload_0_16038;
  reg        [7:0]    _zz_dataOut_payload_0_16039;
  reg        [7:0]    _zz_dataOut_payload_0_16040;
  reg        [7:0]    _zz_dataOut_payload_0_16041;
  reg        [7:0]    _zz_dataOut_payload_0_16042;
  reg        [7:0]    _zz_dataOut_payload_0_16043;
  reg        [7:0]    _zz_dataOut_payload_0_16044;
  reg        [7:0]    _zz_dataOut_payload_0_16045;
  reg        [7:0]    _zz_dataOut_payload_0_16046;
  reg        [7:0]    _zz_dataOut_payload_0_16047;
  reg        [7:0]    _zz_dataOut_payload_0_16048;
  reg        [7:0]    _zz_dataOut_payload_0_16049;
  reg        [7:0]    _zz_dataOut_payload_0_16050;
  reg        [7:0]    _zz_dataOut_payload_0_16051;
  reg        [7:0]    _zz_dataOut_payload_0_16052;
  reg        [7:0]    _zz_dataOut_payload_0_16053;
  reg        [7:0]    _zz_dataOut_payload_0_16054;
  reg        [7:0]    _zz_dataOut_payload_0_16055;
  reg        [7:0]    _zz_dataOut_payload_0_16056;
  reg        [7:0]    _zz_dataOut_payload_0_16057;
  reg        [7:0]    _zz_dataOut_payload_0_16058;
  reg        [7:0]    _zz_dataOut_payload_0_16059;
  reg        [7:0]    _zz_dataOut_payload_0_16060;
  reg        [7:0]    _zz_dataOut_payload_0_16061;
  reg        [7:0]    _zz_dataOut_payload_0_16062;
  reg        [7:0]    _zz_dataOut_payload_0_16063;
  reg        [7:0]    _zz_dataOut_payload_0_16064;
  reg        [7:0]    _zz_dataOut_payload_0_16065;
  reg        [7:0]    _zz_dataOut_payload_0_16066;
  reg        [7:0]    _zz_dataOut_payload_0_16067;
  reg        [7:0]    _zz_dataOut_payload_0_16068;
  reg        [7:0]    _zz_dataOut_payload_0_16069;
  reg        [7:0]    _zz_dataOut_payload_0_16070;
  reg        [7:0]    _zz_dataOut_payload_0_16071;
  reg        [7:0]    _zz_dataOut_payload_0_16072;
  reg        [7:0]    _zz_dataOut_payload_0_16073;
  reg        [7:0]    _zz_dataOut_payload_0_16074;
  reg        [7:0]    _zz_dataOut_payload_0_16075;
  reg        [7:0]    _zz_dataOut_payload_0_16076;
  reg        [7:0]    _zz_dataOut_payload_0_16077;
  reg        [7:0]    _zz_dataOut_payload_0_16078;
  reg        [7:0]    _zz_dataOut_payload_0_16079;
  reg        [7:0]    _zz_dataOut_payload_0_16080;
  reg        [7:0]    _zz_dataOut_payload_0_16081;
  reg        [7:0]    _zz_dataOut_payload_0_16082;
  reg        [7:0]    _zz_dataOut_payload_0_16083;
  reg        [7:0]    _zz_dataOut_payload_0_16084;
  reg        [7:0]    _zz_dataOut_payload_0_16085;
  reg        [7:0]    _zz_dataOut_payload_0_16086;
  reg        [7:0]    _zz_dataOut_payload_0_16087;
  reg        [7:0]    _zz_dataOut_payload_0_16088;
  reg        [7:0]    _zz_dataOut_payload_0_16089;
  reg        [7:0]    _zz_dataOut_payload_0_16090;
  reg        [7:0]    _zz_dataOut_payload_0_16091;
  reg        [7:0]    _zz_dataOut_payload_0_16092;
  reg        [7:0]    _zz_dataOut_payload_0_16093;
  reg        [7:0]    _zz_dataOut_payload_0_16094;
  reg        [7:0]    _zz_dataOut_payload_0_16095;
  reg        [7:0]    _zz_dataOut_payload_0_16096;
  reg        [7:0]    _zz_dataOut_payload_0_16097;
  reg        [7:0]    _zz_dataOut_payload_0_16098;
  reg        [7:0]    _zz_dataOut_payload_0_16099;
  reg        [7:0]    _zz_dataOut_payload_0_16100;
  reg        [7:0]    _zz_dataOut_payload_0_16101;
  reg        [7:0]    _zz_dataOut_payload_0_16102;
  reg        [7:0]    _zz_dataOut_payload_0_16103;
  reg        [7:0]    _zz_dataOut_payload_0_16104;
  reg        [7:0]    _zz_dataOut_payload_0_16105;
  reg        [7:0]    _zz_dataOut_payload_0_16106;
  reg        [7:0]    _zz_dataOut_payload_0_16107;
  reg        [7:0]    _zz_dataOut_payload_0_16108;
  reg        [7:0]    _zz_dataOut_payload_0_16109;
  reg        [7:0]    _zz_dataOut_payload_0_16110;
  reg        [7:0]    _zz_dataOut_payload_0_16111;
  reg        [7:0]    _zz_dataOut_payload_0_16112;
  reg        [7:0]    _zz_dataOut_payload_0_16113;
  reg        [7:0]    _zz_dataOut_payload_0_16114;
  reg        [7:0]    _zz_dataOut_payload_0_16115;
  reg        [7:0]    _zz_dataOut_payload_0_16116;
  reg        [7:0]    _zz_dataOut_payload_0_16117;
  reg        [7:0]    _zz_dataOut_payload_0_16118;
  reg        [7:0]    _zz_dataOut_payload_0_16119;
  reg        [7:0]    _zz_dataOut_payload_0_16120;
  reg        [7:0]    _zz_dataOut_payload_0_16121;
  reg        [7:0]    _zz_dataOut_payload_0_16122;
  reg        [7:0]    _zz_dataOut_payload_0_16123;
  reg        [7:0]    _zz_dataOut_payload_0_16124;
  reg        [7:0]    _zz_dataOut_payload_0_16125;
  reg        [7:0]    _zz_dataOut_payload_0_16126;
  reg        [7:0]    _zz_dataOut_payload_0_16127;
  wire                _zz_dataOut_payload_0_16128;
  wire       [7:0]    _zz_dataOut_payload_0_16129;
  wire       [7:0]    _zz_dataOut_payload_128;
  wire                _zz_dataOut_payload_0_16130;
  wire       [7:0]    _zz_dataOut_payload_0_16131;
  wire       [7:0]    _zz_dataOut_payload_128_1;
  wire                _zz_dataOut_payload_0_16132;
  wire       [7:0]    _zz_dataOut_payload_0_16133;
  wire       [7:0]    _zz_dataOut_payload_128_2;
  wire                _zz_dataOut_payload_0_16134;
  wire       [7:0]    _zz_dataOut_payload_0_16135;
  wire       [7:0]    _zz_dataOut_payload_128_3;
  wire                _zz_dataOut_payload_0_16136;
  wire       [7:0]    _zz_dataOut_payload_0_16137;
  wire       [7:0]    _zz_dataOut_payload_128_4;
  wire                _zz_dataOut_payload_0_16138;
  wire       [7:0]    _zz_dataOut_payload_0_16139;
  wire       [7:0]    _zz_dataOut_payload_128_5;
  wire                _zz_dataOut_payload_0_16140;
  wire       [7:0]    _zz_dataOut_payload_0_16141;
  wire       [7:0]    _zz_dataOut_payload_128_6;
  wire                _zz_dataOut_payload_0_16142;
  wire       [7:0]    _zz_dataOut_payload_0_16143;
  wire       [7:0]    _zz_dataOut_payload_128_7;
  wire                _zz_dataOut_payload_0_16144;
  wire       [7:0]    _zz_dataOut_payload_0_16145;
  wire       [7:0]    _zz_dataOut_payload_128_8;
  wire                _zz_dataOut_payload_0_16146;
  wire       [7:0]    _zz_dataOut_payload_0_16147;
  wire       [7:0]    _zz_dataOut_payload_128_9;
  wire                _zz_dataOut_payload_0_16148;
  wire       [7:0]    _zz_dataOut_payload_0_16149;
  wire       [7:0]    _zz_dataOut_payload_128_10;
  wire                _zz_dataOut_payload_0_16150;
  wire       [7:0]    _zz_dataOut_payload_0_16151;
  wire       [7:0]    _zz_dataOut_payload_128_11;
  wire                _zz_dataOut_payload_0_16152;
  wire       [7:0]    _zz_dataOut_payload_0_16153;
  wire       [7:0]    _zz_dataOut_payload_128_12;
  wire                _zz_dataOut_payload_0_16154;
  wire       [7:0]    _zz_dataOut_payload_0_16155;
  wire       [7:0]    _zz_dataOut_payload_128_13;
  wire                _zz_dataOut_payload_0_16156;
  wire       [7:0]    _zz_dataOut_payload_0_16157;
  wire       [7:0]    _zz_dataOut_payload_128_14;
  wire                _zz_dataOut_payload_0_16158;
  wire       [7:0]    _zz_dataOut_payload_0_16159;
  wire       [7:0]    _zz_dataOut_payload_128_15;
  wire                _zz_dataOut_payload_0_16160;
  wire       [7:0]    _zz_dataOut_payload_0_16161;
  wire       [7:0]    _zz_dataOut_payload_128_16;
  wire                _zz_dataOut_payload_0_16162;
  wire       [7:0]    _zz_dataOut_payload_0_16163;
  wire       [7:0]    _zz_dataOut_payload_128_17;
  wire                _zz_dataOut_payload_0_16164;
  wire       [7:0]    _zz_dataOut_payload_0_16165;
  wire       [7:0]    _zz_dataOut_payload_128_18;
  wire                _zz_dataOut_payload_0_16166;
  wire       [7:0]    _zz_dataOut_payload_0_16167;
  wire       [7:0]    _zz_dataOut_payload_128_19;
  wire                _zz_dataOut_payload_0_16168;
  wire       [7:0]    _zz_dataOut_payload_0_16169;
  wire       [7:0]    _zz_dataOut_payload_128_20;
  wire                _zz_dataOut_payload_0_16170;
  wire       [7:0]    _zz_dataOut_payload_0_16171;
  wire       [7:0]    _zz_dataOut_payload_128_21;
  wire                _zz_dataOut_payload_0_16172;
  wire       [7:0]    _zz_dataOut_payload_0_16173;
  wire       [7:0]    _zz_dataOut_payload_128_22;
  wire                _zz_dataOut_payload_0_16174;
  wire       [7:0]    _zz_dataOut_payload_0_16175;
  wire       [7:0]    _zz_dataOut_payload_128_23;
  wire                _zz_dataOut_payload_0_16176;
  wire       [7:0]    _zz_dataOut_payload_0_16177;
  wire       [7:0]    _zz_dataOut_payload_128_24;
  wire                _zz_dataOut_payload_0_16178;
  wire       [7:0]    _zz_dataOut_payload_0_16179;
  wire       [7:0]    _zz_dataOut_payload_128_25;
  wire                _zz_dataOut_payload_0_16180;
  wire       [7:0]    _zz_dataOut_payload_0_16181;
  wire       [7:0]    _zz_dataOut_payload_128_26;
  wire                _zz_dataOut_payload_0_16182;
  wire       [7:0]    _zz_dataOut_payload_0_16183;
  wire       [7:0]    _zz_dataOut_payload_128_27;
  wire                _zz_dataOut_payload_0_16184;
  wire       [7:0]    _zz_dataOut_payload_0_16185;
  wire       [7:0]    _zz_dataOut_payload_128_28;
  wire                _zz_dataOut_payload_0_16186;
  wire       [7:0]    _zz_dataOut_payload_0_16187;
  wire       [7:0]    _zz_dataOut_payload_128_29;
  wire                _zz_dataOut_payload_0_16188;
  wire       [7:0]    _zz_dataOut_payload_0_16189;
  wire       [7:0]    _zz_dataOut_payload_128_30;
  wire                _zz_dataOut_payload_0_16190;
  wire       [7:0]    _zz_dataOut_payload_0_16191;
  wire       [7:0]    _zz_dataOut_payload_128_31;
  wire                _zz_dataOut_payload_0_16192;
  wire       [7:0]    _zz_dataOut_payload_0_16193;
  wire       [7:0]    _zz_dataOut_payload_128_32;
  wire                _zz_dataOut_payload_0_16194;
  wire       [7:0]    _zz_dataOut_payload_0_16195;
  wire       [7:0]    _zz_dataOut_payload_128_33;
  wire                _zz_dataOut_payload_0_16196;
  wire       [7:0]    _zz_dataOut_payload_0_16197;
  wire       [7:0]    _zz_dataOut_payload_128_34;
  wire                _zz_dataOut_payload_0_16198;
  wire       [7:0]    _zz_dataOut_payload_0_16199;
  wire       [7:0]    _zz_dataOut_payload_128_35;
  wire                _zz_dataOut_payload_0_16200;
  wire       [7:0]    _zz_dataOut_payload_0_16201;
  wire       [7:0]    _zz_dataOut_payload_128_36;
  wire                _zz_dataOut_payload_0_16202;
  wire       [7:0]    _zz_dataOut_payload_0_16203;
  wire       [7:0]    _zz_dataOut_payload_128_37;
  wire                _zz_dataOut_payload_0_16204;
  wire       [7:0]    _zz_dataOut_payload_0_16205;
  wire       [7:0]    _zz_dataOut_payload_128_38;
  wire                _zz_dataOut_payload_0_16206;
  wire       [7:0]    _zz_dataOut_payload_0_16207;
  wire       [7:0]    _zz_dataOut_payload_128_39;
  wire                _zz_dataOut_payload_0_16208;
  wire       [7:0]    _zz_dataOut_payload_0_16209;
  wire       [7:0]    _zz_dataOut_payload_128_40;
  wire                _zz_dataOut_payload_0_16210;
  wire       [7:0]    _zz_dataOut_payload_0_16211;
  wire       [7:0]    _zz_dataOut_payload_128_41;
  wire                _zz_dataOut_payload_0_16212;
  wire       [7:0]    _zz_dataOut_payload_0_16213;
  wire       [7:0]    _zz_dataOut_payload_128_42;
  wire                _zz_dataOut_payload_0_16214;
  wire       [7:0]    _zz_dataOut_payload_0_16215;
  wire       [7:0]    _zz_dataOut_payload_128_43;
  wire                _zz_dataOut_payload_0_16216;
  wire       [7:0]    _zz_dataOut_payload_0_16217;
  wire       [7:0]    _zz_dataOut_payload_128_44;
  wire                _zz_dataOut_payload_0_16218;
  wire       [7:0]    _zz_dataOut_payload_0_16219;
  wire       [7:0]    _zz_dataOut_payload_128_45;
  wire                _zz_dataOut_payload_0_16220;
  wire       [7:0]    _zz_dataOut_payload_0_16221;
  wire       [7:0]    _zz_dataOut_payload_128_46;
  wire                _zz_dataOut_payload_0_16222;
  wire       [7:0]    _zz_dataOut_payload_0_16223;
  wire       [7:0]    _zz_dataOut_payload_128_47;
  wire                _zz_dataOut_payload_0_16224;
  wire       [7:0]    _zz_dataOut_payload_0_16225;
  wire       [7:0]    _zz_dataOut_payload_128_48;
  wire                _zz_dataOut_payload_0_16226;
  wire       [7:0]    _zz_dataOut_payload_0_16227;
  wire       [7:0]    _zz_dataOut_payload_128_49;
  wire                _zz_dataOut_payload_0_16228;
  wire       [7:0]    _zz_dataOut_payload_0_16229;
  wire       [7:0]    _zz_dataOut_payload_128_50;
  wire                _zz_dataOut_payload_0_16230;
  wire       [7:0]    _zz_dataOut_payload_0_16231;
  wire       [7:0]    _zz_dataOut_payload_128_51;
  wire                _zz_dataOut_payload_0_16232;
  wire       [7:0]    _zz_dataOut_payload_0_16233;
  wire       [7:0]    _zz_dataOut_payload_128_52;
  wire                _zz_dataOut_payload_0_16234;
  wire       [7:0]    _zz_dataOut_payload_0_16235;
  wire       [7:0]    _zz_dataOut_payload_128_53;
  wire                _zz_dataOut_payload_0_16236;
  wire       [7:0]    _zz_dataOut_payload_0_16237;
  wire       [7:0]    _zz_dataOut_payload_128_54;
  wire                _zz_dataOut_payload_0_16238;
  wire       [7:0]    _zz_dataOut_payload_0_16239;
  wire       [7:0]    _zz_dataOut_payload_128_55;
  wire                _zz_dataOut_payload_0_16240;
  wire       [7:0]    _zz_dataOut_payload_0_16241;
  wire       [7:0]    _zz_dataOut_payload_128_56;
  wire                _zz_dataOut_payload_0_16242;
  wire       [7:0]    _zz_dataOut_payload_0_16243;
  wire       [7:0]    _zz_dataOut_payload_128_57;
  wire                _zz_dataOut_payload_0_16244;
  wire       [7:0]    _zz_dataOut_payload_0_16245;
  wire       [7:0]    _zz_dataOut_payload_128_58;
  wire                _zz_dataOut_payload_0_16246;
  wire       [7:0]    _zz_dataOut_payload_0_16247;
  wire       [7:0]    _zz_dataOut_payload_128_59;
  wire                _zz_dataOut_payload_0_16248;
  wire       [7:0]    _zz_dataOut_payload_0_16249;
  wire       [7:0]    _zz_dataOut_payload_128_60;
  wire                _zz_dataOut_payload_0_16250;
  wire       [7:0]    _zz_dataOut_payload_0_16251;
  wire       [7:0]    _zz_dataOut_payload_128_61;
  wire                _zz_dataOut_payload_0_16252;
  wire       [7:0]    _zz_dataOut_payload_0_16253;
  wire       [7:0]    _zz_dataOut_payload_128_62;
  wire                _zz_dataOut_payload_0_16254;
  wire       [7:0]    _zz_dataOut_payload_0_16255;
  wire       [7:0]    _zz_dataOut_payload_128_63;
  wire                _zz_dataOut_payload_0_16256;
  wire       [7:0]    _zz_dataOut_payload_0_16257;
  wire       [7:0]    _zz_dataOut_payload_128_64;
  wire                _zz_dataOut_payload_0_16258;
  wire       [7:0]    _zz_dataOut_payload_0_16259;
  wire       [7:0]    _zz_dataOut_payload_128_65;
  wire                _zz_dataOut_payload_0_16260;
  wire       [7:0]    _zz_dataOut_payload_0_16261;
  wire       [7:0]    _zz_dataOut_payload_128_66;
  wire                _zz_dataOut_payload_0_16262;
  wire       [7:0]    _zz_dataOut_payload_0_16263;
  wire       [7:0]    _zz_dataOut_payload_128_67;
  wire                _zz_dataOut_payload_0_16264;
  wire       [7:0]    _zz_dataOut_payload_0_16265;
  wire       [7:0]    _zz_dataOut_payload_128_68;
  wire                _zz_dataOut_payload_0_16266;
  wire       [7:0]    _zz_dataOut_payload_0_16267;
  wire       [7:0]    _zz_dataOut_payload_128_69;
  wire                _zz_dataOut_payload_0_16268;
  wire       [7:0]    _zz_dataOut_payload_0_16269;
  wire       [7:0]    _zz_dataOut_payload_128_70;
  wire                _zz_dataOut_payload_0_16270;
  wire       [7:0]    _zz_dataOut_payload_0_16271;
  wire       [7:0]    _zz_dataOut_payload_128_71;
  wire                _zz_dataOut_payload_0_16272;
  wire       [7:0]    _zz_dataOut_payload_0_16273;
  wire       [7:0]    _zz_dataOut_payload_128_72;
  wire                _zz_dataOut_payload_0_16274;
  wire       [7:0]    _zz_dataOut_payload_0_16275;
  wire       [7:0]    _zz_dataOut_payload_128_73;
  wire                _zz_dataOut_payload_0_16276;
  wire       [7:0]    _zz_dataOut_payload_0_16277;
  wire       [7:0]    _zz_dataOut_payload_128_74;
  wire                _zz_dataOut_payload_0_16278;
  wire       [7:0]    _zz_dataOut_payload_0_16279;
  wire       [7:0]    _zz_dataOut_payload_128_75;
  wire                _zz_dataOut_payload_0_16280;
  wire       [7:0]    _zz_dataOut_payload_0_16281;
  wire       [7:0]    _zz_dataOut_payload_128_76;
  wire                _zz_dataOut_payload_0_16282;
  wire       [7:0]    _zz_dataOut_payload_0_16283;
  wire       [7:0]    _zz_dataOut_payload_128_77;
  wire                _zz_dataOut_payload_0_16284;
  wire       [7:0]    _zz_dataOut_payload_0_16285;
  wire       [7:0]    _zz_dataOut_payload_128_78;
  wire                _zz_dataOut_payload_0_16286;
  wire       [7:0]    _zz_dataOut_payload_0_16287;
  wire       [7:0]    _zz_dataOut_payload_128_79;
  wire                _zz_dataOut_payload_0_16288;
  wire       [7:0]    _zz_dataOut_payload_0_16289;
  wire       [7:0]    _zz_dataOut_payload_128_80;
  wire                _zz_dataOut_payload_0_16290;
  wire       [7:0]    _zz_dataOut_payload_0_16291;
  wire       [7:0]    _zz_dataOut_payload_128_81;
  wire                _zz_dataOut_payload_0_16292;
  wire       [7:0]    _zz_dataOut_payload_0_16293;
  wire       [7:0]    _zz_dataOut_payload_128_82;
  wire                _zz_dataOut_payload_0_16294;
  wire       [7:0]    _zz_dataOut_payload_0_16295;
  wire       [7:0]    _zz_dataOut_payload_128_83;
  wire                _zz_dataOut_payload_0_16296;
  wire       [7:0]    _zz_dataOut_payload_0_16297;
  wire       [7:0]    _zz_dataOut_payload_128_84;
  wire                _zz_dataOut_payload_0_16298;
  wire       [7:0]    _zz_dataOut_payload_0_16299;
  wire       [7:0]    _zz_dataOut_payload_128_85;
  wire                _zz_dataOut_payload_0_16300;
  wire       [7:0]    _zz_dataOut_payload_0_16301;
  wire       [7:0]    _zz_dataOut_payload_128_86;
  wire                _zz_dataOut_payload_0_16302;
  wire       [7:0]    _zz_dataOut_payload_0_16303;
  wire       [7:0]    _zz_dataOut_payload_128_87;
  wire                _zz_dataOut_payload_0_16304;
  wire       [7:0]    _zz_dataOut_payload_0_16305;
  wire       [7:0]    _zz_dataOut_payload_128_88;
  wire                _zz_dataOut_payload_0_16306;
  wire       [7:0]    _zz_dataOut_payload_0_16307;
  wire       [7:0]    _zz_dataOut_payload_128_89;
  wire                _zz_dataOut_payload_0_16308;
  wire       [7:0]    _zz_dataOut_payload_0_16309;
  wire       [7:0]    _zz_dataOut_payload_128_90;
  wire                _zz_dataOut_payload_0_16310;
  wire       [7:0]    _zz_dataOut_payload_0_16311;
  wire       [7:0]    _zz_dataOut_payload_128_91;
  wire                _zz_dataOut_payload_0_16312;
  wire       [7:0]    _zz_dataOut_payload_0_16313;
  wire       [7:0]    _zz_dataOut_payload_128_92;
  wire                _zz_dataOut_payload_0_16314;
  wire       [7:0]    _zz_dataOut_payload_0_16315;
  wire       [7:0]    _zz_dataOut_payload_128_93;
  wire                _zz_dataOut_payload_0_16316;
  wire       [7:0]    _zz_dataOut_payload_0_16317;
  wire       [7:0]    _zz_dataOut_payload_128_94;
  wire                _zz_dataOut_payload_0_16318;
  wire       [7:0]    _zz_dataOut_payload_0_16319;
  wire       [7:0]    _zz_dataOut_payload_128_95;
  wire                _zz_dataOut_payload_0_16320;
  wire       [7:0]    _zz_dataOut_payload_0_16321;
  wire       [7:0]    _zz_dataOut_payload_128_96;
  wire                _zz_dataOut_payload_0_16322;
  wire       [7:0]    _zz_dataOut_payload_0_16323;
  wire       [7:0]    _zz_dataOut_payload_128_97;
  wire                _zz_dataOut_payload_0_16324;
  wire       [7:0]    _zz_dataOut_payload_0_16325;
  wire       [7:0]    _zz_dataOut_payload_128_98;
  wire                _zz_dataOut_payload_0_16326;
  wire       [7:0]    _zz_dataOut_payload_0_16327;
  wire       [7:0]    _zz_dataOut_payload_128_99;
  wire                _zz_dataOut_payload_0_16328;
  wire       [7:0]    _zz_dataOut_payload_0_16329;
  wire       [7:0]    _zz_dataOut_payload_128_100;
  wire                _zz_dataOut_payload_0_16330;
  wire       [7:0]    _zz_dataOut_payload_0_16331;
  wire       [7:0]    _zz_dataOut_payload_128_101;
  wire                _zz_dataOut_payload_0_16332;
  wire       [7:0]    _zz_dataOut_payload_0_16333;
  wire       [7:0]    _zz_dataOut_payload_128_102;
  wire                _zz_dataOut_payload_0_16334;
  wire       [7:0]    _zz_dataOut_payload_0_16335;
  wire       [7:0]    _zz_dataOut_payload_128_103;
  wire                _zz_dataOut_payload_0_16336;
  wire       [7:0]    _zz_dataOut_payload_0_16337;
  wire       [7:0]    _zz_dataOut_payload_128_104;
  wire                _zz_dataOut_payload_0_16338;
  wire       [7:0]    _zz_dataOut_payload_0_16339;
  wire       [7:0]    _zz_dataOut_payload_128_105;
  wire                _zz_dataOut_payload_0_16340;
  wire       [7:0]    _zz_dataOut_payload_0_16341;
  wire       [7:0]    _zz_dataOut_payload_128_106;
  wire                _zz_dataOut_payload_0_16342;
  wire       [7:0]    _zz_dataOut_payload_0_16343;
  wire       [7:0]    _zz_dataOut_payload_128_107;
  wire                _zz_dataOut_payload_0_16344;
  wire       [7:0]    _zz_dataOut_payload_0_16345;
  wire       [7:0]    _zz_dataOut_payload_128_108;
  wire                _zz_dataOut_payload_0_16346;
  wire       [7:0]    _zz_dataOut_payload_0_16347;
  wire       [7:0]    _zz_dataOut_payload_128_109;
  wire                _zz_dataOut_payload_0_16348;
  wire       [7:0]    _zz_dataOut_payload_0_16349;
  wire       [7:0]    _zz_dataOut_payload_128_110;
  wire                _zz_dataOut_payload_0_16350;
  wire       [7:0]    _zz_dataOut_payload_0_16351;
  wire       [7:0]    _zz_dataOut_payload_128_111;
  wire                _zz_dataOut_payload_0_16352;
  wire       [7:0]    _zz_dataOut_payload_0_16353;
  wire       [7:0]    _zz_dataOut_payload_128_112;
  wire                _zz_dataOut_payload_0_16354;
  wire       [7:0]    _zz_dataOut_payload_0_16355;
  wire       [7:0]    _zz_dataOut_payload_128_113;
  wire                _zz_dataOut_payload_0_16356;
  wire       [7:0]    _zz_dataOut_payload_0_16357;
  wire       [7:0]    _zz_dataOut_payload_128_114;
  wire                _zz_dataOut_payload_0_16358;
  wire       [7:0]    _zz_dataOut_payload_0_16359;
  wire       [7:0]    _zz_dataOut_payload_128_115;
  wire                _zz_dataOut_payload_0_16360;
  wire       [7:0]    _zz_dataOut_payload_0_16361;
  wire       [7:0]    _zz_dataOut_payload_128_116;
  wire                _zz_dataOut_payload_0_16362;
  wire       [7:0]    _zz_dataOut_payload_0_16363;
  wire       [7:0]    _zz_dataOut_payload_128_117;
  wire                _zz_dataOut_payload_0_16364;
  wire       [7:0]    _zz_dataOut_payload_0_16365;
  wire       [7:0]    _zz_dataOut_payload_128_118;
  wire                _zz_dataOut_payload_0_16366;
  wire       [7:0]    _zz_dataOut_payload_0_16367;
  wire       [7:0]    _zz_dataOut_payload_128_119;
  wire                _zz_dataOut_payload_0_16368;
  wire       [7:0]    _zz_dataOut_payload_0_16369;
  wire       [7:0]    _zz_dataOut_payload_128_120;
  wire                _zz_dataOut_payload_0_16370;
  wire       [7:0]    _zz_dataOut_payload_0_16371;
  wire       [7:0]    _zz_dataOut_payload_128_121;
  wire                _zz_dataOut_payload_0_16372;
  wire       [7:0]    _zz_dataOut_payload_0_16373;
  wire       [7:0]    _zz_dataOut_payload_128_122;
  wire                _zz_dataOut_payload_0_16374;
  wire       [7:0]    _zz_dataOut_payload_0_16375;
  wire       [7:0]    _zz_dataOut_payload_128_123;
  wire                _zz_dataOut_payload_0_16376;
  wire       [7:0]    _zz_dataOut_payload_0_16377;
  wire       [7:0]    _zz_dataOut_payload_128_124;
  wire                _zz_dataOut_payload_0_16378;
  wire       [7:0]    _zz_dataOut_payload_0_16379;
  wire       [7:0]    _zz_dataOut_payload_128_125;
  wire                _zz_dataOut_payload_0_16380;
  wire       [7:0]    _zz_dataOut_payload_0_16381;
  wire       [7:0]    _zz_dataOut_payload_128_126;
  wire                _zz_dataOut_payload_0_16382;
  wire       [7:0]    _zz_dataOut_payload_0_16383;
  wire       [7:0]    _zz_dataOut_payload_128_127;
  wire                _zz_dataOut_payload_0_16384;
  wire       [7:0]    _zz_dataOut_payload_0_16385;
  wire       [7:0]    _zz_dataOut_payload_64;
  wire                _zz_dataOut_payload_0_16386;
  wire       [7:0]    _zz_dataOut_payload_0_16387;
  wire       [7:0]    _zz_dataOut_payload_64_1;
  wire                _zz_dataOut_payload_0_16388;
  wire       [7:0]    _zz_dataOut_payload_0_16389;
  wire       [7:0]    _zz_dataOut_payload_64_2;
  wire                _zz_dataOut_payload_0_16390;
  wire       [7:0]    _zz_dataOut_payload_0_16391;
  wire       [7:0]    _zz_dataOut_payload_64_3;
  wire                _zz_dataOut_payload_0_16392;
  wire       [7:0]    _zz_dataOut_payload_0_16393;
  wire       [7:0]    _zz_dataOut_payload_64_4;
  wire                _zz_dataOut_payload_0_16394;
  wire       [7:0]    _zz_dataOut_payload_0_16395;
  wire       [7:0]    _zz_dataOut_payload_64_5;
  wire                _zz_dataOut_payload_0_16396;
  wire       [7:0]    _zz_dataOut_payload_0_16397;
  wire       [7:0]    _zz_dataOut_payload_64_6;
  wire                _zz_dataOut_payload_0_16398;
  wire       [7:0]    _zz_dataOut_payload_0_16399;
  wire       [7:0]    _zz_dataOut_payload_64_7;
  wire                _zz_dataOut_payload_0_16400;
  wire       [7:0]    _zz_dataOut_payload_0_16401;
  wire       [7:0]    _zz_dataOut_payload_64_8;
  wire                _zz_dataOut_payload_0_16402;
  wire       [7:0]    _zz_dataOut_payload_0_16403;
  wire       [7:0]    _zz_dataOut_payload_64_9;
  wire                _zz_dataOut_payload_0_16404;
  wire       [7:0]    _zz_dataOut_payload_0_16405;
  wire       [7:0]    _zz_dataOut_payload_64_10;
  wire                _zz_dataOut_payload_0_16406;
  wire       [7:0]    _zz_dataOut_payload_0_16407;
  wire       [7:0]    _zz_dataOut_payload_64_11;
  wire                _zz_dataOut_payload_0_16408;
  wire       [7:0]    _zz_dataOut_payload_0_16409;
  wire       [7:0]    _zz_dataOut_payload_64_12;
  wire                _zz_dataOut_payload_0_16410;
  wire       [7:0]    _zz_dataOut_payload_0_16411;
  wire       [7:0]    _zz_dataOut_payload_64_13;
  wire                _zz_dataOut_payload_0_16412;
  wire       [7:0]    _zz_dataOut_payload_0_16413;
  wire       [7:0]    _zz_dataOut_payload_64_14;
  wire                _zz_dataOut_payload_0_16414;
  wire       [7:0]    _zz_dataOut_payload_0_16415;
  wire       [7:0]    _zz_dataOut_payload_64_15;
  wire                _zz_dataOut_payload_0_16416;
  wire       [7:0]    _zz_dataOut_payload_0_16417;
  wire       [7:0]    _zz_dataOut_payload_64_16;
  wire                _zz_dataOut_payload_0_16418;
  wire       [7:0]    _zz_dataOut_payload_0_16419;
  wire       [7:0]    _zz_dataOut_payload_64_17;
  wire                _zz_dataOut_payload_0_16420;
  wire       [7:0]    _zz_dataOut_payload_0_16421;
  wire       [7:0]    _zz_dataOut_payload_64_18;
  wire                _zz_dataOut_payload_0_16422;
  wire       [7:0]    _zz_dataOut_payload_0_16423;
  wire       [7:0]    _zz_dataOut_payload_64_19;
  wire                _zz_dataOut_payload_0_16424;
  wire       [7:0]    _zz_dataOut_payload_0_16425;
  wire       [7:0]    _zz_dataOut_payload_64_20;
  wire                _zz_dataOut_payload_0_16426;
  wire       [7:0]    _zz_dataOut_payload_0_16427;
  wire       [7:0]    _zz_dataOut_payload_64_21;
  wire                _zz_dataOut_payload_0_16428;
  wire       [7:0]    _zz_dataOut_payload_0_16429;
  wire       [7:0]    _zz_dataOut_payload_64_22;
  wire                _zz_dataOut_payload_0_16430;
  wire       [7:0]    _zz_dataOut_payload_0_16431;
  wire       [7:0]    _zz_dataOut_payload_64_23;
  wire                _zz_dataOut_payload_0_16432;
  wire       [7:0]    _zz_dataOut_payload_0_16433;
  wire       [7:0]    _zz_dataOut_payload_64_24;
  wire                _zz_dataOut_payload_0_16434;
  wire       [7:0]    _zz_dataOut_payload_0_16435;
  wire       [7:0]    _zz_dataOut_payload_64_25;
  wire                _zz_dataOut_payload_0_16436;
  wire       [7:0]    _zz_dataOut_payload_0_16437;
  wire       [7:0]    _zz_dataOut_payload_64_26;
  wire                _zz_dataOut_payload_0_16438;
  wire       [7:0]    _zz_dataOut_payload_0_16439;
  wire       [7:0]    _zz_dataOut_payload_64_27;
  wire                _zz_dataOut_payload_0_16440;
  wire       [7:0]    _zz_dataOut_payload_0_16441;
  wire       [7:0]    _zz_dataOut_payload_64_28;
  wire                _zz_dataOut_payload_0_16442;
  wire       [7:0]    _zz_dataOut_payload_0_16443;
  wire       [7:0]    _zz_dataOut_payload_64_29;
  wire                _zz_dataOut_payload_0_16444;
  wire       [7:0]    _zz_dataOut_payload_0_16445;
  wire       [7:0]    _zz_dataOut_payload_64_30;
  wire                _zz_dataOut_payload_0_16446;
  wire       [7:0]    _zz_dataOut_payload_0_16447;
  wire       [7:0]    _zz_dataOut_payload_64_31;
  wire                _zz_dataOut_payload_0_16448;
  wire       [7:0]    _zz_dataOut_payload_0_16449;
  wire       [7:0]    _zz_dataOut_payload_64_32;
  wire                _zz_dataOut_payload_0_16450;
  wire       [7:0]    _zz_dataOut_payload_0_16451;
  wire       [7:0]    _zz_dataOut_payload_64_33;
  wire                _zz_dataOut_payload_0_16452;
  wire       [7:0]    _zz_dataOut_payload_0_16453;
  wire       [7:0]    _zz_dataOut_payload_64_34;
  wire                _zz_dataOut_payload_0_16454;
  wire       [7:0]    _zz_dataOut_payload_0_16455;
  wire       [7:0]    _zz_dataOut_payload_64_35;
  wire                _zz_dataOut_payload_0_16456;
  wire       [7:0]    _zz_dataOut_payload_0_16457;
  wire       [7:0]    _zz_dataOut_payload_64_36;
  wire                _zz_dataOut_payload_0_16458;
  wire       [7:0]    _zz_dataOut_payload_0_16459;
  wire       [7:0]    _zz_dataOut_payload_64_37;
  wire                _zz_dataOut_payload_0_16460;
  wire       [7:0]    _zz_dataOut_payload_0_16461;
  wire       [7:0]    _zz_dataOut_payload_64_38;
  wire                _zz_dataOut_payload_0_16462;
  wire       [7:0]    _zz_dataOut_payload_0_16463;
  wire       [7:0]    _zz_dataOut_payload_64_39;
  wire                _zz_dataOut_payload_0_16464;
  wire       [7:0]    _zz_dataOut_payload_0_16465;
  wire       [7:0]    _zz_dataOut_payload_64_40;
  wire                _zz_dataOut_payload_0_16466;
  wire       [7:0]    _zz_dataOut_payload_0_16467;
  wire       [7:0]    _zz_dataOut_payload_64_41;
  wire                _zz_dataOut_payload_0_16468;
  wire       [7:0]    _zz_dataOut_payload_0_16469;
  wire       [7:0]    _zz_dataOut_payload_64_42;
  wire                _zz_dataOut_payload_0_16470;
  wire       [7:0]    _zz_dataOut_payload_0_16471;
  wire       [7:0]    _zz_dataOut_payload_64_43;
  wire                _zz_dataOut_payload_0_16472;
  wire       [7:0]    _zz_dataOut_payload_0_16473;
  wire       [7:0]    _zz_dataOut_payload_64_44;
  wire                _zz_dataOut_payload_0_16474;
  wire       [7:0]    _zz_dataOut_payload_0_16475;
  wire       [7:0]    _zz_dataOut_payload_64_45;
  wire                _zz_dataOut_payload_0_16476;
  wire       [7:0]    _zz_dataOut_payload_0_16477;
  wire       [7:0]    _zz_dataOut_payload_64_46;
  wire                _zz_dataOut_payload_0_16478;
  wire       [7:0]    _zz_dataOut_payload_0_16479;
  wire       [7:0]    _zz_dataOut_payload_64_47;
  wire                _zz_dataOut_payload_0_16480;
  wire       [7:0]    _zz_dataOut_payload_0_16481;
  wire       [7:0]    _zz_dataOut_payload_64_48;
  wire                _zz_dataOut_payload_0_16482;
  wire       [7:0]    _zz_dataOut_payload_0_16483;
  wire       [7:0]    _zz_dataOut_payload_64_49;
  wire                _zz_dataOut_payload_0_16484;
  wire       [7:0]    _zz_dataOut_payload_0_16485;
  wire       [7:0]    _zz_dataOut_payload_64_50;
  wire                _zz_dataOut_payload_0_16486;
  wire       [7:0]    _zz_dataOut_payload_0_16487;
  wire       [7:0]    _zz_dataOut_payload_64_51;
  wire                _zz_dataOut_payload_0_16488;
  wire       [7:0]    _zz_dataOut_payload_0_16489;
  wire       [7:0]    _zz_dataOut_payload_64_52;
  wire                _zz_dataOut_payload_0_16490;
  wire       [7:0]    _zz_dataOut_payload_0_16491;
  wire       [7:0]    _zz_dataOut_payload_64_53;
  wire                _zz_dataOut_payload_0_16492;
  wire       [7:0]    _zz_dataOut_payload_0_16493;
  wire       [7:0]    _zz_dataOut_payload_64_54;
  wire                _zz_dataOut_payload_0_16494;
  wire       [7:0]    _zz_dataOut_payload_0_16495;
  wire       [7:0]    _zz_dataOut_payload_64_55;
  wire                _zz_dataOut_payload_0_16496;
  wire       [7:0]    _zz_dataOut_payload_0_16497;
  wire       [7:0]    _zz_dataOut_payload_64_56;
  wire                _zz_dataOut_payload_0_16498;
  wire       [7:0]    _zz_dataOut_payload_0_16499;
  wire       [7:0]    _zz_dataOut_payload_64_57;
  wire                _zz_dataOut_payload_0_16500;
  wire       [7:0]    _zz_dataOut_payload_0_16501;
  wire       [7:0]    _zz_dataOut_payload_64_58;
  wire                _zz_dataOut_payload_0_16502;
  wire       [7:0]    _zz_dataOut_payload_0_16503;
  wire       [7:0]    _zz_dataOut_payload_64_59;
  wire                _zz_dataOut_payload_0_16504;
  wire       [7:0]    _zz_dataOut_payload_0_16505;
  wire       [7:0]    _zz_dataOut_payload_64_60;
  wire                _zz_dataOut_payload_0_16506;
  wire       [7:0]    _zz_dataOut_payload_0_16507;
  wire       [7:0]    _zz_dataOut_payload_64_61;
  wire                _zz_dataOut_payload_0_16508;
  wire       [7:0]    _zz_dataOut_payload_0_16509;
  wire       [7:0]    _zz_dataOut_payload_64_62;
  wire                _zz_dataOut_payload_0_16510;
  wire       [7:0]    _zz_dataOut_payload_0_16511;
  wire       [7:0]    _zz_dataOut_payload_64_63;
  wire                _zz_dataOut_payload_0_16512;
  wire       [7:0]    _zz_dataOut_payload_0_16513;
  wire       [7:0]    _zz_dataOut_payload_32;
  wire                _zz_dataOut_payload_0_16514;
  wire       [7:0]    _zz_dataOut_payload_0_16515;
  wire       [7:0]    _zz_dataOut_payload_32_1;
  wire                _zz_dataOut_payload_0_16516;
  wire       [7:0]    _zz_dataOut_payload_0_16517;
  wire       [7:0]    _zz_dataOut_payload_32_2;
  wire                _zz_dataOut_payload_0_16518;
  wire       [7:0]    _zz_dataOut_payload_0_16519;
  wire       [7:0]    _zz_dataOut_payload_32_3;
  wire                _zz_dataOut_payload_0_16520;
  wire       [7:0]    _zz_dataOut_payload_0_16521;
  wire       [7:0]    _zz_dataOut_payload_32_4;
  wire                _zz_dataOut_payload_0_16522;
  wire       [7:0]    _zz_dataOut_payload_0_16523;
  wire       [7:0]    _zz_dataOut_payload_32_5;
  wire                _zz_dataOut_payload_0_16524;
  wire       [7:0]    _zz_dataOut_payload_0_16525;
  wire       [7:0]    _zz_dataOut_payload_32_6;
  wire                _zz_dataOut_payload_0_16526;
  wire       [7:0]    _zz_dataOut_payload_0_16527;
  wire       [7:0]    _zz_dataOut_payload_32_7;
  wire                _zz_dataOut_payload_0_16528;
  wire       [7:0]    _zz_dataOut_payload_0_16529;
  wire       [7:0]    _zz_dataOut_payload_32_8;
  wire                _zz_dataOut_payload_0_16530;
  wire       [7:0]    _zz_dataOut_payload_0_16531;
  wire       [7:0]    _zz_dataOut_payload_32_9;
  wire                _zz_dataOut_payload_0_16532;
  wire       [7:0]    _zz_dataOut_payload_0_16533;
  wire       [7:0]    _zz_dataOut_payload_32_10;
  wire                _zz_dataOut_payload_0_16534;
  wire       [7:0]    _zz_dataOut_payload_0_16535;
  wire       [7:0]    _zz_dataOut_payload_32_11;
  wire                _zz_dataOut_payload_0_16536;
  wire       [7:0]    _zz_dataOut_payload_0_16537;
  wire       [7:0]    _zz_dataOut_payload_32_12;
  wire                _zz_dataOut_payload_0_16538;
  wire       [7:0]    _zz_dataOut_payload_0_16539;
  wire       [7:0]    _zz_dataOut_payload_32_13;
  wire                _zz_dataOut_payload_0_16540;
  wire       [7:0]    _zz_dataOut_payload_0_16541;
  wire       [7:0]    _zz_dataOut_payload_32_14;
  wire                _zz_dataOut_payload_0_16542;
  wire       [7:0]    _zz_dataOut_payload_0_16543;
  wire       [7:0]    _zz_dataOut_payload_32_15;
  wire                _zz_dataOut_payload_0_16544;
  wire       [7:0]    _zz_dataOut_payload_0_16545;
  wire       [7:0]    _zz_dataOut_payload_32_16;
  wire                _zz_dataOut_payload_0_16546;
  wire       [7:0]    _zz_dataOut_payload_0_16547;
  wire       [7:0]    _zz_dataOut_payload_32_17;
  wire                _zz_dataOut_payload_0_16548;
  wire       [7:0]    _zz_dataOut_payload_0_16549;
  wire       [7:0]    _zz_dataOut_payload_32_18;
  wire                _zz_dataOut_payload_0_16550;
  wire       [7:0]    _zz_dataOut_payload_0_16551;
  wire       [7:0]    _zz_dataOut_payload_32_19;
  wire                _zz_dataOut_payload_0_16552;
  wire       [7:0]    _zz_dataOut_payload_0_16553;
  wire       [7:0]    _zz_dataOut_payload_32_20;
  wire                _zz_dataOut_payload_0_16554;
  wire       [7:0]    _zz_dataOut_payload_0_16555;
  wire       [7:0]    _zz_dataOut_payload_32_21;
  wire                _zz_dataOut_payload_0_16556;
  wire       [7:0]    _zz_dataOut_payload_0_16557;
  wire       [7:0]    _zz_dataOut_payload_32_22;
  wire                _zz_dataOut_payload_0_16558;
  wire       [7:0]    _zz_dataOut_payload_0_16559;
  wire       [7:0]    _zz_dataOut_payload_32_23;
  wire                _zz_dataOut_payload_0_16560;
  wire       [7:0]    _zz_dataOut_payload_0_16561;
  wire       [7:0]    _zz_dataOut_payload_32_24;
  wire                _zz_dataOut_payload_0_16562;
  wire       [7:0]    _zz_dataOut_payload_0_16563;
  wire       [7:0]    _zz_dataOut_payload_32_25;
  wire                _zz_dataOut_payload_0_16564;
  wire       [7:0]    _zz_dataOut_payload_0_16565;
  wire       [7:0]    _zz_dataOut_payload_32_26;
  wire                _zz_dataOut_payload_0_16566;
  wire       [7:0]    _zz_dataOut_payload_0_16567;
  wire       [7:0]    _zz_dataOut_payload_32_27;
  wire                _zz_dataOut_payload_0_16568;
  wire       [7:0]    _zz_dataOut_payload_0_16569;
  wire       [7:0]    _zz_dataOut_payload_32_28;
  wire                _zz_dataOut_payload_0_16570;
  wire       [7:0]    _zz_dataOut_payload_0_16571;
  wire       [7:0]    _zz_dataOut_payload_32_29;
  wire                _zz_dataOut_payload_0_16572;
  wire       [7:0]    _zz_dataOut_payload_0_16573;
  wire       [7:0]    _zz_dataOut_payload_32_30;
  wire                _zz_dataOut_payload_0_16574;
  wire       [7:0]    _zz_dataOut_payload_0_16575;
  wire       [7:0]    _zz_dataOut_payload_32_31;
  wire                _zz_dataOut_payload_0_16576;
  wire       [7:0]    _zz_dataOut_payload_0_16577;
  wire       [7:0]    _zz_dataOut_payload_16;
  wire                _zz_dataOut_payload_0_16578;
  wire       [7:0]    _zz_dataOut_payload_0_16579;
  wire       [7:0]    _zz_dataOut_payload_16_1;
  wire                _zz_dataOut_payload_0_16580;
  wire       [7:0]    _zz_dataOut_payload_0_16581;
  wire       [7:0]    _zz_dataOut_payload_16_2;
  wire                _zz_dataOut_payload_0_16582;
  wire       [7:0]    _zz_dataOut_payload_0_16583;
  wire       [7:0]    _zz_dataOut_payload_16_3;
  wire                _zz_dataOut_payload_0_16584;
  wire       [7:0]    _zz_dataOut_payload_0_16585;
  wire       [7:0]    _zz_dataOut_payload_16_4;
  wire                _zz_dataOut_payload_0_16586;
  wire       [7:0]    _zz_dataOut_payload_0_16587;
  wire       [7:0]    _zz_dataOut_payload_16_5;
  wire                _zz_dataOut_payload_0_16588;
  wire       [7:0]    _zz_dataOut_payload_0_16589;
  wire       [7:0]    _zz_dataOut_payload_16_6;
  wire                _zz_dataOut_payload_0_16590;
  wire       [7:0]    _zz_dataOut_payload_0_16591;
  wire       [7:0]    _zz_dataOut_payload_16_7;
  wire                _zz_dataOut_payload_0_16592;
  wire       [7:0]    _zz_dataOut_payload_0_16593;
  wire       [7:0]    _zz_dataOut_payload_16_8;
  wire                _zz_dataOut_payload_0_16594;
  wire       [7:0]    _zz_dataOut_payload_0_16595;
  wire       [7:0]    _zz_dataOut_payload_16_9;
  wire                _zz_dataOut_payload_0_16596;
  wire       [7:0]    _zz_dataOut_payload_0_16597;
  wire       [7:0]    _zz_dataOut_payload_16_10;
  wire                _zz_dataOut_payload_0_16598;
  wire       [7:0]    _zz_dataOut_payload_0_16599;
  wire       [7:0]    _zz_dataOut_payload_16_11;
  wire                _zz_dataOut_payload_0_16600;
  wire       [7:0]    _zz_dataOut_payload_0_16601;
  wire       [7:0]    _zz_dataOut_payload_16_12;
  wire                _zz_dataOut_payload_0_16602;
  wire       [7:0]    _zz_dataOut_payload_0_16603;
  wire       [7:0]    _zz_dataOut_payload_16_13;
  wire                _zz_dataOut_payload_0_16604;
  wire       [7:0]    _zz_dataOut_payload_0_16605;
  wire       [7:0]    _zz_dataOut_payload_16_14;
  wire                _zz_dataOut_payload_0_16606;
  wire       [7:0]    _zz_dataOut_payload_0_16607;
  wire       [7:0]    _zz_dataOut_payload_16_15;
  wire                _zz_dataOut_payload_0_16608;
  wire       [7:0]    _zz_dataOut_payload_0_16609;
  wire       [7:0]    _zz_dataOut_payload_8;
  wire                _zz_dataOut_payload_0_16610;
  wire       [7:0]    _zz_dataOut_payload_0_16611;
  wire       [7:0]    _zz_dataOut_payload_8_1;
  wire                _zz_dataOut_payload_0_16612;
  wire       [7:0]    _zz_dataOut_payload_0_16613;
  wire       [7:0]    _zz_dataOut_payload_8_2;
  wire                _zz_dataOut_payload_0_16614;
  wire       [7:0]    _zz_dataOut_payload_0_16615;
  wire       [7:0]    _zz_dataOut_payload_8_3;
  wire                _zz_dataOut_payload_0_16616;
  wire       [7:0]    _zz_dataOut_payload_0_16617;
  wire       [7:0]    _zz_dataOut_payload_8_4;
  wire                _zz_dataOut_payload_0_16618;
  wire       [7:0]    _zz_dataOut_payload_0_16619;
  wire       [7:0]    _zz_dataOut_payload_8_5;
  wire                _zz_dataOut_payload_0_16620;
  wire       [7:0]    _zz_dataOut_payload_0_16621;
  wire       [7:0]    _zz_dataOut_payload_8_6;
  wire                _zz_dataOut_payload_0_16622;
  wire       [7:0]    _zz_dataOut_payload_0_16623;
  wire       [7:0]    _zz_dataOut_payload_8_7;
  wire                _zz_dataOut_payload_0_16624;
  wire       [7:0]    _zz_dataOut_payload_0_16625;
  wire       [7:0]    _zz_dataOut_payload_4;
  wire                _zz_dataOut_payload_0_16626;
  wire       [7:0]    _zz_dataOut_payload_0_16627;
  wire       [7:0]    _zz_dataOut_payload_4_1;
  wire                _zz_dataOut_payload_0_16628;
  wire       [7:0]    _zz_dataOut_payload_0_16629;
  wire       [7:0]    _zz_dataOut_payload_4_2;
  wire                _zz_dataOut_payload_0_16630;
  wire       [7:0]    _zz_dataOut_payload_0_16631;
  wire       [7:0]    _zz_dataOut_payload_4_3;
  wire                _zz_dataOut_payload_0_16632;
  wire       [7:0]    _zz_dataOut_payload_0_16633;
  wire       [7:0]    _zz_dataOut_payload_2;
  wire                _zz_dataOut_payload_0_16634;
  wire       [7:0]    _zz_dataOut_payload_0_16635;
  wire       [7:0]    _zz_dataOut_payload_2_1;
  wire                _zz_dataOut_payload_0_16636;
  wire                _zz_dataOut_payload_2_2;
  reg        [7:0]    _zz_dataOut_payload_0_16637;
  reg        [7:0]    _zz_dataOut_payload_1;
  reg        [7:0]    _zz_dataOut_payload_2_3;
  reg        [7:0]    _zz_dataOut_payload_3;
  wire                _zz_dataOut_payload_4_4;
  wire       [7:0]    _zz_dataOut_payload_4_5;
  wire       [7:0]    _zz_dataOut_payload_6;
  wire                _zz_dataOut_payload_4_6;
  wire       [7:0]    _zz_dataOut_payload_4_7;
  wire       [7:0]    _zz_dataOut_payload_6_1;
  wire                _zz_dataOut_payload_4_8;
  wire                _zz_dataOut_payload_6_2;
  reg        [7:0]    _zz_dataOut_payload_4_9;
  reg        [7:0]    _zz_dataOut_payload_5;
  reg        [7:0]    _zz_dataOut_payload_6_3;
  reg        [7:0]    _zz_dataOut_payload_7;
  reg        [7:0]    _zz_dataOut_payload_0_16638;
  reg        [7:0]    _zz_dataOut_payload_1_1;
  reg        [7:0]    _zz_dataOut_payload_2_4;
  reg        [7:0]    _zz_dataOut_payload_3_1;
  reg        [7:0]    _zz_dataOut_payload_4_10;
  reg        [7:0]    _zz_dataOut_payload_5_1;
  reg        [7:0]    _zz_dataOut_payload_6_4;
  reg        [7:0]    _zz_dataOut_payload_7_1;
  wire                _zz_dataOut_payload_8_8;
  wire       [7:0]    _zz_dataOut_payload_8_9;
  wire       [7:0]    _zz_dataOut_payload_12;
  wire                _zz_dataOut_payload_8_10;
  wire       [7:0]    _zz_dataOut_payload_8_11;
  wire       [7:0]    _zz_dataOut_payload_12_1;
  wire                _zz_dataOut_payload_8_12;
  wire       [7:0]    _zz_dataOut_payload_8_13;
  wire       [7:0]    _zz_dataOut_payload_12_2;
  wire                _zz_dataOut_payload_8_14;
  wire       [7:0]    _zz_dataOut_payload_8_15;
  wire       [7:0]    _zz_dataOut_payload_12_3;
  wire                _zz_dataOut_payload_8_16;
  wire       [7:0]    _zz_dataOut_payload_8_17;
  wire       [7:0]    _zz_dataOut_payload_10;
  wire                _zz_dataOut_payload_8_18;
  wire       [7:0]    _zz_dataOut_payload_8_19;
  wire       [7:0]    _zz_dataOut_payload_10_1;
  wire                _zz_dataOut_payload_8_20;
  wire                _zz_dataOut_payload_10_2;
  reg        [7:0]    _zz_dataOut_payload_8_21;
  reg        [7:0]    _zz_dataOut_payload_9;
  reg        [7:0]    _zz_dataOut_payload_10_3;
  reg        [7:0]    _zz_dataOut_payload_11;
  wire                _zz_dataOut_payload_12_4;
  wire       [7:0]    _zz_dataOut_payload_12_5;
  wire       [7:0]    _zz_dataOut_payload_14;
  wire                _zz_dataOut_payload_12_6;
  wire       [7:0]    _zz_dataOut_payload_12_7;
  wire       [7:0]    _zz_dataOut_payload_14_1;
  wire                _zz_dataOut_payload_12_8;
  wire                _zz_dataOut_payload_14_2;
  reg        [7:0]    _zz_dataOut_payload_12_9;
  reg        [7:0]    _zz_dataOut_payload_13;
  reg        [7:0]    _zz_dataOut_payload_14_3;
  reg        [7:0]    _zz_dataOut_payload_15;
  reg        [7:0]    _zz_dataOut_payload_8_22;
  reg        [7:0]    _zz_dataOut_payload_9_1;
  reg        [7:0]    _zz_dataOut_payload_10_4;
  reg        [7:0]    _zz_dataOut_payload_11_1;
  reg        [7:0]    _zz_dataOut_payload_12_10;
  reg        [7:0]    _zz_dataOut_payload_13_1;
  reg        [7:0]    _zz_dataOut_payload_14_4;
  reg        [7:0]    _zz_dataOut_payload_15_1;
  reg        [7:0]    _zz_dataOut_payload_0_16639;
  reg        [7:0]    _zz_dataOut_payload_1_2;
  reg        [7:0]    _zz_dataOut_payload_2_5;
  reg        [7:0]    _zz_dataOut_payload_3_2;
  reg        [7:0]    _zz_dataOut_payload_4_11;
  reg        [7:0]    _zz_dataOut_payload_5_2;
  reg        [7:0]    _zz_dataOut_payload_6_5;
  reg        [7:0]    _zz_dataOut_payload_7_2;
  reg        [7:0]    _zz_dataOut_payload_8_23;
  reg        [7:0]    _zz_dataOut_payload_9_2;
  reg        [7:0]    _zz_dataOut_payload_10_5;
  reg        [7:0]    _zz_dataOut_payload_11_2;
  reg        [7:0]    _zz_dataOut_payload_12_11;
  reg        [7:0]    _zz_dataOut_payload_13_2;
  reg        [7:0]    _zz_dataOut_payload_14_5;
  reg        [7:0]    _zz_dataOut_payload_15_2;
  wire                _zz_dataOut_payload_16_16;
  wire       [7:0]    _zz_dataOut_payload_16_17;
  wire       [7:0]    _zz_dataOut_payload_24;
  wire                _zz_dataOut_payload_16_18;
  wire       [7:0]    _zz_dataOut_payload_16_19;
  wire       [7:0]    _zz_dataOut_payload_24_1;
  wire                _zz_dataOut_payload_16_20;
  wire       [7:0]    _zz_dataOut_payload_16_21;
  wire       [7:0]    _zz_dataOut_payload_24_2;
  wire                _zz_dataOut_payload_16_22;
  wire       [7:0]    _zz_dataOut_payload_16_23;
  wire       [7:0]    _zz_dataOut_payload_24_3;
  wire                _zz_dataOut_payload_16_24;
  wire       [7:0]    _zz_dataOut_payload_16_25;
  wire       [7:0]    _zz_dataOut_payload_24_4;
  wire                _zz_dataOut_payload_16_26;
  wire       [7:0]    _zz_dataOut_payload_16_27;
  wire       [7:0]    _zz_dataOut_payload_24_5;
  wire                _zz_dataOut_payload_16_28;
  wire       [7:0]    _zz_dataOut_payload_16_29;
  wire       [7:0]    _zz_dataOut_payload_24_6;
  wire                _zz_dataOut_payload_16_30;
  wire       [7:0]    _zz_dataOut_payload_16_31;
  wire       [7:0]    _zz_dataOut_payload_24_7;
  wire                _zz_dataOut_payload_16_32;
  wire       [7:0]    _zz_dataOut_payload_16_33;
  wire       [7:0]    _zz_dataOut_payload_20;
  wire                _zz_dataOut_payload_16_34;
  wire       [7:0]    _zz_dataOut_payload_16_35;
  wire       [7:0]    _zz_dataOut_payload_20_1;
  wire                _zz_dataOut_payload_16_36;
  wire       [7:0]    _zz_dataOut_payload_16_37;
  wire       [7:0]    _zz_dataOut_payload_20_2;
  wire                _zz_dataOut_payload_16_38;
  wire       [7:0]    _zz_dataOut_payload_16_39;
  wire       [7:0]    _zz_dataOut_payload_20_3;
  wire                _zz_dataOut_payload_16_40;
  wire       [7:0]    _zz_dataOut_payload_16_41;
  wire       [7:0]    _zz_dataOut_payload_18;
  wire                _zz_dataOut_payload_16_42;
  wire       [7:0]    _zz_dataOut_payload_16_43;
  wire       [7:0]    _zz_dataOut_payload_18_1;
  wire                _zz_dataOut_payload_16_44;
  wire                _zz_dataOut_payload_18_2;
  reg        [7:0]    _zz_dataOut_payload_16_45;
  reg        [7:0]    _zz_dataOut_payload_17;
  reg        [7:0]    _zz_dataOut_payload_18_3;
  reg        [7:0]    _zz_dataOut_payload_19;
  wire                _zz_dataOut_payload_20_4;
  wire       [7:0]    _zz_dataOut_payload_20_5;
  wire       [7:0]    _zz_dataOut_payload_22;
  wire                _zz_dataOut_payload_20_6;
  wire       [7:0]    _zz_dataOut_payload_20_7;
  wire       [7:0]    _zz_dataOut_payload_22_1;
  wire                _zz_dataOut_payload_20_8;
  wire                _zz_dataOut_payload_22_2;
  reg        [7:0]    _zz_dataOut_payload_20_9;
  reg        [7:0]    _zz_dataOut_payload_21;
  reg        [7:0]    _zz_dataOut_payload_22_3;
  reg        [7:0]    _zz_dataOut_payload_23;
  reg        [7:0]    _zz_dataOut_payload_16_46;
  reg        [7:0]    _zz_dataOut_payload_17_1;
  reg        [7:0]    _zz_dataOut_payload_18_4;
  reg        [7:0]    _zz_dataOut_payload_19_1;
  reg        [7:0]    _zz_dataOut_payload_20_10;
  reg        [7:0]    _zz_dataOut_payload_21_1;
  reg        [7:0]    _zz_dataOut_payload_22_4;
  reg        [7:0]    _zz_dataOut_payload_23_1;
  wire                _zz_dataOut_payload_24_8;
  wire       [7:0]    _zz_dataOut_payload_24_9;
  wire       [7:0]    _zz_dataOut_payload_28;
  wire                _zz_dataOut_payload_24_10;
  wire       [7:0]    _zz_dataOut_payload_24_11;
  wire       [7:0]    _zz_dataOut_payload_28_1;
  wire                _zz_dataOut_payload_24_12;
  wire       [7:0]    _zz_dataOut_payload_24_13;
  wire       [7:0]    _zz_dataOut_payload_28_2;
  wire                _zz_dataOut_payload_24_14;
  wire       [7:0]    _zz_dataOut_payload_24_15;
  wire       [7:0]    _zz_dataOut_payload_28_3;
  wire                _zz_dataOut_payload_24_16;
  wire       [7:0]    _zz_dataOut_payload_24_17;
  wire       [7:0]    _zz_dataOut_payload_26;
  wire                _zz_dataOut_payload_24_18;
  wire       [7:0]    _zz_dataOut_payload_24_19;
  wire       [7:0]    _zz_dataOut_payload_26_1;
  wire                _zz_dataOut_payload_24_20;
  wire                _zz_dataOut_payload_26_2;
  reg        [7:0]    _zz_dataOut_payload_24_21;
  reg        [7:0]    _zz_dataOut_payload_25;
  reg        [7:0]    _zz_dataOut_payload_26_3;
  reg        [7:0]    _zz_dataOut_payload_27;
  wire                _zz_dataOut_payload_28_4;
  wire       [7:0]    _zz_dataOut_payload_28_5;
  wire       [7:0]    _zz_dataOut_payload_30;
  wire                _zz_dataOut_payload_28_6;
  wire       [7:0]    _zz_dataOut_payload_28_7;
  wire       [7:0]    _zz_dataOut_payload_30_1;
  wire                _zz_dataOut_payload_28_8;
  wire                _zz_dataOut_payload_30_2;
  reg        [7:0]    _zz_dataOut_payload_28_9;
  reg        [7:0]    _zz_dataOut_payload_29;
  reg        [7:0]    _zz_dataOut_payload_30_3;
  reg        [7:0]    _zz_dataOut_payload_31;
  reg        [7:0]    _zz_dataOut_payload_24_22;
  reg        [7:0]    _zz_dataOut_payload_25_1;
  reg        [7:0]    _zz_dataOut_payload_26_4;
  reg        [7:0]    _zz_dataOut_payload_27_1;
  reg        [7:0]    _zz_dataOut_payload_28_10;
  reg        [7:0]    _zz_dataOut_payload_29_1;
  reg        [7:0]    _zz_dataOut_payload_30_4;
  reg        [7:0]    _zz_dataOut_payload_31_1;
  reg        [7:0]    _zz_dataOut_payload_16_47;
  reg        [7:0]    _zz_dataOut_payload_17_2;
  reg        [7:0]    _zz_dataOut_payload_18_5;
  reg        [7:0]    _zz_dataOut_payload_19_2;
  reg        [7:0]    _zz_dataOut_payload_20_11;
  reg        [7:0]    _zz_dataOut_payload_21_2;
  reg        [7:0]    _zz_dataOut_payload_22_5;
  reg        [7:0]    _zz_dataOut_payload_23_2;
  reg        [7:0]    _zz_dataOut_payload_24_23;
  reg        [7:0]    _zz_dataOut_payload_25_2;
  reg        [7:0]    _zz_dataOut_payload_26_5;
  reg        [7:0]    _zz_dataOut_payload_27_2;
  reg        [7:0]    _zz_dataOut_payload_28_11;
  reg        [7:0]    _zz_dataOut_payload_29_2;
  reg        [7:0]    _zz_dataOut_payload_30_5;
  reg        [7:0]    _zz_dataOut_payload_31_2;
  reg        [7:0]    _zz_dataOut_payload_0_16640;
  reg        [7:0]    _zz_dataOut_payload_1_3;
  reg        [7:0]    _zz_dataOut_payload_2_6;
  reg        [7:0]    _zz_dataOut_payload_3_3;
  reg        [7:0]    _zz_dataOut_payload_4_12;
  reg        [7:0]    _zz_dataOut_payload_5_3;
  reg        [7:0]    _zz_dataOut_payload_6_6;
  reg        [7:0]    _zz_dataOut_payload_7_3;
  reg        [7:0]    _zz_dataOut_payload_8_24;
  reg        [7:0]    _zz_dataOut_payload_9_3;
  reg        [7:0]    _zz_dataOut_payload_10_6;
  reg        [7:0]    _zz_dataOut_payload_11_3;
  reg        [7:0]    _zz_dataOut_payload_12_12;
  reg        [7:0]    _zz_dataOut_payload_13_3;
  reg        [7:0]    _zz_dataOut_payload_14_6;
  reg        [7:0]    _zz_dataOut_payload_15_3;
  reg        [7:0]    _zz_dataOut_payload_16_48;
  reg        [7:0]    _zz_dataOut_payload_17_3;
  reg        [7:0]    _zz_dataOut_payload_18_6;
  reg        [7:0]    _zz_dataOut_payload_19_3;
  reg        [7:0]    _zz_dataOut_payload_20_12;
  reg        [7:0]    _zz_dataOut_payload_21_3;
  reg        [7:0]    _zz_dataOut_payload_22_6;
  reg        [7:0]    _zz_dataOut_payload_23_3;
  reg        [7:0]    _zz_dataOut_payload_24_24;
  reg        [7:0]    _zz_dataOut_payload_25_3;
  reg        [7:0]    _zz_dataOut_payload_26_6;
  reg        [7:0]    _zz_dataOut_payload_27_3;
  reg        [7:0]    _zz_dataOut_payload_28_12;
  reg        [7:0]    _zz_dataOut_payload_29_3;
  reg        [7:0]    _zz_dataOut_payload_30_6;
  reg        [7:0]    _zz_dataOut_payload_31_3;
  wire                _zz_dataOut_payload_32_32;
  wire       [7:0]    _zz_dataOut_payload_32_33;
  wire       [7:0]    _zz_dataOut_payload_48;
  wire                _zz_dataOut_payload_32_34;
  wire       [7:0]    _zz_dataOut_payload_32_35;
  wire       [7:0]    _zz_dataOut_payload_48_1;
  wire                _zz_dataOut_payload_32_36;
  wire       [7:0]    _zz_dataOut_payload_32_37;
  wire       [7:0]    _zz_dataOut_payload_48_2;
  wire                _zz_dataOut_payload_32_38;
  wire       [7:0]    _zz_dataOut_payload_32_39;
  wire       [7:0]    _zz_dataOut_payload_48_3;
  wire                _zz_dataOut_payload_32_40;
  wire       [7:0]    _zz_dataOut_payload_32_41;
  wire       [7:0]    _zz_dataOut_payload_48_4;
  wire                _zz_dataOut_payload_32_42;
  wire       [7:0]    _zz_dataOut_payload_32_43;
  wire       [7:0]    _zz_dataOut_payload_48_5;
  wire                _zz_dataOut_payload_32_44;
  wire       [7:0]    _zz_dataOut_payload_32_45;
  wire       [7:0]    _zz_dataOut_payload_48_6;
  wire                _zz_dataOut_payload_32_46;
  wire       [7:0]    _zz_dataOut_payload_32_47;
  wire       [7:0]    _zz_dataOut_payload_48_7;
  wire                _zz_dataOut_payload_32_48;
  wire       [7:0]    _zz_dataOut_payload_32_49;
  wire       [7:0]    _zz_dataOut_payload_48_8;
  wire                _zz_dataOut_payload_32_50;
  wire       [7:0]    _zz_dataOut_payload_32_51;
  wire       [7:0]    _zz_dataOut_payload_48_9;
  wire                _zz_dataOut_payload_32_52;
  wire       [7:0]    _zz_dataOut_payload_32_53;
  wire       [7:0]    _zz_dataOut_payload_48_10;
  wire                _zz_dataOut_payload_32_54;
  wire       [7:0]    _zz_dataOut_payload_32_55;
  wire       [7:0]    _zz_dataOut_payload_48_11;
  wire                _zz_dataOut_payload_32_56;
  wire       [7:0]    _zz_dataOut_payload_32_57;
  wire       [7:0]    _zz_dataOut_payload_48_12;
  wire                _zz_dataOut_payload_32_58;
  wire       [7:0]    _zz_dataOut_payload_32_59;
  wire       [7:0]    _zz_dataOut_payload_48_13;
  wire                _zz_dataOut_payload_32_60;
  wire       [7:0]    _zz_dataOut_payload_32_61;
  wire       [7:0]    _zz_dataOut_payload_48_14;
  wire                _zz_dataOut_payload_32_62;
  wire       [7:0]    _zz_dataOut_payload_32_63;
  wire       [7:0]    _zz_dataOut_payload_48_15;
  wire                _zz_dataOut_payload_32_64;
  wire       [7:0]    _zz_dataOut_payload_32_65;
  wire       [7:0]    _zz_dataOut_payload_40;
  wire                _zz_dataOut_payload_32_66;
  wire       [7:0]    _zz_dataOut_payload_32_67;
  wire       [7:0]    _zz_dataOut_payload_40_1;
  wire                _zz_dataOut_payload_32_68;
  wire       [7:0]    _zz_dataOut_payload_32_69;
  wire       [7:0]    _zz_dataOut_payload_40_2;
  wire                _zz_dataOut_payload_32_70;
  wire       [7:0]    _zz_dataOut_payload_32_71;
  wire       [7:0]    _zz_dataOut_payload_40_3;
  wire                _zz_dataOut_payload_32_72;
  wire       [7:0]    _zz_dataOut_payload_32_73;
  wire       [7:0]    _zz_dataOut_payload_40_4;
  wire                _zz_dataOut_payload_32_74;
  wire       [7:0]    _zz_dataOut_payload_32_75;
  wire       [7:0]    _zz_dataOut_payload_40_5;
  wire                _zz_dataOut_payload_32_76;
  wire       [7:0]    _zz_dataOut_payload_32_77;
  wire       [7:0]    _zz_dataOut_payload_40_6;
  wire                _zz_dataOut_payload_32_78;
  wire       [7:0]    _zz_dataOut_payload_32_79;
  wire       [7:0]    _zz_dataOut_payload_40_7;
  wire                _zz_dataOut_payload_32_80;
  wire       [7:0]    _zz_dataOut_payload_32_81;
  wire       [7:0]    _zz_dataOut_payload_36;
  wire                _zz_dataOut_payload_32_82;
  wire       [7:0]    _zz_dataOut_payload_32_83;
  wire       [7:0]    _zz_dataOut_payload_36_1;
  wire                _zz_dataOut_payload_32_84;
  wire       [7:0]    _zz_dataOut_payload_32_85;
  wire       [7:0]    _zz_dataOut_payload_36_2;
  wire                _zz_dataOut_payload_32_86;
  wire       [7:0]    _zz_dataOut_payload_32_87;
  wire       [7:0]    _zz_dataOut_payload_36_3;
  wire                _zz_dataOut_payload_32_88;
  wire       [7:0]    _zz_dataOut_payload_32_89;
  wire       [7:0]    _zz_dataOut_payload_34;
  wire                _zz_dataOut_payload_32_90;
  wire       [7:0]    _zz_dataOut_payload_32_91;
  wire       [7:0]    _zz_dataOut_payload_34_1;
  wire                _zz_dataOut_payload_32_92;
  wire                _zz_dataOut_payload_34_2;
  reg        [7:0]    _zz_dataOut_payload_32_93;
  reg        [7:0]    _zz_dataOut_payload_33;
  reg        [7:0]    _zz_dataOut_payload_34_3;
  reg        [7:0]    _zz_dataOut_payload_35;
  wire                _zz_dataOut_payload_36_4;
  wire       [7:0]    _zz_dataOut_payload_36_5;
  wire       [7:0]    _zz_dataOut_payload_38;
  wire                _zz_dataOut_payload_36_6;
  wire       [7:0]    _zz_dataOut_payload_36_7;
  wire       [7:0]    _zz_dataOut_payload_38_1;
  wire                _zz_dataOut_payload_36_8;
  wire                _zz_dataOut_payload_38_2;
  reg        [7:0]    _zz_dataOut_payload_36_9;
  reg        [7:0]    _zz_dataOut_payload_37;
  reg        [7:0]    _zz_dataOut_payload_38_3;
  reg        [7:0]    _zz_dataOut_payload_39;
  reg        [7:0]    _zz_dataOut_payload_32_94;
  reg        [7:0]    _zz_dataOut_payload_33_1;
  reg        [7:0]    _zz_dataOut_payload_34_4;
  reg        [7:0]    _zz_dataOut_payload_35_1;
  reg        [7:0]    _zz_dataOut_payload_36_10;
  reg        [7:0]    _zz_dataOut_payload_37_1;
  reg        [7:0]    _zz_dataOut_payload_38_4;
  reg        [7:0]    _zz_dataOut_payload_39_1;
  wire                _zz_dataOut_payload_40_8;
  wire       [7:0]    _zz_dataOut_payload_40_9;
  wire       [7:0]    _zz_dataOut_payload_44;
  wire                _zz_dataOut_payload_40_10;
  wire       [7:0]    _zz_dataOut_payload_40_11;
  wire       [7:0]    _zz_dataOut_payload_44_1;
  wire                _zz_dataOut_payload_40_12;
  wire       [7:0]    _zz_dataOut_payload_40_13;
  wire       [7:0]    _zz_dataOut_payload_44_2;
  wire                _zz_dataOut_payload_40_14;
  wire       [7:0]    _zz_dataOut_payload_40_15;
  wire       [7:0]    _zz_dataOut_payload_44_3;
  wire                _zz_dataOut_payload_40_16;
  wire       [7:0]    _zz_dataOut_payload_40_17;
  wire       [7:0]    _zz_dataOut_payload_42;
  wire                _zz_dataOut_payload_40_18;
  wire       [7:0]    _zz_dataOut_payload_40_19;
  wire       [7:0]    _zz_dataOut_payload_42_1;
  wire                _zz_dataOut_payload_40_20;
  wire                _zz_dataOut_payload_42_2;
  reg        [7:0]    _zz_dataOut_payload_40_21;
  reg        [7:0]    _zz_dataOut_payload_41;
  reg        [7:0]    _zz_dataOut_payload_42_3;
  reg        [7:0]    _zz_dataOut_payload_43;
  wire                _zz_dataOut_payload_44_4;
  wire       [7:0]    _zz_dataOut_payload_44_5;
  wire       [7:0]    _zz_dataOut_payload_46;
  wire                _zz_dataOut_payload_44_6;
  wire       [7:0]    _zz_dataOut_payload_44_7;
  wire       [7:0]    _zz_dataOut_payload_46_1;
  wire                _zz_dataOut_payload_44_8;
  wire                _zz_dataOut_payload_46_2;
  reg        [7:0]    _zz_dataOut_payload_44_9;
  reg        [7:0]    _zz_dataOut_payload_45;
  reg        [7:0]    _zz_dataOut_payload_46_3;
  reg        [7:0]    _zz_dataOut_payload_47;
  reg        [7:0]    _zz_dataOut_payload_40_22;
  reg        [7:0]    _zz_dataOut_payload_41_1;
  reg        [7:0]    _zz_dataOut_payload_42_4;
  reg        [7:0]    _zz_dataOut_payload_43_1;
  reg        [7:0]    _zz_dataOut_payload_44_10;
  reg        [7:0]    _zz_dataOut_payload_45_1;
  reg        [7:0]    _zz_dataOut_payload_46_4;
  reg        [7:0]    _zz_dataOut_payload_47_1;
  reg        [7:0]    _zz_dataOut_payload_32_95;
  reg        [7:0]    _zz_dataOut_payload_33_2;
  reg        [7:0]    _zz_dataOut_payload_34_5;
  reg        [7:0]    _zz_dataOut_payload_35_2;
  reg        [7:0]    _zz_dataOut_payload_36_11;
  reg        [7:0]    _zz_dataOut_payload_37_2;
  reg        [7:0]    _zz_dataOut_payload_38_5;
  reg        [7:0]    _zz_dataOut_payload_39_2;
  reg        [7:0]    _zz_dataOut_payload_40_23;
  reg        [7:0]    _zz_dataOut_payload_41_2;
  reg        [7:0]    _zz_dataOut_payload_42_5;
  reg        [7:0]    _zz_dataOut_payload_43_2;
  reg        [7:0]    _zz_dataOut_payload_44_11;
  reg        [7:0]    _zz_dataOut_payload_45_2;
  reg        [7:0]    _zz_dataOut_payload_46_5;
  reg        [7:0]    _zz_dataOut_payload_47_2;
  wire                _zz_dataOut_payload_48_16;
  wire       [7:0]    _zz_dataOut_payload_48_17;
  wire       [7:0]    _zz_dataOut_payload_56;
  wire                _zz_dataOut_payload_48_18;
  wire       [7:0]    _zz_dataOut_payload_48_19;
  wire       [7:0]    _zz_dataOut_payload_56_1;
  wire                _zz_dataOut_payload_48_20;
  wire       [7:0]    _zz_dataOut_payload_48_21;
  wire       [7:0]    _zz_dataOut_payload_56_2;
  wire                _zz_dataOut_payload_48_22;
  wire       [7:0]    _zz_dataOut_payload_48_23;
  wire       [7:0]    _zz_dataOut_payload_56_3;
  wire                _zz_dataOut_payload_48_24;
  wire       [7:0]    _zz_dataOut_payload_48_25;
  wire       [7:0]    _zz_dataOut_payload_56_4;
  wire                _zz_dataOut_payload_48_26;
  wire       [7:0]    _zz_dataOut_payload_48_27;
  wire       [7:0]    _zz_dataOut_payload_56_5;
  wire                _zz_dataOut_payload_48_28;
  wire       [7:0]    _zz_dataOut_payload_48_29;
  wire       [7:0]    _zz_dataOut_payload_56_6;
  wire                _zz_dataOut_payload_48_30;
  wire       [7:0]    _zz_dataOut_payload_48_31;
  wire       [7:0]    _zz_dataOut_payload_56_7;
  wire                _zz_dataOut_payload_48_32;
  wire       [7:0]    _zz_dataOut_payload_48_33;
  wire       [7:0]    _zz_dataOut_payload_52;
  wire                _zz_dataOut_payload_48_34;
  wire       [7:0]    _zz_dataOut_payload_48_35;
  wire       [7:0]    _zz_dataOut_payload_52_1;
  wire                _zz_dataOut_payload_48_36;
  wire       [7:0]    _zz_dataOut_payload_48_37;
  wire       [7:0]    _zz_dataOut_payload_52_2;
  wire                _zz_dataOut_payload_48_38;
  wire       [7:0]    _zz_dataOut_payload_48_39;
  wire       [7:0]    _zz_dataOut_payload_52_3;
  wire                _zz_dataOut_payload_48_40;
  wire       [7:0]    _zz_dataOut_payload_48_41;
  wire       [7:0]    _zz_dataOut_payload_50;
  wire                _zz_dataOut_payload_48_42;
  wire       [7:0]    _zz_dataOut_payload_48_43;
  wire       [7:0]    _zz_dataOut_payload_50_1;
  wire                _zz_dataOut_payload_48_44;
  wire                _zz_dataOut_payload_50_2;
  reg        [7:0]    _zz_dataOut_payload_48_45;
  reg        [7:0]    _zz_dataOut_payload_49;
  reg        [7:0]    _zz_dataOut_payload_50_3;
  reg        [7:0]    _zz_dataOut_payload_51;
  wire                _zz_dataOut_payload_52_4;
  wire       [7:0]    _zz_dataOut_payload_52_5;
  wire       [7:0]    _zz_dataOut_payload_54;
  wire                _zz_dataOut_payload_52_6;
  wire       [7:0]    _zz_dataOut_payload_52_7;
  wire       [7:0]    _zz_dataOut_payload_54_1;
  wire                _zz_dataOut_payload_52_8;
  wire                _zz_dataOut_payload_54_2;
  reg        [7:0]    _zz_dataOut_payload_52_9;
  reg        [7:0]    _zz_dataOut_payload_53;
  reg        [7:0]    _zz_dataOut_payload_54_3;
  reg        [7:0]    _zz_dataOut_payload_55;
  reg        [7:0]    _zz_dataOut_payload_48_46;
  reg        [7:0]    _zz_dataOut_payload_49_1;
  reg        [7:0]    _zz_dataOut_payload_50_4;
  reg        [7:0]    _zz_dataOut_payload_51_1;
  reg        [7:0]    _zz_dataOut_payload_52_10;
  reg        [7:0]    _zz_dataOut_payload_53_1;
  reg        [7:0]    _zz_dataOut_payload_54_4;
  reg        [7:0]    _zz_dataOut_payload_55_1;
  wire                _zz_dataOut_payload_56_8;
  wire       [7:0]    _zz_dataOut_payload_56_9;
  wire       [7:0]    _zz_dataOut_payload_60;
  wire                _zz_dataOut_payload_56_10;
  wire       [7:0]    _zz_dataOut_payload_56_11;
  wire       [7:0]    _zz_dataOut_payload_60_1;
  wire                _zz_dataOut_payload_56_12;
  wire       [7:0]    _zz_dataOut_payload_56_13;
  wire       [7:0]    _zz_dataOut_payload_60_2;
  wire                _zz_dataOut_payload_56_14;
  wire       [7:0]    _zz_dataOut_payload_56_15;
  wire       [7:0]    _zz_dataOut_payload_60_3;
  wire                _zz_dataOut_payload_56_16;
  wire       [7:0]    _zz_dataOut_payload_56_17;
  wire       [7:0]    _zz_dataOut_payload_58;
  wire                _zz_dataOut_payload_56_18;
  wire       [7:0]    _zz_dataOut_payload_56_19;
  wire       [7:0]    _zz_dataOut_payload_58_1;
  wire                _zz_dataOut_payload_56_20;
  wire                _zz_dataOut_payload_58_2;
  reg        [7:0]    _zz_dataOut_payload_56_21;
  reg        [7:0]    _zz_dataOut_payload_57;
  reg        [7:0]    _zz_dataOut_payload_58_3;
  reg        [7:0]    _zz_dataOut_payload_59;
  wire                _zz_dataOut_payload_60_4;
  wire       [7:0]    _zz_dataOut_payload_60_5;
  wire       [7:0]    _zz_dataOut_payload_62;
  wire                _zz_dataOut_payload_60_6;
  wire       [7:0]    _zz_dataOut_payload_60_7;
  wire       [7:0]    _zz_dataOut_payload_62_1;
  wire                _zz_dataOut_payload_60_8;
  wire                _zz_dataOut_payload_62_2;
  reg        [7:0]    _zz_dataOut_payload_60_9;
  reg        [7:0]    _zz_dataOut_payload_61;
  reg        [7:0]    _zz_dataOut_payload_62_3;
  reg        [7:0]    _zz_dataOut_payload_63;
  reg        [7:0]    _zz_dataOut_payload_56_22;
  reg        [7:0]    _zz_dataOut_payload_57_1;
  reg        [7:0]    _zz_dataOut_payload_58_4;
  reg        [7:0]    _zz_dataOut_payload_59_1;
  reg        [7:0]    _zz_dataOut_payload_60_10;
  reg        [7:0]    _zz_dataOut_payload_61_1;
  reg        [7:0]    _zz_dataOut_payload_62_4;
  reg        [7:0]    _zz_dataOut_payload_63_1;
  reg        [7:0]    _zz_dataOut_payload_48_47;
  reg        [7:0]    _zz_dataOut_payload_49_2;
  reg        [7:0]    _zz_dataOut_payload_50_5;
  reg        [7:0]    _zz_dataOut_payload_51_2;
  reg        [7:0]    _zz_dataOut_payload_52_11;
  reg        [7:0]    _zz_dataOut_payload_53_2;
  reg        [7:0]    _zz_dataOut_payload_54_5;
  reg        [7:0]    _zz_dataOut_payload_55_2;
  reg        [7:0]    _zz_dataOut_payload_56_23;
  reg        [7:0]    _zz_dataOut_payload_57_2;
  reg        [7:0]    _zz_dataOut_payload_58_5;
  reg        [7:0]    _zz_dataOut_payload_59_2;
  reg        [7:0]    _zz_dataOut_payload_60_11;
  reg        [7:0]    _zz_dataOut_payload_61_2;
  reg        [7:0]    _zz_dataOut_payload_62_5;
  reg        [7:0]    _zz_dataOut_payload_63_2;
  reg        [7:0]    _zz_dataOut_payload_32_96;
  reg        [7:0]    _zz_dataOut_payload_33_3;
  reg        [7:0]    _zz_dataOut_payload_34_6;
  reg        [7:0]    _zz_dataOut_payload_35_3;
  reg        [7:0]    _zz_dataOut_payload_36_12;
  reg        [7:0]    _zz_dataOut_payload_37_3;
  reg        [7:0]    _zz_dataOut_payload_38_6;
  reg        [7:0]    _zz_dataOut_payload_39_3;
  reg        [7:0]    _zz_dataOut_payload_40_24;
  reg        [7:0]    _zz_dataOut_payload_41_3;
  reg        [7:0]    _zz_dataOut_payload_42_6;
  reg        [7:0]    _zz_dataOut_payload_43_3;
  reg        [7:0]    _zz_dataOut_payload_44_12;
  reg        [7:0]    _zz_dataOut_payload_45_3;
  reg        [7:0]    _zz_dataOut_payload_46_6;
  reg        [7:0]    _zz_dataOut_payload_47_3;
  reg        [7:0]    _zz_dataOut_payload_48_48;
  reg        [7:0]    _zz_dataOut_payload_49_3;
  reg        [7:0]    _zz_dataOut_payload_50_6;
  reg        [7:0]    _zz_dataOut_payload_51_3;
  reg        [7:0]    _zz_dataOut_payload_52_12;
  reg        [7:0]    _zz_dataOut_payload_53_3;
  reg        [7:0]    _zz_dataOut_payload_54_6;
  reg        [7:0]    _zz_dataOut_payload_55_3;
  reg        [7:0]    _zz_dataOut_payload_56_24;
  reg        [7:0]    _zz_dataOut_payload_57_3;
  reg        [7:0]    _zz_dataOut_payload_58_6;
  reg        [7:0]    _zz_dataOut_payload_59_3;
  reg        [7:0]    _zz_dataOut_payload_60_12;
  reg        [7:0]    _zz_dataOut_payload_61_3;
  reg        [7:0]    _zz_dataOut_payload_62_6;
  reg        [7:0]    _zz_dataOut_payload_63_3;
  reg        [7:0]    _zz_dataOut_payload_0_16641;
  reg        [7:0]    _zz_dataOut_payload_1_4;
  reg        [7:0]    _zz_dataOut_payload_2_7;
  reg        [7:0]    _zz_dataOut_payload_3_4;
  reg        [7:0]    _zz_dataOut_payload_4_13;
  reg        [7:0]    _zz_dataOut_payload_5_4;
  reg        [7:0]    _zz_dataOut_payload_6_7;
  reg        [7:0]    _zz_dataOut_payload_7_4;
  reg        [7:0]    _zz_dataOut_payload_8_25;
  reg        [7:0]    _zz_dataOut_payload_9_4;
  reg        [7:0]    _zz_dataOut_payload_10_7;
  reg        [7:0]    _zz_dataOut_payload_11_4;
  reg        [7:0]    _zz_dataOut_payload_12_13;
  reg        [7:0]    _zz_dataOut_payload_13_4;
  reg        [7:0]    _zz_dataOut_payload_14_7;
  reg        [7:0]    _zz_dataOut_payload_15_4;
  reg        [7:0]    _zz_dataOut_payload_16_49;
  reg        [7:0]    _zz_dataOut_payload_17_4;
  reg        [7:0]    _zz_dataOut_payload_18_7;
  reg        [7:0]    _zz_dataOut_payload_19_4;
  reg        [7:0]    _zz_dataOut_payload_20_13;
  reg        [7:0]    _zz_dataOut_payload_21_4;
  reg        [7:0]    _zz_dataOut_payload_22_7;
  reg        [7:0]    _zz_dataOut_payload_23_4;
  reg        [7:0]    _zz_dataOut_payload_24_25;
  reg        [7:0]    _zz_dataOut_payload_25_4;
  reg        [7:0]    _zz_dataOut_payload_26_7;
  reg        [7:0]    _zz_dataOut_payload_27_4;
  reg        [7:0]    _zz_dataOut_payload_28_13;
  reg        [7:0]    _zz_dataOut_payload_29_4;
  reg        [7:0]    _zz_dataOut_payload_30_7;
  reg        [7:0]    _zz_dataOut_payload_31_4;
  reg        [7:0]    _zz_dataOut_payload_32_97;
  reg        [7:0]    _zz_dataOut_payload_33_4;
  reg        [7:0]    _zz_dataOut_payload_34_7;
  reg        [7:0]    _zz_dataOut_payload_35_4;
  reg        [7:0]    _zz_dataOut_payload_36_13;
  reg        [7:0]    _zz_dataOut_payload_37_4;
  reg        [7:0]    _zz_dataOut_payload_38_7;
  reg        [7:0]    _zz_dataOut_payload_39_4;
  reg        [7:0]    _zz_dataOut_payload_40_25;
  reg        [7:0]    _zz_dataOut_payload_41_4;
  reg        [7:0]    _zz_dataOut_payload_42_7;
  reg        [7:0]    _zz_dataOut_payload_43_4;
  reg        [7:0]    _zz_dataOut_payload_44_13;
  reg        [7:0]    _zz_dataOut_payload_45_4;
  reg        [7:0]    _zz_dataOut_payload_46_7;
  reg        [7:0]    _zz_dataOut_payload_47_4;
  reg        [7:0]    _zz_dataOut_payload_48_49;
  reg        [7:0]    _zz_dataOut_payload_49_4;
  reg        [7:0]    _zz_dataOut_payload_50_7;
  reg        [7:0]    _zz_dataOut_payload_51_4;
  reg        [7:0]    _zz_dataOut_payload_52_13;
  reg        [7:0]    _zz_dataOut_payload_53_4;
  reg        [7:0]    _zz_dataOut_payload_54_7;
  reg        [7:0]    _zz_dataOut_payload_55_4;
  reg        [7:0]    _zz_dataOut_payload_56_25;
  reg        [7:0]    _zz_dataOut_payload_57_4;
  reg        [7:0]    _zz_dataOut_payload_58_7;
  reg        [7:0]    _zz_dataOut_payload_59_4;
  reg        [7:0]    _zz_dataOut_payload_60_13;
  reg        [7:0]    _zz_dataOut_payload_61_4;
  reg        [7:0]    _zz_dataOut_payload_62_7;
  reg        [7:0]    _zz_dataOut_payload_63_4;
  wire                _zz_dataOut_payload_64_64;
  wire       [7:0]    _zz_dataOut_payload_64_65;
  wire       [7:0]    _zz_dataOut_payload_96;
  wire                _zz_dataOut_payload_64_66;
  wire       [7:0]    _zz_dataOut_payload_64_67;
  wire       [7:0]    _zz_dataOut_payload_96_1;
  wire                _zz_dataOut_payload_64_68;
  wire       [7:0]    _zz_dataOut_payload_64_69;
  wire       [7:0]    _zz_dataOut_payload_96_2;
  wire                _zz_dataOut_payload_64_70;
  wire       [7:0]    _zz_dataOut_payload_64_71;
  wire       [7:0]    _zz_dataOut_payload_96_3;
  wire                _zz_dataOut_payload_64_72;
  wire       [7:0]    _zz_dataOut_payload_64_73;
  wire       [7:0]    _zz_dataOut_payload_96_4;
  wire                _zz_dataOut_payload_64_74;
  wire       [7:0]    _zz_dataOut_payload_64_75;
  wire       [7:0]    _zz_dataOut_payload_96_5;
  wire                _zz_dataOut_payload_64_76;
  wire       [7:0]    _zz_dataOut_payload_64_77;
  wire       [7:0]    _zz_dataOut_payload_96_6;
  wire                _zz_dataOut_payload_64_78;
  wire       [7:0]    _zz_dataOut_payload_64_79;
  wire       [7:0]    _zz_dataOut_payload_96_7;
  wire                _zz_dataOut_payload_64_80;
  wire       [7:0]    _zz_dataOut_payload_64_81;
  wire       [7:0]    _zz_dataOut_payload_96_8;
  wire                _zz_dataOut_payload_64_82;
  wire       [7:0]    _zz_dataOut_payload_64_83;
  wire       [7:0]    _zz_dataOut_payload_96_9;
  wire                _zz_dataOut_payload_64_84;
  wire       [7:0]    _zz_dataOut_payload_64_85;
  wire       [7:0]    _zz_dataOut_payload_96_10;
  wire                _zz_dataOut_payload_64_86;
  wire       [7:0]    _zz_dataOut_payload_64_87;
  wire       [7:0]    _zz_dataOut_payload_96_11;
  wire                _zz_dataOut_payload_64_88;
  wire       [7:0]    _zz_dataOut_payload_64_89;
  wire       [7:0]    _zz_dataOut_payload_96_12;
  wire                _zz_dataOut_payload_64_90;
  wire       [7:0]    _zz_dataOut_payload_64_91;
  wire       [7:0]    _zz_dataOut_payload_96_13;
  wire                _zz_dataOut_payload_64_92;
  wire       [7:0]    _zz_dataOut_payload_64_93;
  wire       [7:0]    _zz_dataOut_payload_96_14;
  wire                _zz_dataOut_payload_64_94;
  wire       [7:0]    _zz_dataOut_payload_64_95;
  wire       [7:0]    _zz_dataOut_payload_96_15;
  wire                _zz_dataOut_payload_64_96;
  wire       [7:0]    _zz_dataOut_payload_64_97;
  wire       [7:0]    _zz_dataOut_payload_96_16;
  wire                _zz_dataOut_payload_64_98;
  wire       [7:0]    _zz_dataOut_payload_64_99;
  wire       [7:0]    _zz_dataOut_payload_96_17;
  wire                _zz_dataOut_payload_64_100;
  wire       [7:0]    _zz_dataOut_payload_64_101;
  wire       [7:0]    _zz_dataOut_payload_96_18;
  wire                _zz_dataOut_payload_64_102;
  wire       [7:0]    _zz_dataOut_payload_64_103;
  wire       [7:0]    _zz_dataOut_payload_96_19;
  wire                _zz_dataOut_payload_64_104;
  wire       [7:0]    _zz_dataOut_payload_64_105;
  wire       [7:0]    _zz_dataOut_payload_96_20;
  wire                _zz_dataOut_payload_64_106;
  wire       [7:0]    _zz_dataOut_payload_64_107;
  wire       [7:0]    _zz_dataOut_payload_96_21;
  wire                _zz_dataOut_payload_64_108;
  wire       [7:0]    _zz_dataOut_payload_64_109;
  wire       [7:0]    _zz_dataOut_payload_96_22;
  wire                _zz_dataOut_payload_64_110;
  wire       [7:0]    _zz_dataOut_payload_64_111;
  wire       [7:0]    _zz_dataOut_payload_96_23;
  wire                _zz_dataOut_payload_64_112;
  wire       [7:0]    _zz_dataOut_payload_64_113;
  wire       [7:0]    _zz_dataOut_payload_96_24;
  wire                _zz_dataOut_payload_64_114;
  wire       [7:0]    _zz_dataOut_payload_64_115;
  wire       [7:0]    _zz_dataOut_payload_96_25;
  wire                _zz_dataOut_payload_64_116;
  wire       [7:0]    _zz_dataOut_payload_64_117;
  wire       [7:0]    _zz_dataOut_payload_96_26;
  wire                _zz_dataOut_payload_64_118;
  wire       [7:0]    _zz_dataOut_payload_64_119;
  wire       [7:0]    _zz_dataOut_payload_96_27;
  wire                _zz_dataOut_payload_64_120;
  wire       [7:0]    _zz_dataOut_payload_64_121;
  wire       [7:0]    _zz_dataOut_payload_96_28;
  wire                _zz_dataOut_payload_64_122;
  wire       [7:0]    _zz_dataOut_payload_64_123;
  wire       [7:0]    _zz_dataOut_payload_96_29;
  wire                _zz_dataOut_payload_64_124;
  wire       [7:0]    _zz_dataOut_payload_64_125;
  wire       [7:0]    _zz_dataOut_payload_96_30;
  wire                _zz_dataOut_payload_64_126;
  wire       [7:0]    _zz_dataOut_payload_64_127;
  wire       [7:0]    _zz_dataOut_payload_96_31;
  wire                _zz_dataOut_payload_64_128;
  wire       [7:0]    _zz_dataOut_payload_64_129;
  wire       [7:0]    _zz_dataOut_payload_80;
  wire                _zz_dataOut_payload_64_130;
  wire       [7:0]    _zz_dataOut_payload_64_131;
  wire       [7:0]    _zz_dataOut_payload_80_1;
  wire                _zz_dataOut_payload_64_132;
  wire       [7:0]    _zz_dataOut_payload_64_133;
  wire       [7:0]    _zz_dataOut_payload_80_2;
  wire                _zz_dataOut_payload_64_134;
  wire       [7:0]    _zz_dataOut_payload_64_135;
  wire       [7:0]    _zz_dataOut_payload_80_3;
  wire                _zz_dataOut_payload_64_136;
  wire       [7:0]    _zz_dataOut_payload_64_137;
  wire       [7:0]    _zz_dataOut_payload_80_4;
  wire                _zz_dataOut_payload_64_138;
  wire       [7:0]    _zz_dataOut_payload_64_139;
  wire       [7:0]    _zz_dataOut_payload_80_5;
  wire                _zz_dataOut_payload_64_140;
  wire       [7:0]    _zz_dataOut_payload_64_141;
  wire       [7:0]    _zz_dataOut_payload_80_6;
  wire                _zz_dataOut_payload_64_142;
  wire       [7:0]    _zz_dataOut_payload_64_143;
  wire       [7:0]    _zz_dataOut_payload_80_7;
  wire                _zz_dataOut_payload_64_144;
  wire       [7:0]    _zz_dataOut_payload_64_145;
  wire       [7:0]    _zz_dataOut_payload_80_8;
  wire                _zz_dataOut_payload_64_146;
  wire       [7:0]    _zz_dataOut_payload_64_147;
  wire       [7:0]    _zz_dataOut_payload_80_9;
  wire                _zz_dataOut_payload_64_148;
  wire       [7:0]    _zz_dataOut_payload_64_149;
  wire       [7:0]    _zz_dataOut_payload_80_10;
  wire                _zz_dataOut_payload_64_150;
  wire       [7:0]    _zz_dataOut_payload_64_151;
  wire       [7:0]    _zz_dataOut_payload_80_11;
  wire                _zz_dataOut_payload_64_152;
  wire       [7:0]    _zz_dataOut_payload_64_153;
  wire       [7:0]    _zz_dataOut_payload_80_12;
  wire                _zz_dataOut_payload_64_154;
  wire       [7:0]    _zz_dataOut_payload_64_155;
  wire       [7:0]    _zz_dataOut_payload_80_13;
  wire                _zz_dataOut_payload_64_156;
  wire       [7:0]    _zz_dataOut_payload_64_157;
  wire       [7:0]    _zz_dataOut_payload_80_14;
  wire                _zz_dataOut_payload_64_158;
  wire       [7:0]    _zz_dataOut_payload_64_159;
  wire       [7:0]    _zz_dataOut_payload_80_15;
  wire                _zz_dataOut_payload_64_160;
  wire       [7:0]    _zz_dataOut_payload_64_161;
  wire       [7:0]    _zz_dataOut_payload_72;
  wire                _zz_dataOut_payload_64_162;
  wire       [7:0]    _zz_dataOut_payload_64_163;
  wire       [7:0]    _zz_dataOut_payload_72_1;
  wire                _zz_dataOut_payload_64_164;
  wire       [7:0]    _zz_dataOut_payload_64_165;
  wire       [7:0]    _zz_dataOut_payload_72_2;
  wire                _zz_dataOut_payload_64_166;
  wire       [7:0]    _zz_dataOut_payload_64_167;
  wire       [7:0]    _zz_dataOut_payload_72_3;
  wire                _zz_dataOut_payload_64_168;
  wire       [7:0]    _zz_dataOut_payload_64_169;
  wire       [7:0]    _zz_dataOut_payload_72_4;
  wire                _zz_dataOut_payload_64_170;
  wire       [7:0]    _zz_dataOut_payload_64_171;
  wire       [7:0]    _zz_dataOut_payload_72_5;
  wire                _zz_dataOut_payload_64_172;
  wire       [7:0]    _zz_dataOut_payload_64_173;
  wire       [7:0]    _zz_dataOut_payload_72_6;
  wire                _zz_dataOut_payload_64_174;
  wire       [7:0]    _zz_dataOut_payload_64_175;
  wire       [7:0]    _zz_dataOut_payload_72_7;
  wire                _zz_dataOut_payload_64_176;
  wire       [7:0]    _zz_dataOut_payload_64_177;
  wire       [7:0]    _zz_dataOut_payload_68;
  wire                _zz_dataOut_payload_64_178;
  wire       [7:0]    _zz_dataOut_payload_64_179;
  wire       [7:0]    _zz_dataOut_payload_68_1;
  wire                _zz_dataOut_payload_64_180;
  wire       [7:0]    _zz_dataOut_payload_64_181;
  wire       [7:0]    _zz_dataOut_payload_68_2;
  wire                _zz_dataOut_payload_64_182;
  wire       [7:0]    _zz_dataOut_payload_64_183;
  wire       [7:0]    _zz_dataOut_payload_68_3;
  wire                _zz_dataOut_payload_64_184;
  wire       [7:0]    _zz_dataOut_payload_64_185;
  wire       [7:0]    _zz_dataOut_payload_66;
  wire                _zz_dataOut_payload_64_186;
  wire       [7:0]    _zz_dataOut_payload_64_187;
  wire       [7:0]    _zz_dataOut_payload_66_1;
  wire                _zz_dataOut_payload_64_188;
  wire                _zz_dataOut_payload_66_2;
  reg        [7:0]    _zz_dataOut_payload_64_189;
  reg        [7:0]    _zz_dataOut_payload_65;
  reg        [7:0]    _zz_dataOut_payload_66_3;
  reg        [7:0]    _zz_dataOut_payload_67;
  wire                _zz_dataOut_payload_68_4;
  wire       [7:0]    _zz_dataOut_payload_68_5;
  wire       [7:0]    _zz_dataOut_payload_70;
  wire                _zz_dataOut_payload_68_6;
  wire       [7:0]    _zz_dataOut_payload_68_7;
  wire       [7:0]    _zz_dataOut_payload_70_1;
  wire                _zz_dataOut_payload_68_8;
  wire                _zz_dataOut_payload_70_2;
  reg        [7:0]    _zz_dataOut_payload_68_9;
  reg        [7:0]    _zz_dataOut_payload_69;
  reg        [7:0]    _zz_dataOut_payload_70_3;
  reg        [7:0]    _zz_dataOut_payload_71;
  reg        [7:0]    _zz_dataOut_payload_64_190;
  reg        [7:0]    _zz_dataOut_payload_65_1;
  reg        [7:0]    _zz_dataOut_payload_66_4;
  reg        [7:0]    _zz_dataOut_payload_67_1;
  reg        [7:0]    _zz_dataOut_payload_68_10;
  reg        [7:0]    _zz_dataOut_payload_69_1;
  reg        [7:0]    _zz_dataOut_payload_70_4;
  reg        [7:0]    _zz_dataOut_payload_71_1;
  wire                _zz_dataOut_payload_72_8;
  wire       [7:0]    _zz_dataOut_payload_72_9;
  wire       [7:0]    _zz_dataOut_payload_76;
  wire                _zz_dataOut_payload_72_10;
  wire       [7:0]    _zz_dataOut_payload_72_11;
  wire       [7:0]    _zz_dataOut_payload_76_1;
  wire                _zz_dataOut_payload_72_12;
  wire       [7:0]    _zz_dataOut_payload_72_13;
  wire       [7:0]    _zz_dataOut_payload_76_2;
  wire                _zz_dataOut_payload_72_14;
  wire       [7:0]    _zz_dataOut_payload_72_15;
  wire       [7:0]    _zz_dataOut_payload_76_3;
  wire                _zz_dataOut_payload_72_16;
  wire       [7:0]    _zz_dataOut_payload_72_17;
  wire       [7:0]    _zz_dataOut_payload_74;
  wire                _zz_dataOut_payload_72_18;
  wire       [7:0]    _zz_dataOut_payload_72_19;
  wire       [7:0]    _zz_dataOut_payload_74_1;
  wire                _zz_dataOut_payload_72_20;
  wire                _zz_dataOut_payload_74_2;
  reg        [7:0]    _zz_dataOut_payload_72_21;
  reg        [7:0]    _zz_dataOut_payload_73;
  reg        [7:0]    _zz_dataOut_payload_74_3;
  reg        [7:0]    _zz_dataOut_payload_75;
  wire                _zz_dataOut_payload_76_4;
  wire       [7:0]    _zz_dataOut_payload_76_5;
  wire       [7:0]    _zz_dataOut_payload_78;
  wire                _zz_dataOut_payload_76_6;
  wire       [7:0]    _zz_dataOut_payload_76_7;
  wire       [7:0]    _zz_dataOut_payload_78_1;
  wire                _zz_dataOut_payload_76_8;
  wire                _zz_dataOut_payload_78_2;
  reg        [7:0]    _zz_dataOut_payload_76_9;
  reg        [7:0]    _zz_dataOut_payload_77;
  reg        [7:0]    _zz_dataOut_payload_78_3;
  reg        [7:0]    _zz_dataOut_payload_79;
  reg        [7:0]    _zz_dataOut_payload_72_22;
  reg        [7:0]    _zz_dataOut_payload_73_1;
  reg        [7:0]    _zz_dataOut_payload_74_4;
  reg        [7:0]    _zz_dataOut_payload_75_1;
  reg        [7:0]    _zz_dataOut_payload_76_10;
  reg        [7:0]    _zz_dataOut_payload_77_1;
  reg        [7:0]    _zz_dataOut_payload_78_4;
  reg        [7:0]    _zz_dataOut_payload_79_1;
  reg        [7:0]    _zz_dataOut_payload_64_191;
  reg        [7:0]    _zz_dataOut_payload_65_2;
  reg        [7:0]    _zz_dataOut_payload_66_5;
  reg        [7:0]    _zz_dataOut_payload_67_2;
  reg        [7:0]    _zz_dataOut_payload_68_11;
  reg        [7:0]    _zz_dataOut_payload_69_2;
  reg        [7:0]    _zz_dataOut_payload_70_5;
  reg        [7:0]    _zz_dataOut_payload_71_2;
  reg        [7:0]    _zz_dataOut_payload_72_23;
  reg        [7:0]    _zz_dataOut_payload_73_2;
  reg        [7:0]    _zz_dataOut_payload_74_5;
  reg        [7:0]    _zz_dataOut_payload_75_2;
  reg        [7:0]    _zz_dataOut_payload_76_11;
  reg        [7:0]    _zz_dataOut_payload_77_2;
  reg        [7:0]    _zz_dataOut_payload_78_5;
  reg        [7:0]    _zz_dataOut_payload_79_2;
  wire                _zz_dataOut_payload_80_16;
  wire       [7:0]    _zz_dataOut_payload_80_17;
  wire       [7:0]    _zz_dataOut_payload_88;
  wire                _zz_dataOut_payload_80_18;
  wire       [7:0]    _zz_dataOut_payload_80_19;
  wire       [7:0]    _zz_dataOut_payload_88_1;
  wire                _zz_dataOut_payload_80_20;
  wire       [7:0]    _zz_dataOut_payload_80_21;
  wire       [7:0]    _zz_dataOut_payload_88_2;
  wire                _zz_dataOut_payload_80_22;
  wire       [7:0]    _zz_dataOut_payload_80_23;
  wire       [7:0]    _zz_dataOut_payload_88_3;
  wire                _zz_dataOut_payload_80_24;
  wire       [7:0]    _zz_dataOut_payload_80_25;
  wire       [7:0]    _zz_dataOut_payload_88_4;
  wire                _zz_dataOut_payload_80_26;
  wire       [7:0]    _zz_dataOut_payload_80_27;
  wire       [7:0]    _zz_dataOut_payload_88_5;
  wire                _zz_dataOut_payload_80_28;
  wire       [7:0]    _zz_dataOut_payload_80_29;
  wire       [7:0]    _zz_dataOut_payload_88_6;
  wire                _zz_dataOut_payload_80_30;
  wire       [7:0]    _zz_dataOut_payload_80_31;
  wire       [7:0]    _zz_dataOut_payload_88_7;
  wire                _zz_dataOut_payload_80_32;
  wire       [7:0]    _zz_dataOut_payload_80_33;
  wire       [7:0]    _zz_dataOut_payload_84;
  wire                _zz_dataOut_payload_80_34;
  wire       [7:0]    _zz_dataOut_payload_80_35;
  wire       [7:0]    _zz_dataOut_payload_84_1;
  wire                _zz_dataOut_payload_80_36;
  wire       [7:0]    _zz_dataOut_payload_80_37;
  wire       [7:0]    _zz_dataOut_payload_84_2;
  wire                _zz_dataOut_payload_80_38;
  wire       [7:0]    _zz_dataOut_payload_80_39;
  wire       [7:0]    _zz_dataOut_payload_84_3;
  wire                _zz_dataOut_payload_80_40;
  wire       [7:0]    _zz_dataOut_payload_80_41;
  wire       [7:0]    _zz_dataOut_payload_82;
  wire                _zz_dataOut_payload_80_42;
  wire       [7:0]    _zz_dataOut_payload_80_43;
  wire       [7:0]    _zz_dataOut_payload_82_1;
  wire                _zz_dataOut_payload_80_44;
  wire                _zz_dataOut_payload_82_2;
  reg        [7:0]    _zz_dataOut_payload_80_45;
  reg        [7:0]    _zz_dataOut_payload_81;
  reg        [7:0]    _zz_dataOut_payload_82_3;
  reg        [7:0]    _zz_dataOut_payload_83;
  wire                _zz_dataOut_payload_84_4;
  wire       [7:0]    _zz_dataOut_payload_84_5;
  wire       [7:0]    _zz_dataOut_payload_86;
  wire                _zz_dataOut_payload_84_6;
  wire       [7:0]    _zz_dataOut_payload_84_7;
  wire       [7:0]    _zz_dataOut_payload_86_1;
  wire                _zz_dataOut_payload_84_8;
  wire                _zz_dataOut_payload_86_2;
  reg        [7:0]    _zz_dataOut_payload_84_9;
  reg        [7:0]    _zz_dataOut_payload_85;
  reg        [7:0]    _zz_dataOut_payload_86_3;
  reg        [7:0]    _zz_dataOut_payload_87;
  reg        [7:0]    _zz_dataOut_payload_80_46;
  reg        [7:0]    _zz_dataOut_payload_81_1;
  reg        [7:0]    _zz_dataOut_payload_82_4;
  reg        [7:0]    _zz_dataOut_payload_83_1;
  reg        [7:0]    _zz_dataOut_payload_84_10;
  reg        [7:0]    _zz_dataOut_payload_85_1;
  reg        [7:0]    _zz_dataOut_payload_86_4;
  reg        [7:0]    _zz_dataOut_payload_87_1;
  wire                _zz_dataOut_payload_88_8;
  wire       [7:0]    _zz_dataOut_payload_88_9;
  wire       [7:0]    _zz_dataOut_payload_92;
  wire                _zz_dataOut_payload_88_10;
  wire       [7:0]    _zz_dataOut_payload_88_11;
  wire       [7:0]    _zz_dataOut_payload_92_1;
  wire                _zz_dataOut_payload_88_12;
  wire       [7:0]    _zz_dataOut_payload_88_13;
  wire       [7:0]    _zz_dataOut_payload_92_2;
  wire                _zz_dataOut_payload_88_14;
  wire       [7:0]    _zz_dataOut_payload_88_15;
  wire       [7:0]    _zz_dataOut_payload_92_3;
  wire                _zz_dataOut_payload_88_16;
  wire       [7:0]    _zz_dataOut_payload_88_17;
  wire       [7:0]    _zz_dataOut_payload_90;
  wire                _zz_dataOut_payload_88_18;
  wire       [7:0]    _zz_dataOut_payload_88_19;
  wire       [7:0]    _zz_dataOut_payload_90_1;
  wire                _zz_dataOut_payload_88_20;
  wire                _zz_dataOut_payload_90_2;
  reg        [7:0]    _zz_dataOut_payload_88_21;
  reg        [7:0]    _zz_dataOut_payload_89;
  reg        [7:0]    _zz_dataOut_payload_90_3;
  reg        [7:0]    _zz_dataOut_payload_91;
  wire                _zz_dataOut_payload_92_4;
  wire       [7:0]    _zz_dataOut_payload_92_5;
  wire       [7:0]    _zz_dataOut_payload_94;
  wire                _zz_dataOut_payload_92_6;
  wire       [7:0]    _zz_dataOut_payload_92_7;
  wire       [7:0]    _zz_dataOut_payload_94_1;
  wire                _zz_dataOut_payload_92_8;
  wire                _zz_dataOut_payload_94_2;
  reg        [7:0]    _zz_dataOut_payload_92_9;
  reg        [7:0]    _zz_dataOut_payload_93;
  reg        [7:0]    _zz_dataOut_payload_94_3;
  reg        [7:0]    _zz_dataOut_payload_95;
  reg        [7:0]    _zz_dataOut_payload_88_22;
  reg        [7:0]    _zz_dataOut_payload_89_1;
  reg        [7:0]    _zz_dataOut_payload_90_4;
  reg        [7:0]    _zz_dataOut_payload_91_1;
  reg        [7:0]    _zz_dataOut_payload_92_10;
  reg        [7:0]    _zz_dataOut_payload_93_1;
  reg        [7:0]    _zz_dataOut_payload_94_4;
  reg        [7:0]    _zz_dataOut_payload_95_1;
  reg        [7:0]    _zz_dataOut_payload_80_47;
  reg        [7:0]    _zz_dataOut_payload_81_2;
  reg        [7:0]    _zz_dataOut_payload_82_5;
  reg        [7:0]    _zz_dataOut_payload_83_2;
  reg        [7:0]    _zz_dataOut_payload_84_11;
  reg        [7:0]    _zz_dataOut_payload_85_2;
  reg        [7:0]    _zz_dataOut_payload_86_5;
  reg        [7:0]    _zz_dataOut_payload_87_2;
  reg        [7:0]    _zz_dataOut_payload_88_23;
  reg        [7:0]    _zz_dataOut_payload_89_2;
  reg        [7:0]    _zz_dataOut_payload_90_5;
  reg        [7:0]    _zz_dataOut_payload_91_2;
  reg        [7:0]    _zz_dataOut_payload_92_11;
  reg        [7:0]    _zz_dataOut_payload_93_2;
  reg        [7:0]    _zz_dataOut_payload_94_5;
  reg        [7:0]    _zz_dataOut_payload_95_2;
  reg        [7:0]    _zz_dataOut_payload_64_192;
  reg        [7:0]    _zz_dataOut_payload_65_3;
  reg        [7:0]    _zz_dataOut_payload_66_6;
  reg        [7:0]    _zz_dataOut_payload_67_3;
  reg        [7:0]    _zz_dataOut_payload_68_12;
  reg        [7:0]    _zz_dataOut_payload_69_3;
  reg        [7:0]    _zz_dataOut_payload_70_6;
  reg        [7:0]    _zz_dataOut_payload_71_3;
  reg        [7:0]    _zz_dataOut_payload_72_24;
  reg        [7:0]    _zz_dataOut_payload_73_3;
  reg        [7:0]    _zz_dataOut_payload_74_6;
  reg        [7:0]    _zz_dataOut_payload_75_3;
  reg        [7:0]    _zz_dataOut_payload_76_12;
  reg        [7:0]    _zz_dataOut_payload_77_3;
  reg        [7:0]    _zz_dataOut_payload_78_6;
  reg        [7:0]    _zz_dataOut_payload_79_3;
  reg        [7:0]    _zz_dataOut_payload_80_48;
  reg        [7:0]    _zz_dataOut_payload_81_3;
  reg        [7:0]    _zz_dataOut_payload_82_6;
  reg        [7:0]    _zz_dataOut_payload_83_3;
  reg        [7:0]    _zz_dataOut_payload_84_12;
  reg        [7:0]    _zz_dataOut_payload_85_3;
  reg        [7:0]    _zz_dataOut_payload_86_6;
  reg        [7:0]    _zz_dataOut_payload_87_3;
  reg        [7:0]    _zz_dataOut_payload_88_24;
  reg        [7:0]    _zz_dataOut_payload_89_3;
  reg        [7:0]    _zz_dataOut_payload_90_6;
  reg        [7:0]    _zz_dataOut_payload_91_3;
  reg        [7:0]    _zz_dataOut_payload_92_12;
  reg        [7:0]    _zz_dataOut_payload_93_3;
  reg        [7:0]    _zz_dataOut_payload_94_6;
  reg        [7:0]    _zz_dataOut_payload_95_3;
  wire                _zz_dataOut_payload_96_32;
  wire       [7:0]    _zz_dataOut_payload_96_33;
  wire       [7:0]    _zz_dataOut_payload_112;
  wire                _zz_dataOut_payload_96_34;
  wire       [7:0]    _zz_dataOut_payload_96_35;
  wire       [7:0]    _zz_dataOut_payload_112_1;
  wire                _zz_dataOut_payload_96_36;
  wire       [7:0]    _zz_dataOut_payload_96_37;
  wire       [7:0]    _zz_dataOut_payload_112_2;
  wire                _zz_dataOut_payload_96_38;
  wire       [7:0]    _zz_dataOut_payload_96_39;
  wire       [7:0]    _zz_dataOut_payload_112_3;
  wire                _zz_dataOut_payload_96_40;
  wire       [7:0]    _zz_dataOut_payload_96_41;
  wire       [7:0]    _zz_dataOut_payload_112_4;
  wire                _zz_dataOut_payload_96_42;
  wire       [7:0]    _zz_dataOut_payload_96_43;
  wire       [7:0]    _zz_dataOut_payload_112_5;
  wire                _zz_dataOut_payload_96_44;
  wire       [7:0]    _zz_dataOut_payload_96_45;
  wire       [7:0]    _zz_dataOut_payload_112_6;
  wire                _zz_dataOut_payload_96_46;
  wire       [7:0]    _zz_dataOut_payload_96_47;
  wire       [7:0]    _zz_dataOut_payload_112_7;
  wire                _zz_dataOut_payload_96_48;
  wire       [7:0]    _zz_dataOut_payload_96_49;
  wire       [7:0]    _zz_dataOut_payload_112_8;
  wire                _zz_dataOut_payload_96_50;
  wire       [7:0]    _zz_dataOut_payload_96_51;
  wire       [7:0]    _zz_dataOut_payload_112_9;
  wire                _zz_dataOut_payload_96_52;
  wire       [7:0]    _zz_dataOut_payload_96_53;
  wire       [7:0]    _zz_dataOut_payload_112_10;
  wire                _zz_dataOut_payload_96_54;
  wire       [7:0]    _zz_dataOut_payload_96_55;
  wire       [7:0]    _zz_dataOut_payload_112_11;
  wire                _zz_dataOut_payload_96_56;
  wire       [7:0]    _zz_dataOut_payload_96_57;
  wire       [7:0]    _zz_dataOut_payload_112_12;
  wire                _zz_dataOut_payload_96_58;
  wire       [7:0]    _zz_dataOut_payload_96_59;
  wire       [7:0]    _zz_dataOut_payload_112_13;
  wire                _zz_dataOut_payload_96_60;
  wire       [7:0]    _zz_dataOut_payload_96_61;
  wire       [7:0]    _zz_dataOut_payload_112_14;
  wire                _zz_dataOut_payload_96_62;
  wire       [7:0]    _zz_dataOut_payload_96_63;
  wire       [7:0]    _zz_dataOut_payload_112_15;
  wire                _zz_dataOut_payload_96_64;
  wire       [7:0]    _zz_dataOut_payload_96_65;
  wire       [7:0]    _zz_dataOut_payload_104;
  wire                _zz_dataOut_payload_96_66;
  wire       [7:0]    _zz_dataOut_payload_96_67;
  wire       [7:0]    _zz_dataOut_payload_104_1;
  wire                _zz_dataOut_payload_96_68;
  wire       [7:0]    _zz_dataOut_payload_96_69;
  wire       [7:0]    _zz_dataOut_payload_104_2;
  wire                _zz_dataOut_payload_96_70;
  wire       [7:0]    _zz_dataOut_payload_96_71;
  wire       [7:0]    _zz_dataOut_payload_104_3;
  wire                _zz_dataOut_payload_96_72;
  wire       [7:0]    _zz_dataOut_payload_96_73;
  wire       [7:0]    _zz_dataOut_payload_104_4;
  wire                _zz_dataOut_payload_96_74;
  wire       [7:0]    _zz_dataOut_payload_96_75;
  wire       [7:0]    _zz_dataOut_payload_104_5;
  wire                _zz_dataOut_payload_96_76;
  wire       [7:0]    _zz_dataOut_payload_96_77;
  wire       [7:0]    _zz_dataOut_payload_104_6;
  wire                _zz_dataOut_payload_96_78;
  wire       [7:0]    _zz_dataOut_payload_96_79;
  wire       [7:0]    _zz_dataOut_payload_104_7;
  wire                _zz_dataOut_payload_96_80;
  wire       [7:0]    _zz_dataOut_payload_96_81;
  wire       [7:0]    _zz_dataOut_payload_100;
  wire                _zz_dataOut_payload_96_82;
  wire       [7:0]    _zz_dataOut_payload_96_83;
  wire       [7:0]    _zz_dataOut_payload_100_1;
  wire                _zz_dataOut_payload_96_84;
  wire       [7:0]    _zz_dataOut_payload_96_85;
  wire       [7:0]    _zz_dataOut_payload_100_2;
  wire                _zz_dataOut_payload_96_86;
  wire       [7:0]    _zz_dataOut_payload_96_87;
  wire       [7:0]    _zz_dataOut_payload_100_3;
  wire                _zz_dataOut_payload_96_88;
  wire       [7:0]    _zz_dataOut_payload_96_89;
  wire       [7:0]    _zz_dataOut_payload_98;
  wire                _zz_dataOut_payload_96_90;
  wire       [7:0]    _zz_dataOut_payload_96_91;
  wire       [7:0]    _zz_dataOut_payload_98_1;
  wire                _zz_dataOut_payload_96_92;
  wire                _zz_dataOut_payload_98_2;
  reg        [7:0]    _zz_dataOut_payload_96_93;
  reg        [7:0]    _zz_dataOut_payload_97;
  reg        [7:0]    _zz_dataOut_payload_98_3;
  reg        [7:0]    _zz_dataOut_payload_99;
  wire                _zz_dataOut_payload_100_4;
  wire       [7:0]    _zz_dataOut_payload_100_5;
  wire       [7:0]    _zz_dataOut_payload_102;
  wire                _zz_dataOut_payload_100_6;
  wire       [7:0]    _zz_dataOut_payload_100_7;
  wire       [7:0]    _zz_dataOut_payload_102_1;
  wire                _zz_dataOut_payload_100_8;
  wire                _zz_dataOut_payload_102_2;
  reg        [7:0]    _zz_dataOut_payload_100_9;
  reg        [7:0]    _zz_dataOut_payload_101;
  reg        [7:0]    _zz_dataOut_payload_102_3;
  reg        [7:0]    _zz_dataOut_payload_103;
  reg        [7:0]    _zz_dataOut_payload_96_94;
  reg        [7:0]    _zz_dataOut_payload_97_1;
  reg        [7:0]    _zz_dataOut_payload_98_4;
  reg        [7:0]    _zz_dataOut_payload_99_1;
  reg        [7:0]    _zz_dataOut_payload_100_10;
  reg        [7:0]    _zz_dataOut_payload_101_1;
  reg        [7:0]    _zz_dataOut_payload_102_4;
  reg        [7:0]    _zz_dataOut_payload_103_1;
  wire                _zz_dataOut_payload_104_8;
  wire       [7:0]    _zz_dataOut_payload_104_9;
  wire       [7:0]    _zz_dataOut_payload_108;
  wire                _zz_dataOut_payload_104_10;
  wire       [7:0]    _zz_dataOut_payload_104_11;
  wire       [7:0]    _zz_dataOut_payload_108_1;
  wire                _zz_dataOut_payload_104_12;
  wire       [7:0]    _zz_dataOut_payload_104_13;
  wire       [7:0]    _zz_dataOut_payload_108_2;
  wire                _zz_dataOut_payload_104_14;
  wire       [7:0]    _zz_dataOut_payload_104_15;
  wire       [7:0]    _zz_dataOut_payload_108_3;
  wire                _zz_dataOut_payload_104_16;
  wire       [7:0]    _zz_dataOut_payload_104_17;
  wire       [7:0]    _zz_dataOut_payload_106;
  wire                _zz_dataOut_payload_104_18;
  wire       [7:0]    _zz_dataOut_payload_104_19;
  wire       [7:0]    _zz_dataOut_payload_106_1;
  wire                _zz_dataOut_payload_104_20;
  wire                _zz_dataOut_payload_106_2;
  reg        [7:0]    _zz_dataOut_payload_104_21;
  reg        [7:0]    _zz_dataOut_payload_105;
  reg        [7:0]    _zz_dataOut_payload_106_3;
  reg        [7:0]    _zz_dataOut_payload_107;
  wire                _zz_dataOut_payload_108_4;
  wire       [7:0]    _zz_dataOut_payload_108_5;
  wire       [7:0]    _zz_dataOut_payload_110;
  wire                _zz_dataOut_payload_108_6;
  wire       [7:0]    _zz_dataOut_payload_108_7;
  wire       [7:0]    _zz_dataOut_payload_110_1;
  wire                _zz_dataOut_payload_108_8;
  wire                _zz_dataOut_payload_110_2;
  reg        [7:0]    _zz_dataOut_payload_108_9;
  reg        [7:0]    _zz_dataOut_payload_109;
  reg        [7:0]    _zz_dataOut_payload_110_3;
  reg        [7:0]    _zz_dataOut_payload_111;
  reg        [7:0]    _zz_dataOut_payload_104_22;
  reg        [7:0]    _zz_dataOut_payload_105_1;
  reg        [7:0]    _zz_dataOut_payload_106_4;
  reg        [7:0]    _zz_dataOut_payload_107_1;
  reg        [7:0]    _zz_dataOut_payload_108_10;
  reg        [7:0]    _zz_dataOut_payload_109_1;
  reg        [7:0]    _zz_dataOut_payload_110_4;
  reg        [7:0]    _zz_dataOut_payload_111_1;
  reg        [7:0]    _zz_dataOut_payload_96_95;
  reg        [7:0]    _zz_dataOut_payload_97_2;
  reg        [7:0]    _zz_dataOut_payload_98_5;
  reg        [7:0]    _zz_dataOut_payload_99_2;
  reg        [7:0]    _zz_dataOut_payload_100_11;
  reg        [7:0]    _zz_dataOut_payload_101_2;
  reg        [7:0]    _zz_dataOut_payload_102_5;
  reg        [7:0]    _zz_dataOut_payload_103_2;
  reg        [7:0]    _zz_dataOut_payload_104_23;
  reg        [7:0]    _zz_dataOut_payload_105_2;
  reg        [7:0]    _zz_dataOut_payload_106_5;
  reg        [7:0]    _zz_dataOut_payload_107_2;
  reg        [7:0]    _zz_dataOut_payload_108_11;
  reg        [7:0]    _zz_dataOut_payload_109_2;
  reg        [7:0]    _zz_dataOut_payload_110_5;
  reg        [7:0]    _zz_dataOut_payload_111_2;
  wire                _zz_dataOut_payload_112_16;
  wire       [7:0]    _zz_dataOut_payload_112_17;
  wire       [7:0]    _zz_dataOut_payload_120;
  wire                _zz_dataOut_payload_112_18;
  wire       [7:0]    _zz_dataOut_payload_112_19;
  wire       [7:0]    _zz_dataOut_payload_120_1;
  wire                _zz_dataOut_payload_112_20;
  wire       [7:0]    _zz_dataOut_payload_112_21;
  wire       [7:0]    _zz_dataOut_payload_120_2;
  wire                _zz_dataOut_payload_112_22;
  wire       [7:0]    _zz_dataOut_payload_112_23;
  wire       [7:0]    _zz_dataOut_payload_120_3;
  wire                _zz_dataOut_payload_112_24;
  wire       [7:0]    _zz_dataOut_payload_112_25;
  wire       [7:0]    _zz_dataOut_payload_120_4;
  wire                _zz_dataOut_payload_112_26;
  wire       [7:0]    _zz_dataOut_payload_112_27;
  wire       [7:0]    _zz_dataOut_payload_120_5;
  wire                _zz_dataOut_payload_112_28;
  wire       [7:0]    _zz_dataOut_payload_112_29;
  wire       [7:0]    _zz_dataOut_payload_120_6;
  wire                _zz_dataOut_payload_112_30;
  wire       [7:0]    _zz_dataOut_payload_112_31;
  wire       [7:0]    _zz_dataOut_payload_120_7;
  wire                _zz_dataOut_payload_112_32;
  wire       [7:0]    _zz_dataOut_payload_112_33;
  wire       [7:0]    _zz_dataOut_payload_116;
  wire                _zz_dataOut_payload_112_34;
  wire       [7:0]    _zz_dataOut_payload_112_35;
  wire       [7:0]    _zz_dataOut_payload_116_1;
  wire                _zz_dataOut_payload_112_36;
  wire       [7:0]    _zz_dataOut_payload_112_37;
  wire       [7:0]    _zz_dataOut_payload_116_2;
  wire                _zz_dataOut_payload_112_38;
  wire       [7:0]    _zz_dataOut_payload_112_39;
  wire       [7:0]    _zz_dataOut_payload_116_3;
  wire                _zz_dataOut_payload_112_40;
  wire       [7:0]    _zz_dataOut_payload_112_41;
  wire       [7:0]    _zz_dataOut_payload_114;
  wire                _zz_dataOut_payload_112_42;
  wire       [7:0]    _zz_dataOut_payload_112_43;
  wire       [7:0]    _zz_dataOut_payload_114_1;
  wire                _zz_dataOut_payload_112_44;
  wire                _zz_dataOut_payload_114_2;
  reg        [7:0]    _zz_dataOut_payload_112_45;
  reg        [7:0]    _zz_dataOut_payload_113;
  reg        [7:0]    _zz_dataOut_payload_114_3;
  reg        [7:0]    _zz_dataOut_payload_115;
  wire                _zz_dataOut_payload_116_4;
  wire       [7:0]    _zz_dataOut_payload_116_5;
  wire       [7:0]    _zz_dataOut_payload_118;
  wire                _zz_dataOut_payload_116_6;
  wire       [7:0]    _zz_dataOut_payload_116_7;
  wire       [7:0]    _zz_dataOut_payload_118_1;
  wire                _zz_dataOut_payload_116_8;
  wire                _zz_dataOut_payload_118_2;
  reg        [7:0]    _zz_dataOut_payload_116_9;
  reg        [7:0]    _zz_dataOut_payload_117;
  reg        [7:0]    _zz_dataOut_payload_118_3;
  reg        [7:0]    _zz_dataOut_payload_119;
  reg        [7:0]    _zz_dataOut_payload_112_46;
  reg        [7:0]    _zz_dataOut_payload_113_1;
  reg        [7:0]    _zz_dataOut_payload_114_4;
  reg        [7:0]    _zz_dataOut_payload_115_1;
  reg        [7:0]    _zz_dataOut_payload_116_10;
  reg        [7:0]    _zz_dataOut_payload_117_1;
  reg        [7:0]    _zz_dataOut_payload_118_4;
  reg        [7:0]    _zz_dataOut_payload_119_1;
  wire                _zz_dataOut_payload_120_8;
  wire       [7:0]    _zz_dataOut_payload_120_9;
  wire       [7:0]    _zz_dataOut_payload_124;
  wire                _zz_dataOut_payload_120_10;
  wire       [7:0]    _zz_dataOut_payload_120_11;
  wire       [7:0]    _zz_dataOut_payload_124_1;
  wire                _zz_dataOut_payload_120_12;
  wire       [7:0]    _zz_dataOut_payload_120_13;
  wire       [7:0]    _zz_dataOut_payload_124_2;
  wire                _zz_dataOut_payload_120_14;
  wire       [7:0]    _zz_dataOut_payload_120_15;
  wire       [7:0]    _zz_dataOut_payload_124_3;
  wire                _zz_dataOut_payload_120_16;
  wire       [7:0]    _zz_dataOut_payload_120_17;
  wire       [7:0]    _zz_dataOut_payload_122;
  wire                _zz_dataOut_payload_120_18;
  wire       [7:0]    _zz_dataOut_payload_120_19;
  wire       [7:0]    _zz_dataOut_payload_122_1;
  wire                _zz_dataOut_payload_120_20;
  wire                _zz_dataOut_payload_122_2;
  reg        [7:0]    _zz_dataOut_payload_120_21;
  reg        [7:0]    _zz_dataOut_payload_121;
  reg        [7:0]    _zz_dataOut_payload_122_3;
  reg        [7:0]    _zz_dataOut_payload_123;
  wire                _zz_dataOut_payload_124_4;
  wire       [7:0]    _zz_dataOut_payload_124_5;
  wire       [7:0]    _zz_dataOut_payload_126;
  wire                _zz_dataOut_payload_124_6;
  wire       [7:0]    _zz_dataOut_payload_124_7;
  wire       [7:0]    _zz_dataOut_payload_126_1;
  wire                _zz_dataOut_payload_124_8;
  wire                _zz_dataOut_payload_126_2;
  reg        [7:0]    _zz_dataOut_payload_124_9;
  reg        [7:0]    _zz_dataOut_payload_125;
  reg        [7:0]    _zz_dataOut_payload_126_3;
  reg        [7:0]    _zz_dataOut_payload_127;
  reg        [7:0]    _zz_dataOut_payload_120_22;
  reg        [7:0]    _zz_dataOut_payload_121_1;
  reg        [7:0]    _zz_dataOut_payload_122_4;
  reg        [7:0]    _zz_dataOut_payload_123_1;
  reg        [7:0]    _zz_dataOut_payload_124_10;
  reg        [7:0]    _zz_dataOut_payload_125_1;
  reg        [7:0]    _zz_dataOut_payload_126_4;
  reg        [7:0]    _zz_dataOut_payload_127_1;
  reg        [7:0]    _zz_dataOut_payload_112_47;
  reg        [7:0]    _zz_dataOut_payload_113_2;
  reg        [7:0]    _zz_dataOut_payload_114_5;
  reg        [7:0]    _zz_dataOut_payload_115_2;
  reg        [7:0]    _zz_dataOut_payload_116_11;
  reg        [7:0]    _zz_dataOut_payload_117_2;
  reg        [7:0]    _zz_dataOut_payload_118_5;
  reg        [7:0]    _zz_dataOut_payload_119_2;
  reg        [7:0]    _zz_dataOut_payload_120_23;
  reg        [7:0]    _zz_dataOut_payload_121_2;
  reg        [7:0]    _zz_dataOut_payload_122_5;
  reg        [7:0]    _zz_dataOut_payload_123_2;
  reg        [7:0]    _zz_dataOut_payload_124_11;
  reg        [7:0]    _zz_dataOut_payload_125_2;
  reg        [7:0]    _zz_dataOut_payload_126_5;
  reg        [7:0]    _zz_dataOut_payload_127_2;
  reg        [7:0]    _zz_dataOut_payload_96_96;
  reg        [7:0]    _zz_dataOut_payload_97_3;
  reg        [7:0]    _zz_dataOut_payload_98_6;
  reg        [7:0]    _zz_dataOut_payload_99_3;
  reg        [7:0]    _zz_dataOut_payload_100_12;
  reg        [7:0]    _zz_dataOut_payload_101_3;
  reg        [7:0]    _zz_dataOut_payload_102_6;
  reg        [7:0]    _zz_dataOut_payload_103_3;
  reg        [7:0]    _zz_dataOut_payload_104_24;
  reg        [7:0]    _zz_dataOut_payload_105_3;
  reg        [7:0]    _zz_dataOut_payload_106_6;
  reg        [7:0]    _zz_dataOut_payload_107_3;
  reg        [7:0]    _zz_dataOut_payload_108_12;
  reg        [7:0]    _zz_dataOut_payload_109_3;
  reg        [7:0]    _zz_dataOut_payload_110_6;
  reg        [7:0]    _zz_dataOut_payload_111_3;
  reg        [7:0]    _zz_dataOut_payload_112_48;
  reg        [7:0]    _zz_dataOut_payload_113_3;
  reg        [7:0]    _zz_dataOut_payload_114_6;
  reg        [7:0]    _zz_dataOut_payload_115_3;
  reg        [7:0]    _zz_dataOut_payload_116_12;
  reg        [7:0]    _zz_dataOut_payload_117_3;
  reg        [7:0]    _zz_dataOut_payload_118_6;
  reg        [7:0]    _zz_dataOut_payload_119_3;
  reg        [7:0]    _zz_dataOut_payload_120_24;
  reg        [7:0]    _zz_dataOut_payload_121_3;
  reg        [7:0]    _zz_dataOut_payload_122_6;
  reg        [7:0]    _zz_dataOut_payload_123_3;
  reg        [7:0]    _zz_dataOut_payload_124_12;
  reg        [7:0]    _zz_dataOut_payload_125_3;
  reg        [7:0]    _zz_dataOut_payload_126_6;
  reg        [7:0]    _zz_dataOut_payload_127_3;
  reg        [7:0]    _zz_dataOut_payload_64_193;
  reg        [7:0]    _zz_dataOut_payload_65_4;
  reg        [7:0]    _zz_dataOut_payload_66_7;
  reg        [7:0]    _zz_dataOut_payload_67_4;
  reg        [7:0]    _zz_dataOut_payload_68_13;
  reg        [7:0]    _zz_dataOut_payload_69_4;
  reg        [7:0]    _zz_dataOut_payload_70_7;
  reg        [7:0]    _zz_dataOut_payload_71_4;
  reg        [7:0]    _zz_dataOut_payload_72_25;
  reg        [7:0]    _zz_dataOut_payload_73_4;
  reg        [7:0]    _zz_dataOut_payload_74_7;
  reg        [7:0]    _zz_dataOut_payload_75_4;
  reg        [7:0]    _zz_dataOut_payload_76_13;
  reg        [7:0]    _zz_dataOut_payload_77_4;
  reg        [7:0]    _zz_dataOut_payload_78_7;
  reg        [7:0]    _zz_dataOut_payload_79_4;
  reg        [7:0]    _zz_dataOut_payload_80_49;
  reg        [7:0]    _zz_dataOut_payload_81_4;
  reg        [7:0]    _zz_dataOut_payload_82_7;
  reg        [7:0]    _zz_dataOut_payload_83_4;
  reg        [7:0]    _zz_dataOut_payload_84_13;
  reg        [7:0]    _zz_dataOut_payload_85_4;
  reg        [7:0]    _zz_dataOut_payload_86_7;
  reg        [7:0]    _zz_dataOut_payload_87_4;
  reg        [7:0]    _zz_dataOut_payload_88_25;
  reg        [7:0]    _zz_dataOut_payload_89_4;
  reg        [7:0]    _zz_dataOut_payload_90_7;
  reg        [7:0]    _zz_dataOut_payload_91_4;
  reg        [7:0]    _zz_dataOut_payload_92_13;
  reg        [7:0]    _zz_dataOut_payload_93_4;
  reg        [7:0]    _zz_dataOut_payload_94_7;
  reg        [7:0]    _zz_dataOut_payload_95_4;
  reg        [7:0]    _zz_dataOut_payload_96_97;
  reg        [7:0]    _zz_dataOut_payload_97_4;
  reg        [7:0]    _zz_dataOut_payload_98_7;
  reg        [7:0]    _zz_dataOut_payload_99_4;
  reg        [7:0]    _zz_dataOut_payload_100_13;
  reg        [7:0]    _zz_dataOut_payload_101_4;
  reg        [7:0]    _zz_dataOut_payload_102_7;
  reg        [7:0]    _zz_dataOut_payload_103_4;
  reg        [7:0]    _zz_dataOut_payload_104_25;
  reg        [7:0]    _zz_dataOut_payload_105_4;
  reg        [7:0]    _zz_dataOut_payload_106_7;
  reg        [7:0]    _zz_dataOut_payload_107_4;
  reg        [7:0]    _zz_dataOut_payload_108_13;
  reg        [7:0]    _zz_dataOut_payload_109_4;
  reg        [7:0]    _zz_dataOut_payload_110_7;
  reg        [7:0]    _zz_dataOut_payload_111_4;
  reg        [7:0]    _zz_dataOut_payload_112_49;
  reg        [7:0]    _zz_dataOut_payload_113_4;
  reg        [7:0]    _zz_dataOut_payload_114_7;
  reg        [7:0]    _zz_dataOut_payload_115_4;
  reg        [7:0]    _zz_dataOut_payload_116_13;
  reg        [7:0]    _zz_dataOut_payload_117_4;
  reg        [7:0]    _zz_dataOut_payload_118_7;
  reg        [7:0]    _zz_dataOut_payload_119_4;
  reg        [7:0]    _zz_dataOut_payload_120_25;
  reg        [7:0]    _zz_dataOut_payload_121_4;
  reg        [7:0]    _zz_dataOut_payload_122_7;
  reg        [7:0]    _zz_dataOut_payload_123_4;
  reg        [7:0]    _zz_dataOut_payload_124_13;
  reg        [7:0]    _zz_dataOut_payload_125_4;
  reg        [7:0]    _zz_dataOut_payload_126_7;
  reg        [7:0]    _zz_dataOut_payload_127_4;
  reg        [7:0]    _zz_dataOut_payload_0_16642;
  reg        [7:0]    _zz_dataOut_payload_1_5;
  reg        [7:0]    _zz_dataOut_payload_2_8;
  reg        [7:0]    _zz_dataOut_payload_3_5;
  reg        [7:0]    _zz_dataOut_payload_4_14;
  reg        [7:0]    _zz_dataOut_payload_5_5;
  reg        [7:0]    _zz_dataOut_payload_6_8;
  reg        [7:0]    _zz_dataOut_payload_7_5;
  reg        [7:0]    _zz_dataOut_payload_8_26;
  reg        [7:0]    _zz_dataOut_payload_9_5;
  reg        [7:0]    _zz_dataOut_payload_10_8;
  reg        [7:0]    _zz_dataOut_payload_11_5;
  reg        [7:0]    _zz_dataOut_payload_12_14;
  reg        [7:0]    _zz_dataOut_payload_13_5;
  reg        [7:0]    _zz_dataOut_payload_14_8;
  reg        [7:0]    _zz_dataOut_payload_15_5;
  reg        [7:0]    _zz_dataOut_payload_16_50;
  reg        [7:0]    _zz_dataOut_payload_17_5;
  reg        [7:0]    _zz_dataOut_payload_18_8;
  reg        [7:0]    _zz_dataOut_payload_19_5;
  reg        [7:0]    _zz_dataOut_payload_20_14;
  reg        [7:0]    _zz_dataOut_payload_21_5;
  reg        [7:0]    _zz_dataOut_payload_22_8;
  reg        [7:0]    _zz_dataOut_payload_23_5;
  reg        [7:0]    _zz_dataOut_payload_24_26;
  reg        [7:0]    _zz_dataOut_payload_25_5;
  reg        [7:0]    _zz_dataOut_payload_26_8;
  reg        [7:0]    _zz_dataOut_payload_27_5;
  reg        [7:0]    _zz_dataOut_payload_28_14;
  reg        [7:0]    _zz_dataOut_payload_29_5;
  reg        [7:0]    _zz_dataOut_payload_30_8;
  reg        [7:0]    _zz_dataOut_payload_31_5;
  reg        [7:0]    _zz_dataOut_payload_32_98;
  reg        [7:0]    _zz_dataOut_payload_33_5;
  reg        [7:0]    _zz_dataOut_payload_34_8;
  reg        [7:0]    _zz_dataOut_payload_35_5;
  reg        [7:0]    _zz_dataOut_payload_36_14;
  reg        [7:0]    _zz_dataOut_payload_37_5;
  reg        [7:0]    _zz_dataOut_payload_38_8;
  reg        [7:0]    _zz_dataOut_payload_39_5;
  reg        [7:0]    _zz_dataOut_payload_40_26;
  reg        [7:0]    _zz_dataOut_payload_41_5;
  reg        [7:0]    _zz_dataOut_payload_42_8;
  reg        [7:0]    _zz_dataOut_payload_43_5;
  reg        [7:0]    _zz_dataOut_payload_44_14;
  reg        [7:0]    _zz_dataOut_payload_45_5;
  reg        [7:0]    _zz_dataOut_payload_46_8;
  reg        [7:0]    _zz_dataOut_payload_47_5;
  reg        [7:0]    _zz_dataOut_payload_48_50;
  reg        [7:0]    _zz_dataOut_payload_49_5;
  reg        [7:0]    _zz_dataOut_payload_50_8;
  reg        [7:0]    _zz_dataOut_payload_51_5;
  reg        [7:0]    _zz_dataOut_payload_52_14;
  reg        [7:0]    _zz_dataOut_payload_53_5;
  reg        [7:0]    _zz_dataOut_payload_54_8;
  reg        [7:0]    _zz_dataOut_payload_55_5;
  reg        [7:0]    _zz_dataOut_payload_56_26;
  reg        [7:0]    _zz_dataOut_payload_57_5;
  reg        [7:0]    _zz_dataOut_payload_58_8;
  reg        [7:0]    _zz_dataOut_payload_59_5;
  reg        [7:0]    _zz_dataOut_payload_60_14;
  reg        [7:0]    _zz_dataOut_payload_61_5;
  reg        [7:0]    _zz_dataOut_payload_62_8;
  reg        [7:0]    _zz_dataOut_payload_63_5;
  reg        [7:0]    _zz_dataOut_payload_64_194;
  reg        [7:0]    _zz_dataOut_payload_65_5;
  reg        [7:0]    _zz_dataOut_payload_66_8;
  reg        [7:0]    _zz_dataOut_payload_67_5;
  reg        [7:0]    _zz_dataOut_payload_68_14;
  reg        [7:0]    _zz_dataOut_payload_69_5;
  reg        [7:0]    _zz_dataOut_payload_70_8;
  reg        [7:0]    _zz_dataOut_payload_71_5;
  reg        [7:0]    _zz_dataOut_payload_72_26;
  reg        [7:0]    _zz_dataOut_payload_73_5;
  reg        [7:0]    _zz_dataOut_payload_74_8;
  reg        [7:0]    _zz_dataOut_payload_75_5;
  reg        [7:0]    _zz_dataOut_payload_76_14;
  reg        [7:0]    _zz_dataOut_payload_77_5;
  reg        [7:0]    _zz_dataOut_payload_78_8;
  reg        [7:0]    _zz_dataOut_payload_79_5;
  reg        [7:0]    _zz_dataOut_payload_80_50;
  reg        [7:0]    _zz_dataOut_payload_81_5;
  reg        [7:0]    _zz_dataOut_payload_82_8;
  reg        [7:0]    _zz_dataOut_payload_83_5;
  reg        [7:0]    _zz_dataOut_payload_84_14;
  reg        [7:0]    _zz_dataOut_payload_85_5;
  reg        [7:0]    _zz_dataOut_payload_86_8;
  reg        [7:0]    _zz_dataOut_payload_87_5;
  reg        [7:0]    _zz_dataOut_payload_88_26;
  reg        [7:0]    _zz_dataOut_payload_89_5;
  reg        [7:0]    _zz_dataOut_payload_90_8;
  reg        [7:0]    _zz_dataOut_payload_91_5;
  reg        [7:0]    _zz_dataOut_payload_92_14;
  reg        [7:0]    _zz_dataOut_payload_93_5;
  reg        [7:0]    _zz_dataOut_payload_94_8;
  reg        [7:0]    _zz_dataOut_payload_95_5;
  reg        [7:0]    _zz_dataOut_payload_96_98;
  reg        [7:0]    _zz_dataOut_payload_97_5;
  reg        [7:0]    _zz_dataOut_payload_98_8;
  reg        [7:0]    _zz_dataOut_payload_99_5;
  reg        [7:0]    _zz_dataOut_payload_100_14;
  reg        [7:0]    _zz_dataOut_payload_101_5;
  reg        [7:0]    _zz_dataOut_payload_102_8;
  reg        [7:0]    _zz_dataOut_payload_103_5;
  reg        [7:0]    _zz_dataOut_payload_104_26;
  reg        [7:0]    _zz_dataOut_payload_105_5;
  reg        [7:0]    _zz_dataOut_payload_106_8;
  reg        [7:0]    _zz_dataOut_payload_107_5;
  reg        [7:0]    _zz_dataOut_payload_108_14;
  reg        [7:0]    _zz_dataOut_payload_109_5;
  reg        [7:0]    _zz_dataOut_payload_110_8;
  reg        [7:0]    _zz_dataOut_payload_111_5;
  reg        [7:0]    _zz_dataOut_payload_112_50;
  reg        [7:0]    _zz_dataOut_payload_113_5;
  reg        [7:0]    _zz_dataOut_payload_114_8;
  reg        [7:0]    _zz_dataOut_payload_115_5;
  reg        [7:0]    _zz_dataOut_payload_116_14;
  reg        [7:0]    _zz_dataOut_payload_117_5;
  reg        [7:0]    _zz_dataOut_payload_118_8;
  reg        [7:0]    _zz_dataOut_payload_119_5;
  reg        [7:0]    _zz_dataOut_payload_120_26;
  reg        [7:0]    _zz_dataOut_payload_121_5;
  reg        [7:0]    _zz_dataOut_payload_122_8;
  reg        [7:0]    _zz_dataOut_payload_123_5;
  reg        [7:0]    _zz_dataOut_payload_124_14;
  reg        [7:0]    _zz_dataOut_payload_125_5;
  reg        [7:0]    _zz_dataOut_payload_126_8;
  reg        [7:0]    _zz_dataOut_payload_127_5;
  wire                _zz_dataOut_payload_128_128;
  wire       [7:0]    _zz_dataOut_payload_128_129;
  wire       [7:0]    _zz_dataOut_payload_192;
  wire                _zz_dataOut_payload_128_130;
  wire       [7:0]    _zz_dataOut_payload_128_131;
  wire       [7:0]    _zz_dataOut_payload_192_1;
  wire                _zz_dataOut_payload_128_132;
  wire       [7:0]    _zz_dataOut_payload_128_133;
  wire       [7:0]    _zz_dataOut_payload_192_2;
  wire                _zz_dataOut_payload_128_134;
  wire       [7:0]    _zz_dataOut_payload_128_135;
  wire       [7:0]    _zz_dataOut_payload_192_3;
  wire                _zz_dataOut_payload_128_136;
  wire       [7:0]    _zz_dataOut_payload_128_137;
  wire       [7:0]    _zz_dataOut_payload_192_4;
  wire                _zz_dataOut_payload_128_138;
  wire       [7:0]    _zz_dataOut_payload_128_139;
  wire       [7:0]    _zz_dataOut_payload_192_5;
  wire                _zz_dataOut_payload_128_140;
  wire       [7:0]    _zz_dataOut_payload_128_141;
  wire       [7:0]    _zz_dataOut_payload_192_6;
  wire                _zz_dataOut_payload_128_142;
  wire       [7:0]    _zz_dataOut_payload_128_143;
  wire       [7:0]    _zz_dataOut_payload_192_7;
  wire                _zz_dataOut_payload_128_144;
  wire       [7:0]    _zz_dataOut_payload_128_145;
  wire       [7:0]    _zz_dataOut_payload_192_8;
  wire                _zz_dataOut_payload_128_146;
  wire       [7:0]    _zz_dataOut_payload_128_147;
  wire       [7:0]    _zz_dataOut_payload_192_9;
  wire                _zz_dataOut_payload_128_148;
  wire       [7:0]    _zz_dataOut_payload_128_149;
  wire       [7:0]    _zz_dataOut_payload_192_10;
  wire                _zz_dataOut_payload_128_150;
  wire       [7:0]    _zz_dataOut_payload_128_151;
  wire       [7:0]    _zz_dataOut_payload_192_11;
  wire                _zz_dataOut_payload_128_152;
  wire       [7:0]    _zz_dataOut_payload_128_153;
  wire       [7:0]    _zz_dataOut_payload_192_12;
  wire                _zz_dataOut_payload_128_154;
  wire       [7:0]    _zz_dataOut_payload_128_155;
  wire       [7:0]    _zz_dataOut_payload_192_13;
  wire                _zz_dataOut_payload_128_156;
  wire       [7:0]    _zz_dataOut_payload_128_157;
  wire       [7:0]    _zz_dataOut_payload_192_14;
  wire                _zz_dataOut_payload_128_158;
  wire       [7:0]    _zz_dataOut_payload_128_159;
  wire       [7:0]    _zz_dataOut_payload_192_15;
  wire                _zz_dataOut_payload_128_160;
  wire       [7:0]    _zz_dataOut_payload_128_161;
  wire       [7:0]    _zz_dataOut_payload_192_16;
  wire                _zz_dataOut_payload_128_162;
  wire       [7:0]    _zz_dataOut_payload_128_163;
  wire       [7:0]    _zz_dataOut_payload_192_17;
  wire                _zz_dataOut_payload_128_164;
  wire       [7:0]    _zz_dataOut_payload_128_165;
  wire       [7:0]    _zz_dataOut_payload_192_18;
  wire                _zz_dataOut_payload_128_166;
  wire       [7:0]    _zz_dataOut_payload_128_167;
  wire       [7:0]    _zz_dataOut_payload_192_19;
  wire                _zz_dataOut_payload_128_168;
  wire       [7:0]    _zz_dataOut_payload_128_169;
  wire       [7:0]    _zz_dataOut_payload_192_20;
  wire                _zz_dataOut_payload_128_170;
  wire       [7:0]    _zz_dataOut_payload_128_171;
  wire       [7:0]    _zz_dataOut_payload_192_21;
  wire                _zz_dataOut_payload_128_172;
  wire       [7:0]    _zz_dataOut_payload_128_173;
  wire       [7:0]    _zz_dataOut_payload_192_22;
  wire                _zz_dataOut_payload_128_174;
  wire       [7:0]    _zz_dataOut_payload_128_175;
  wire       [7:0]    _zz_dataOut_payload_192_23;
  wire                _zz_dataOut_payload_128_176;
  wire       [7:0]    _zz_dataOut_payload_128_177;
  wire       [7:0]    _zz_dataOut_payload_192_24;
  wire                _zz_dataOut_payload_128_178;
  wire       [7:0]    _zz_dataOut_payload_128_179;
  wire       [7:0]    _zz_dataOut_payload_192_25;
  wire                _zz_dataOut_payload_128_180;
  wire       [7:0]    _zz_dataOut_payload_128_181;
  wire       [7:0]    _zz_dataOut_payload_192_26;
  wire                _zz_dataOut_payload_128_182;
  wire       [7:0]    _zz_dataOut_payload_128_183;
  wire       [7:0]    _zz_dataOut_payload_192_27;
  wire                _zz_dataOut_payload_128_184;
  wire       [7:0]    _zz_dataOut_payload_128_185;
  wire       [7:0]    _zz_dataOut_payload_192_28;
  wire                _zz_dataOut_payload_128_186;
  wire       [7:0]    _zz_dataOut_payload_128_187;
  wire       [7:0]    _zz_dataOut_payload_192_29;
  wire                _zz_dataOut_payload_128_188;
  wire       [7:0]    _zz_dataOut_payload_128_189;
  wire       [7:0]    _zz_dataOut_payload_192_30;
  wire                _zz_dataOut_payload_128_190;
  wire       [7:0]    _zz_dataOut_payload_128_191;
  wire       [7:0]    _zz_dataOut_payload_192_31;
  wire                _zz_dataOut_payload_128_192;
  wire       [7:0]    _zz_dataOut_payload_128_193;
  wire       [7:0]    _zz_dataOut_payload_192_32;
  wire                _zz_dataOut_payload_128_194;
  wire       [7:0]    _zz_dataOut_payload_128_195;
  wire       [7:0]    _zz_dataOut_payload_192_33;
  wire                _zz_dataOut_payload_128_196;
  wire       [7:0]    _zz_dataOut_payload_128_197;
  wire       [7:0]    _zz_dataOut_payload_192_34;
  wire                _zz_dataOut_payload_128_198;
  wire       [7:0]    _zz_dataOut_payload_128_199;
  wire       [7:0]    _zz_dataOut_payload_192_35;
  wire                _zz_dataOut_payload_128_200;
  wire       [7:0]    _zz_dataOut_payload_128_201;
  wire       [7:0]    _zz_dataOut_payload_192_36;
  wire                _zz_dataOut_payload_128_202;
  wire       [7:0]    _zz_dataOut_payload_128_203;
  wire       [7:0]    _zz_dataOut_payload_192_37;
  wire                _zz_dataOut_payload_128_204;
  wire       [7:0]    _zz_dataOut_payload_128_205;
  wire       [7:0]    _zz_dataOut_payload_192_38;
  wire                _zz_dataOut_payload_128_206;
  wire       [7:0]    _zz_dataOut_payload_128_207;
  wire       [7:0]    _zz_dataOut_payload_192_39;
  wire                _zz_dataOut_payload_128_208;
  wire       [7:0]    _zz_dataOut_payload_128_209;
  wire       [7:0]    _zz_dataOut_payload_192_40;
  wire                _zz_dataOut_payload_128_210;
  wire       [7:0]    _zz_dataOut_payload_128_211;
  wire       [7:0]    _zz_dataOut_payload_192_41;
  wire                _zz_dataOut_payload_128_212;
  wire       [7:0]    _zz_dataOut_payload_128_213;
  wire       [7:0]    _zz_dataOut_payload_192_42;
  wire                _zz_dataOut_payload_128_214;
  wire       [7:0]    _zz_dataOut_payload_128_215;
  wire       [7:0]    _zz_dataOut_payload_192_43;
  wire                _zz_dataOut_payload_128_216;
  wire       [7:0]    _zz_dataOut_payload_128_217;
  wire       [7:0]    _zz_dataOut_payload_192_44;
  wire                _zz_dataOut_payload_128_218;
  wire       [7:0]    _zz_dataOut_payload_128_219;
  wire       [7:0]    _zz_dataOut_payload_192_45;
  wire                _zz_dataOut_payload_128_220;
  wire       [7:0]    _zz_dataOut_payload_128_221;
  wire       [7:0]    _zz_dataOut_payload_192_46;
  wire                _zz_dataOut_payload_128_222;
  wire       [7:0]    _zz_dataOut_payload_128_223;
  wire       [7:0]    _zz_dataOut_payload_192_47;
  wire                _zz_dataOut_payload_128_224;
  wire       [7:0]    _zz_dataOut_payload_128_225;
  wire       [7:0]    _zz_dataOut_payload_192_48;
  wire                _zz_dataOut_payload_128_226;
  wire       [7:0]    _zz_dataOut_payload_128_227;
  wire       [7:0]    _zz_dataOut_payload_192_49;
  wire                _zz_dataOut_payload_128_228;
  wire       [7:0]    _zz_dataOut_payload_128_229;
  wire       [7:0]    _zz_dataOut_payload_192_50;
  wire                _zz_dataOut_payload_128_230;
  wire       [7:0]    _zz_dataOut_payload_128_231;
  wire       [7:0]    _zz_dataOut_payload_192_51;
  wire                _zz_dataOut_payload_128_232;
  wire       [7:0]    _zz_dataOut_payload_128_233;
  wire       [7:0]    _zz_dataOut_payload_192_52;
  wire                _zz_dataOut_payload_128_234;
  wire       [7:0]    _zz_dataOut_payload_128_235;
  wire       [7:0]    _zz_dataOut_payload_192_53;
  wire                _zz_dataOut_payload_128_236;
  wire       [7:0]    _zz_dataOut_payload_128_237;
  wire       [7:0]    _zz_dataOut_payload_192_54;
  wire                _zz_dataOut_payload_128_238;
  wire       [7:0]    _zz_dataOut_payload_128_239;
  wire       [7:0]    _zz_dataOut_payload_192_55;
  wire                _zz_dataOut_payload_128_240;
  wire       [7:0]    _zz_dataOut_payload_128_241;
  wire       [7:0]    _zz_dataOut_payload_192_56;
  wire                _zz_dataOut_payload_128_242;
  wire       [7:0]    _zz_dataOut_payload_128_243;
  wire       [7:0]    _zz_dataOut_payload_192_57;
  wire                _zz_dataOut_payload_128_244;
  wire       [7:0]    _zz_dataOut_payload_128_245;
  wire       [7:0]    _zz_dataOut_payload_192_58;
  wire                _zz_dataOut_payload_128_246;
  wire       [7:0]    _zz_dataOut_payload_128_247;
  wire       [7:0]    _zz_dataOut_payload_192_59;
  wire                _zz_dataOut_payload_128_248;
  wire       [7:0]    _zz_dataOut_payload_128_249;
  wire       [7:0]    _zz_dataOut_payload_192_60;
  wire                _zz_dataOut_payload_128_250;
  wire       [7:0]    _zz_dataOut_payload_128_251;
  wire       [7:0]    _zz_dataOut_payload_192_61;
  wire                _zz_dataOut_payload_128_252;
  wire       [7:0]    _zz_dataOut_payload_128_253;
  wire       [7:0]    _zz_dataOut_payload_192_62;
  wire                _zz_dataOut_payload_128_254;
  wire       [7:0]    _zz_dataOut_payload_128_255;
  wire       [7:0]    _zz_dataOut_payload_192_63;
  wire                _zz_dataOut_payload_128_256;
  wire       [7:0]    _zz_dataOut_payload_128_257;
  wire       [7:0]    _zz_dataOut_payload_160;
  wire                _zz_dataOut_payload_128_258;
  wire       [7:0]    _zz_dataOut_payload_128_259;
  wire       [7:0]    _zz_dataOut_payload_160_1;
  wire                _zz_dataOut_payload_128_260;
  wire       [7:0]    _zz_dataOut_payload_128_261;
  wire       [7:0]    _zz_dataOut_payload_160_2;
  wire                _zz_dataOut_payload_128_262;
  wire       [7:0]    _zz_dataOut_payload_128_263;
  wire       [7:0]    _zz_dataOut_payload_160_3;
  wire                _zz_dataOut_payload_128_264;
  wire       [7:0]    _zz_dataOut_payload_128_265;
  wire       [7:0]    _zz_dataOut_payload_160_4;
  wire                _zz_dataOut_payload_128_266;
  wire       [7:0]    _zz_dataOut_payload_128_267;
  wire       [7:0]    _zz_dataOut_payload_160_5;
  wire                _zz_dataOut_payload_128_268;
  wire       [7:0]    _zz_dataOut_payload_128_269;
  wire       [7:0]    _zz_dataOut_payload_160_6;
  wire                _zz_dataOut_payload_128_270;
  wire       [7:0]    _zz_dataOut_payload_128_271;
  wire       [7:0]    _zz_dataOut_payload_160_7;
  wire                _zz_dataOut_payload_128_272;
  wire       [7:0]    _zz_dataOut_payload_128_273;
  wire       [7:0]    _zz_dataOut_payload_160_8;
  wire                _zz_dataOut_payload_128_274;
  wire       [7:0]    _zz_dataOut_payload_128_275;
  wire       [7:0]    _zz_dataOut_payload_160_9;
  wire                _zz_dataOut_payload_128_276;
  wire       [7:0]    _zz_dataOut_payload_128_277;
  wire       [7:0]    _zz_dataOut_payload_160_10;
  wire                _zz_dataOut_payload_128_278;
  wire       [7:0]    _zz_dataOut_payload_128_279;
  wire       [7:0]    _zz_dataOut_payload_160_11;
  wire                _zz_dataOut_payload_128_280;
  wire       [7:0]    _zz_dataOut_payload_128_281;
  wire       [7:0]    _zz_dataOut_payload_160_12;
  wire                _zz_dataOut_payload_128_282;
  wire       [7:0]    _zz_dataOut_payload_128_283;
  wire       [7:0]    _zz_dataOut_payload_160_13;
  wire                _zz_dataOut_payload_128_284;
  wire       [7:0]    _zz_dataOut_payload_128_285;
  wire       [7:0]    _zz_dataOut_payload_160_14;
  wire                _zz_dataOut_payload_128_286;
  wire       [7:0]    _zz_dataOut_payload_128_287;
  wire       [7:0]    _zz_dataOut_payload_160_15;
  wire                _zz_dataOut_payload_128_288;
  wire       [7:0]    _zz_dataOut_payload_128_289;
  wire       [7:0]    _zz_dataOut_payload_160_16;
  wire                _zz_dataOut_payload_128_290;
  wire       [7:0]    _zz_dataOut_payload_128_291;
  wire       [7:0]    _zz_dataOut_payload_160_17;
  wire                _zz_dataOut_payload_128_292;
  wire       [7:0]    _zz_dataOut_payload_128_293;
  wire       [7:0]    _zz_dataOut_payload_160_18;
  wire                _zz_dataOut_payload_128_294;
  wire       [7:0]    _zz_dataOut_payload_128_295;
  wire       [7:0]    _zz_dataOut_payload_160_19;
  wire                _zz_dataOut_payload_128_296;
  wire       [7:0]    _zz_dataOut_payload_128_297;
  wire       [7:0]    _zz_dataOut_payload_160_20;
  wire                _zz_dataOut_payload_128_298;
  wire       [7:0]    _zz_dataOut_payload_128_299;
  wire       [7:0]    _zz_dataOut_payload_160_21;
  wire                _zz_dataOut_payload_128_300;
  wire       [7:0]    _zz_dataOut_payload_128_301;
  wire       [7:0]    _zz_dataOut_payload_160_22;
  wire                _zz_dataOut_payload_128_302;
  wire       [7:0]    _zz_dataOut_payload_128_303;
  wire       [7:0]    _zz_dataOut_payload_160_23;
  wire                _zz_dataOut_payload_128_304;
  wire       [7:0]    _zz_dataOut_payload_128_305;
  wire       [7:0]    _zz_dataOut_payload_160_24;
  wire                _zz_dataOut_payload_128_306;
  wire       [7:0]    _zz_dataOut_payload_128_307;
  wire       [7:0]    _zz_dataOut_payload_160_25;
  wire                _zz_dataOut_payload_128_308;
  wire       [7:0]    _zz_dataOut_payload_128_309;
  wire       [7:0]    _zz_dataOut_payload_160_26;
  wire                _zz_dataOut_payload_128_310;
  wire       [7:0]    _zz_dataOut_payload_128_311;
  wire       [7:0]    _zz_dataOut_payload_160_27;
  wire                _zz_dataOut_payload_128_312;
  wire       [7:0]    _zz_dataOut_payload_128_313;
  wire       [7:0]    _zz_dataOut_payload_160_28;
  wire                _zz_dataOut_payload_128_314;
  wire       [7:0]    _zz_dataOut_payload_128_315;
  wire       [7:0]    _zz_dataOut_payload_160_29;
  wire                _zz_dataOut_payload_128_316;
  wire       [7:0]    _zz_dataOut_payload_128_317;
  wire       [7:0]    _zz_dataOut_payload_160_30;
  wire                _zz_dataOut_payload_128_318;
  wire       [7:0]    _zz_dataOut_payload_128_319;
  wire       [7:0]    _zz_dataOut_payload_160_31;
  wire                _zz_dataOut_payload_128_320;
  wire       [7:0]    _zz_dataOut_payload_128_321;
  wire       [7:0]    _zz_dataOut_payload_144;
  wire                _zz_dataOut_payload_128_322;
  wire       [7:0]    _zz_dataOut_payload_128_323;
  wire       [7:0]    _zz_dataOut_payload_144_1;
  wire                _zz_dataOut_payload_128_324;
  wire       [7:0]    _zz_dataOut_payload_128_325;
  wire       [7:0]    _zz_dataOut_payload_144_2;
  wire                _zz_dataOut_payload_128_326;
  wire       [7:0]    _zz_dataOut_payload_128_327;
  wire       [7:0]    _zz_dataOut_payload_144_3;
  wire                _zz_dataOut_payload_128_328;
  wire       [7:0]    _zz_dataOut_payload_128_329;
  wire       [7:0]    _zz_dataOut_payload_144_4;
  wire                _zz_dataOut_payload_128_330;
  wire       [7:0]    _zz_dataOut_payload_128_331;
  wire       [7:0]    _zz_dataOut_payload_144_5;
  wire                _zz_dataOut_payload_128_332;
  wire       [7:0]    _zz_dataOut_payload_128_333;
  wire       [7:0]    _zz_dataOut_payload_144_6;
  wire                _zz_dataOut_payload_128_334;
  wire       [7:0]    _zz_dataOut_payload_128_335;
  wire       [7:0]    _zz_dataOut_payload_144_7;
  wire                _zz_dataOut_payload_128_336;
  wire       [7:0]    _zz_dataOut_payload_128_337;
  wire       [7:0]    _zz_dataOut_payload_144_8;
  wire                _zz_dataOut_payload_128_338;
  wire       [7:0]    _zz_dataOut_payload_128_339;
  wire       [7:0]    _zz_dataOut_payload_144_9;
  wire                _zz_dataOut_payload_128_340;
  wire       [7:0]    _zz_dataOut_payload_128_341;
  wire       [7:0]    _zz_dataOut_payload_144_10;
  wire                _zz_dataOut_payload_128_342;
  wire       [7:0]    _zz_dataOut_payload_128_343;
  wire       [7:0]    _zz_dataOut_payload_144_11;
  wire                _zz_dataOut_payload_128_344;
  wire       [7:0]    _zz_dataOut_payload_128_345;
  wire       [7:0]    _zz_dataOut_payload_144_12;
  wire                _zz_dataOut_payload_128_346;
  wire       [7:0]    _zz_dataOut_payload_128_347;
  wire       [7:0]    _zz_dataOut_payload_144_13;
  wire                _zz_dataOut_payload_128_348;
  wire       [7:0]    _zz_dataOut_payload_128_349;
  wire       [7:0]    _zz_dataOut_payload_144_14;
  wire                _zz_dataOut_payload_128_350;
  wire       [7:0]    _zz_dataOut_payload_128_351;
  wire       [7:0]    _zz_dataOut_payload_144_15;
  wire                _zz_dataOut_payload_128_352;
  wire       [7:0]    _zz_dataOut_payload_128_353;
  wire       [7:0]    _zz_dataOut_payload_136;
  wire                _zz_dataOut_payload_128_354;
  wire       [7:0]    _zz_dataOut_payload_128_355;
  wire       [7:0]    _zz_dataOut_payload_136_1;
  wire                _zz_dataOut_payload_128_356;
  wire       [7:0]    _zz_dataOut_payload_128_357;
  wire       [7:0]    _zz_dataOut_payload_136_2;
  wire                _zz_dataOut_payload_128_358;
  wire       [7:0]    _zz_dataOut_payload_128_359;
  wire       [7:0]    _zz_dataOut_payload_136_3;
  wire                _zz_dataOut_payload_128_360;
  wire       [7:0]    _zz_dataOut_payload_128_361;
  wire       [7:0]    _zz_dataOut_payload_136_4;
  wire                _zz_dataOut_payload_128_362;
  wire       [7:0]    _zz_dataOut_payload_128_363;
  wire       [7:0]    _zz_dataOut_payload_136_5;
  wire                _zz_dataOut_payload_128_364;
  wire       [7:0]    _zz_dataOut_payload_128_365;
  wire       [7:0]    _zz_dataOut_payload_136_6;
  wire                _zz_dataOut_payload_128_366;
  wire       [7:0]    _zz_dataOut_payload_128_367;
  wire       [7:0]    _zz_dataOut_payload_136_7;
  wire                _zz_dataOut_payload_128_368;
  wire       [7:0]    _zz_dataOut_payload_128_369;
  wire       [7:0]    _zz_dataOut_payload_132;
  wire                _zz_dataOut_payload_128_370;
  wire       [7:0]    _zz_dataOut_payload_128_371;
  wire       [7:0]    _zz_dataOut_payload_132_1;
  wire                _zz_dataOut_payload_128_372;
  wire       [7:0]    _zz_dataOut_payload_128_373;
  wire       [7:0]    _zz_dataOut_payload_132_2;
  wire                _zz_dataOut_payload_128_374;
  wire       [7:0]    _zz_dataOut_payload_128_375;
  wire       [7:0]    _zz_dataOut_payload_132_3;
  wire                _zz_dataOut_payload_128_376;
  wire       [7:0]    _zz_dataOut_payload_128_377;
  wire       [7:0]    _zz_dataOut_payload_130;
  wire                _zz_dataOut_payload_128_378;
  wire       [7:0]    _zz_dataOut_payload_128_379;
  wire       [7:0]    _zz_dataOut_payload_130_1;
  wire                _zz_dataOut_payload_128_380;
  wire                _zz_dataOut_payload_130_2;
  reg        [7:0]    _zz_dataOut_payload_128_381;
  reg        [7:0]    _zz_dataOut_payload_129;
  reg        [7:0]    _zz_dataOut_payload_130_3;
  reg        [7:0]    _zz_dataOut_payload_131;
  wire                _zz_dataOut_payload_132_4;
  wire       [7:0]    _zz_dataOut_payload_132_5;
  wire       [7:0]    _zz_dataOut_payload_134;
  wire                _zz_dataOut_payload_132_6;
  wire       [7:0]    _zz_dataOut_payload_132_7;
  wire       [7:0]    _zz_dataOut_payload_134_1;
  wire                _zz_dataOut_payload_132_8;
  wire                _zz_dataOut_payload_134_2;
  reg        [7:0]    _zz_dataOut_payload_132_9;
  reg        [7:0]    _zz_dataOut_payload_133;
  reg        [7:0]    _zz_dataOut_payload_134_3;
  reg        [7:0]    _zz_dataOut_payload_135;
  reg        [7:0]    _zz_dataOut_payload_128_382;
  reg        [7:0]    _zz_dataOut_payload_129_1;
  reg        [7:0]    _zz_dataOut_payload_130_4;
  reg        [7:0]    _zz_dataOut_payload_131_1;
  reg        [7:0]    _zz_dataOut_payload_132_10;
  reg        [7:0]    _zz_dataOut_payload_133_1;
  reg        [7:0]    _zz_dataOut_payload_134_4;
  reg        [7:0]    _zz_dataOut_payload_135_1;
  wire                _zz_dataOut_payload_136_8;
  wire       [7:0]    _zz_dataOut_payload_136_9;
  wire       [7:0]    _zz_dataOut_payload_140;
  wire                _zz_dataOut_payload_136_10;
  wire       [7:0]    _zz_dataOut_payload_136_11;
  wire       [7:0]    _zz_dataOut_payload_140_1;
  wire                _zz_dataOut_payload_136_12;
  wire       [7:0]    _zz_dataOut_payload_136_13;
  wire       [7:0]    _zz_dataOut_payload_140_2;
  wire                _zz_dataOut_payload_136_14;
  wire       [7:0]    _zz_dataOut_payload_136_15;
  wire       [7:0]    _zz_dataOut_payload_140_3;
  wire                _zz_dataOut_payload_136_16;
  wire       [7:0]    _zz_dataOut_payload_136_17;
  wire       [7:0]    _zz_dataOut_payload_138;
  wire                _zz_dataOut_payload_136_18;
  wire       [7:0]    _zz_dataOut_payload_136_19;
  wire       [7:0]    _zz_dataOut_payload_138_1;
  wire                _zz_dataOut_payload_136_20;
  wire                _zz_dataOut_payload_138_2;
  reg        [7:0]    _zz_dataOut_payload_136_21;
  reg        [7:0]    _zz_dataOut_payload_137;
  reg        [7:0]    _zz_dataOut_payload_138_3;
  reg        [7:0]    _zz_dataOut_payload_139;
  wire                _zz_dataOut_payload_140_4;
  wire       [7:0]    _zz_dataOut_payload_140_5;
  wire       [7:0]    _zz_dataOut_payload_142;
  wire                _zz_dataOut_payload_140_6;
  wire       [7:0]    _zz_dataOut_payload_140_7;
  wire       [7:0]    _zz_dataOut_payload_142_1;
  wire                _zz_dataOut_payload_140_8;
  wire                _zz_dataOut_payload_142_2;
  reg        [7:0]    _zz_dataOut_payload_140_9;
  reg        [7:0]    _zz_dataOut_payload_141;
  reg        [7:0]    _zz_dataOut_payload_142_3;
  reg        [7:0]    _zz_dataOut_payload_143;
  reg        [7:0]    _zz_dataOut_payload_136_22;
  reg        [7:0]    _zz_dataOut_payload_137_1;
  reg        [7:0]    _zz_dataOut_payload_138_4;
  reg        [7:0]    _zz_dataOut_payload_139_1;
  reg        [7:0]    _zz_dataOut_payload_140_10;
  reg        [7:0]    _zz_dataOut_payload_141_1;
  reg        [7:0]    _zz_dataOut_payload_142_4;
  reg        [7:0]    _zz_dataOut_payload_143_1;
  reg        [7:0]    _zz_dataOut_payload_128_383;
  reg        [7:0]    _zz_dataOut_payload_129_2;
  reg        [7:0]    _zz_dataOut_payload_130_5;
  reg        [7:0]    _zz_dataOut_payload_131_2;
  reg        [7:0]    _zz_dataOut_payload_132_11;
  reg        [7:0]    _zz_dataOut_payload_133_2;
  reg        [7:0]    _zz_dataOut_payload_134_5;
  reg        [7:0]    _zz_dataOut_payload_135_2;
  reg        [7:0]    _zz_dataOut_payload_136_23;
  reg        [7:0]    _zz_dataOut_payload_137_2;
  reg        [7:0]    _zz_dataOut_payload_138_5;
  reg        [7:0]    _zz_dataOut_payload_139_2;
  reg        [7:0]    _zz_dataOut_payload_140_11;
  reg        [7:0]    _zz_dataOut_payload_141_2;
  reg        [7:0]    _zz_dataOut_payload_142_5;
  reg        [7:0]    _zz_dataOut_payload_143_2;
  wire                _zz_dataOut_payload_144_16;
  wire       [7:0]    _zz_dataOut_payload_144_17;
  wire       [7:0]    _zz_dataOut_payload_152;
  wire                _zz_dataOut_payload_144_18;
  wire       [7:0]    _zz_dataOut_payload_144_19;
  wire       [7:0]    _zz_dataOut_payload_152_1;
  wire                _zz_dataOut_payload_144_20;
  wire       [7:0]    _zz_dataOut_payload_144_21;
  wire       [7:0]    _zz_dataOut_payload_152_2;
  wire                _zz_dataOut_payload_144_22;
  wire       [7:0]    _zz_dataOut_payload_144_23;
  wire       [7:0]    _zz_dataOut_payload_152_3;
  wire                _zz_dataOut_payload_144_24;
  wire       [7:0]    _zz_dataOut_payload_144_25;
  wire       [7:0]    _zz_dataOut_payload_152_4;
  wire                _zz_dataOut_payload_144_26;
  wire       [7:0]    _zz_dataOut_payload_144_27;
  wire       [7:0]    _zz_dataOut_payload_152_5;
  wire                _zz_dataOut_payload_144_28;
  wire       [7:0]    _zz_dataOut_payload_144_29;
  wire       [7:0]    _zz_dataOut_payload_152_6;
  wire                _zz_dataOut_payload_144_30;
  wire       [7:0]    _zz_dataOut_payload_144_31;
  wire       [7:0]    _zz_dataOut_payload_152_7;
  wire                _zz_dataOut_payload_144_32;
  wire       [7:0]    _zz_dataOut_payload_144_33;
  wire       [7:0]    _zz_dataOut_payload_148;
  wire                _zz_dataOut_payload_144_34;
  wire       [7:0]    _zz_dataOut_payload_144_35;
  wire       [7:0]    _zz_dataOut_payload_148_1;
  wire                _zz_dataOut_payload_144_36;
  wire       [7:0]    _zz_dataOut_payload_144_37;
  wire       [7:0]    _zz_dataOut_payload_148_2;
  wire                _zz_dataOut_payload_144_38;
  wire       [7:0]    _zz_dataOut_payload_144_39;
  wire       [7:0]    _zz_dataOut_payload_148_3;
  wire                _zz_dataOut_payload_144_40;
  wire       [7:0]    _zz_dataOut_payload_144_41;
  wire       [7:0]    _zz_dataOut_payload_146;
  wire                _zz_dataOut_payload_144_42;
  wire       [7:0]    _zz_dataOut_payload_144_43;
  wire       [7:0]    _zz_dataOut_payload_146_1;
  wire                _zz_dataOut_payload_144_44;
  wire                _zz_dataOut_payload_146_2;
  reg        [7:0]    _zz_dataOut_payload_144_45;
  reg        [7:0]    _zz_dataOut_payload_145;
  reg        [7:0]    _zz_dataOut_payload_146_3;
  reg        [7:0]    _zz_dataOut_payload_147;
  wire                _zz_dataOut_payload_148_4;
  wire       [7:0]    _zz_dataOut_payload_148_5;
  wire       [7:0]    _zz_dataOut_payload_150;
  wire                _zz_dataOut_payload_148_6;
  wire       [7:0]    _zz_dataOut_payload_148_7;
  wire       [7:0]    _zz_dataOut_payload_150_1;
  wire                _zz_dataOut_payload_148_8;
  wire                _zz_dataOut_payload_150_2;
  reg        [7:0]    _zz_dataOut_payload_148_9;
  reg        [7:0]    _zz_dataOut_payload_149;
  reg        [7:0]    _zz_dataOut_payload_150_3;
  reg        [7:0]    _zz_dataOut_payload_151;
  reg        [7:0]    _zz_dataOut_payload_144_46;
  reg        [7:0]    _zz_dataOut_payload_145_1;
  reg        [7:0]    _zz_dataOut_payload_146_4;
  reg        [7:0]    _zz_dataOut_payload_147_1;
  reg        [7:0]    _zz_dataOut_payload_148_10;
  reg        [7:0]    _zz_dataOut_payload_149_1;
  reg        [7:0]    _zz_dataOut_payload_150_4;
  reg        [7:0]    _zz_dataOut_payload_151_1;
  wire                _zz_dataOut_payload_152_8;
  wire       [7:0]    _zz_dataOut_payload_152_9;
  wire       [7:0]    _zz_dataOut_payload_156;
  wire                _zz_dataOut_payload_152_10;
  wire       [7:0]    _zz_dataOut_payload_152_11;
  wire       [7:0]    _zz_dataOut_payload_156_1;
  wire                _zz_dataOut_payload_152_12;
  wire       [7:0]    _zz_dataOut_payload_152_13;
  wire       [7:0]    _zz_dataOut_payload_156_2;
  wire                _zz_dataOut_payload_152_14;
  wire       [7:0]    _zz_dataOut_payload_152_15;
  wire       [7:0]    _zz_dataOut_payload_156_3;
  wire                _zz_dataOut_payload_152_16;
  wire       [7:0]    _zz_dataOut_payload_152_17;
  wire       [7:0]    _zz_dataOut_payload_154;
  wire                _zz_dataOut_payload_152_18;
  wire       [7:0]    _zz_dataOut_payload_152_19;
  wire       [7:0]    _zz_dataOut_payload_154_1;
  wire                _zz_dataOut_payload_152_20;
  wire                _zz_dataOut_payload_154_2;
  reg        [7:0]    _zz_dataOut_payload_152_21;
  reg        [7:0]    _zz_dataOut_payload_153;
  reg        [7:0]    _zz_dataOut_payload_154_3;
  reg        [7:0]    _zz_dataOut_payload_155;
  wire                _zz_dataOut_payload_156_4;
  wire       [7:0]    _zz_dataOut_payload_156_5;
  wire       [7:0]    _zz_dataOut_payload_158;
  wire                _zz_dataOut_payload_156_6;
  wire       [7:0]    _zz_dataOut_payload_156_7;
  wire       [7:0]    _zz_dataOut_payload_158_1;
  wire                _zz_dataOut_payload_156_8;
  wire                _zz_dataOut_payload_158_2;
  reg        [7:0]    _zz_dataOut_payload_156_9;
  reg        [7:0]    _zz_dataOut_payload_157;
  reg        [7:0]    _zz_dataOut_payload_158_3;
  reg        [7:0]    _zz_dataOut_payload_159;
  reg        [7:0]    _zz_dataOut_payload_152_22;
  reg        [7:0]    _zz_dataOut_payload_153_1;
  reg        [7:0]    _zz_dataOut_payload_154_4;
  reg        [7:0]    _zz_dataOut_payload_155_1;
  reg        [7:0]    _zz_dataOut_payload_156_10;
  reg        [7:0]    _zz_dataOut_payload_157_1;
  reg        [7:0]    _zz_dataOut_payload_158_4;
  reg        [7:0]    _zz_dataOut_payload_159_1;
  reg        [7:0]    _zz_dataOut_payload_144_47;
  reg        [7:0]    _zz_dataOut_payload_145_2;
  reg        [7:0]    _zz_dataOut_payload_146_5;
  reg        [7:0]    _zz_dataOut_payload_147_2;
  reg        [7:0]    _zz_dataOut_payload_148_11;
  reg        [7:0]    _zz_dataOut_payload_149_2;
  reg        [7:0]    _zz_dataOut_payload_150_5;
  reg        [7:0]    _zz_dataOut_payload_151_2;
  reg        [7:0]    _zz_dataOut_payload_152_23;
  reg        [7:0]    _zz_dataOut_payload_153_2;
  reg        [7:0]    _zz_dataOut_payload_154_5;
  reg        [7:0]    _zz_dataOut_payload_155_2;
  reg        [7:0]    _zz_dataOut_payload_156_11;
  reg        [7:0]    _zz_dataOut_payload_157_2;
  reg        [7:0]    _zz_dataOut_payload_158_5;
  reg        [7:0]    _zz_dataOut_payload_159_2;
  reg        [7:0]    _zz_dataOut_payload_128_384;
  reg        [7:0]    _zz_dataOut_payload_129_3;
  reg        [7:0]    _zz_dataOut_payload_130_6;
  reg        [7:0]    _zz_dataOut_payload_131_3;
  reg        [7:0]    _zz_dataOut_payload_132_12;
  reg        [7:0]    _zz_dataOut_payload_133_3;
  reg        [7:0]    _zz_dataOut_payload_134_6;
  reg        [7:0]    _zz_dataOut_payload_135_3;
  reg        [7:0]    _zz_dataOut_payload_136_24;
  reg        [7:0]    _zz_dataOut_payload_137_3;
  reg        [7:0]    _zz_dataOut_payload_138_6;
  reg        [7:0]    _zz_dataOut_payload_139_3;
  reg        [7:0]    _zz_dataOut_payload_140_12;
  reg        [7:0]    _zz_dataOut_payload_141_3;
  reg        [7:0]    _zz_dataOut_payload_142_6;
  reg        [7:0]    _zz_dataOut_payload_143_3;
  reg        [7:0]    _zz_dataOut_payload_144_48;
  reg        [7:0]    _zz_dataOut_payload_145_3;
  reg        [7:0]    _zz_dataOut_payload_146_6;
  reg        [7:0]    _zz_dataOut_payload_147_3;
  reg        [7:0]    _zz_dataOut_payload_148_12;
  reg        [7:0]    _zz_dataOut_payload_149_3;
  reg        [7:0]    _zz_dataOut_payload_150_6;
  reg        [7:0]    _zz_dataOut_payload_151_3;
  reg        [7:0]    _zz_dataOut_payload_152_24;
  reg        [7:0]    _zz_dataOut_payload_153_3;
  reg        [7:0]    _zz_dataOut_payload_154_6;
  reg        [7:0]    _zz_dataOut_payload_155_3;
  reg        [7:0]    _zz_dataOut_payload_156_12;
  reg        [7:0]    _zz_dataOut_payload_157_3;
  reg        [7:0]    _zz_dataOut_payload_158_6;
  reg        [7:0]    _zz_dataOut_payload_159_3;
  wire                _zz_dataOut_payload_160_32;
  wire       [7:0]    _zz_dataOut_payload_160_33;
  wire       [7:0]    _zz_dataOut_payload_176;
  wire                _zz_dataOut_payload_160_34;
  wire       [7:0]    _zz_dataOut_payload_160_35;
  wire       [7:0]    _zz_dataOut_payload_176_1;
  wire                _zz_dataOut_payload_160_36;
  wire       [7:0]    _zz_dataOut_payload_160_37;
  wire       [7:0]    _zz_dataOut_payload_176_2;
  wire                _zz_dataOut_payload_160_38;
  wire       [7:0]    _zz_dataOut_payload_160_39;
  wire       [7:0]    _zz_dataOut_payload_176_3;
  wire                _zz_dataOut_payload_160_40;
  wire       [7:0]    _zz_dataOut_payload_160_41;
  wire       [7:0]    _zz_dataOut_payload_176_4;
  wire                _zz_dataOut_payload_160_42;
  wire       [7:0]    _zz_dataOut_payload_160_43;
  wire       [7:0]    _zz_dataOut_payload_176_5;
  wire                _zz_dataOut_payload_160_44;
  wire       [7:0]    _zz_dataOut_payload_160_45;
  wire       [7:0]    _zz_dataOut_payload_176_6;
  wire                _zz_dataOut_payload_160_46;
  wire       [7:0]    _zz_dataOut_payload_160_47;
  wire       [7:0]    _zz_dataOut_payload_176_7;
  wire                _zz_dataOut_payload_160_48;
  wire       [7:0]    _zz_dataOut_payload_160_49;
  wire       [7:0]    _zz_dataOut_payload_176_8;
  wire                _zz_dataOut_payload_160_50;
  wire       [7:0]    _zz_dataOut_payload_160_51;
  wire       [7:0]    _zz_dataOut_payload_176_9;
  wire                _zz_dataOut_payload_160_52;
  wire       [7:0]    _zz_dataOut_payload_160_53;
  wire       [7:0]    _zz_dataOut_payload_176_10;
  wire                _zz_dataOut_payload_160_54;
  wire       [7:0]    _zz_dataOut_payload_160_55;
  wire       [7:0]    _zz_dataOut_payload_176_11;
  wire                _zz_dataOut_payload_160_56;
  wire       [7:0]    _zz_dataOut_payload_160_57;
  wire       [7:0]    _zz_dataOut_payload_176_12;
  wire                _zz_dataOut_payload_160_58;
  wire       [7:0]    _zz_dataOut_payload_160_59;
  wire       [7:0]    _zz_dataOut_payload_176_13;
  wire                _zz_dataOut_payload_160_60;
  wire       [7:0]    _zz_dataOut_payload_160_61;
  wire       [7:0]    _zz_dataOut_payload_176_14;
  wire                _zz_dataOut_payload_160_62;
  wire       [7:0]    _zz_dataOut_payload_160_63;
  wire       [7:0]    _zz_dataOut_payload_176_15;
  wire                _zz_dataOut_payload_160_64;
  wire       [7:0]    _zz_dataOut_payload_160_65;
  wire       [7:0]    _zz_dataOut_payload_168;
  wire                _zz_dataOut_payload_160_66;
  wire       [7:0]    _zz_dataOut_payload_160_67;
  wire       [7:0]    _zz_dataOut_payload_168_1;
  wire                _zz_dataOut_payload_160_68;
  wire       [7:0]    _zz_dataOut_payload_160_69;
  wire       [7:0]    _zz_dataOut_payload_168_2;
  wire                _zz_dataOut_payload_160_70;
  wire       [7:0]    _zz_dataOut_payload_160_71;
  wire       [7:0]    _zz_dataOut_payload_168_3;
  wire                _zz_dataOut_payload_160_72;
  wire       [7:0]    _zz_dataOut_payload_160_73;
  wire       [7:0]    _zz_dataOut_payload_168_4;
  wire                _zz_dataOut_payload_160_74;
  wire       [7:0]    _zz_dataOut_payload_160_75;
  wire       [7:0]    _zz_dataOut_payload_168_5;
  wire                _zz_dataOut_payload_160_76;
  wire       [7:0]    _zz_dataOut_payload_160_77;
  wire       [7:0]    _zz_dataOut_payload_168_6;
  wire                _zz_dataOut_payload_160_78;
  wire       [7:0]    _zz_dataOut_payload_160_79;
  wire       [7:0]    _zz_dataOut_payload_168_7;
  wire                _zz_dataOut_payload_160_80;
  wire       [7:0]    _zz_dataOut_payload_160_81;
  wire       [7:0]    _zz_dataOut_payload_164;
  wire                _zz_dataOut_payload_160_82;
  wire       [7:0]    _zz_dataOut_payload_160_83;
  wire       [7:0]    _zz_dataOut_payload_164_1;
  wire                _zz_dataOut_payload_160_84;
  wire       [7:0]    _zz_dataOut_payload_160_85;
  wire       [7:0]    _zz_dataOut_payload_164_2;
  wire                _zz_dataOut_payload_160_86;
  wire       [7:0]    _zz_dataOut_payload_160_87;
  wire       [7:0]    _zz_dataOut_payload_164_3;
  wire                _zz_dataOut_payload_160_88;
  wire       [7:0]    _zz_dataOut_payload_160_89;
  wire       [7:0]    _zz_dataOut_payload_162;
  wire                _zz_dataOut_payload_160_90;
  wire       [7:0]    _zz_dataOut_payload_160_91;
  wire       [7:0]    _zz_dataOut_payload_162_1;
  wire                _zz_dataOut_payload_160_92;
  wire                _zz_dataOut_payload_162_2;
  reg        [7:0]    _zz_dataOut_payload_160_93;
  reg        [7:0]    _zz_dataOut_payload_161;
  reg        [7:0]    _zz_dataOut_payload_162_3;
  reg        [7:0]    _zz_dataOut_payload_163;
  wire                _zz_dataOut_payload_164_4;
  wire       [7:0]    _zz_dataOut_payload_164_5;
  wire       [7:0]    _zz_dataOut_payload_166;
  wire                _zz_dataOut_payload_164_6;
  wire       [7:0]    _zz_dataOut_payload_164_7;
  wire       [7:0]    _zz_dataOut_payload_166_1;
  wire                _zz_dataOut_payload_164_8;
  wire                _zz_dataOut_payload_166_2;
  reg        [7:0]    _zz_dataOut_payload_164_9;
  reg        [7:0]    _zz_dataOut_payload_165;
  reg        [7:0]    _zz_dataOut_payload_166_3;
  reg        [7:0]    _zz_dataOut_payload_167;
  reg        [7:0]    _zz_dataOut_payload_160_94;
  reg        [7:0]    _zz_dataOut_payload_161_1;
  reg        [7:0]    _zz_dataOut_payload_162_4;
  reg        [7:0]    _zz_dataOut_payload_163_1;
  reg        [7:0]    _zz_dataOut_payload_164_10;
  reg        [7:0]    _zz_dataOut_payload_165_1;
  reg        [7:0]    _zz_dataOut_payload_166_4;
  reg        [7:0]    _zz_dataOut_payload_167_1;
  wire                _zz_dataOut_payload_168_8;
  wire       [7:0]    _zz_dataOut_payload_168_9;
  wire       [7:0]    _zz_dataOut_payload_172;
  wire                _zz_dataOut_payload_168_10;
  wire       [7:0]    _zz_dataOut_payload_168_11;
  wire       [7:0]    _zz_dataOut_payload_172_1;
  wire                _zz_dataOut_payload_168_12;
  wire       [7:0]    _zz_dataOut_payload_168_13;
  wire       [7:0]    _zz_dataOut_payload_172_2;
  wire                _zz_dataOut_payload_168_14;
  wire       [7:0]    _zz_dataOut_payload_168_15;
  wire       [7:0]    _zz_dataOut_payload_172_3;
  wire                _zz_dataOut_payload_168_16;
  wire       [7:0]    _zz_dataOut_payload_168_17;
  wire       [7:0]    _zz_dataOut_payload_170;
  wire                _zz_dataOut_payload_168_18;
  wire       [7:0]    _zz_dataOut_payload_168_19;
  wire       [7:0]    _zz_dataOut_payload_170_1;
  wire                _zz_dataOut_payload_168_20;
  wire                _zz_dataOut_payload_170_2;
  reg        [7:0]    _zz_dataOut_payload_168_21;
  reg        [7:0]    _zz_dataOut_payload_169;
  reg        [7:0]    _zz_dataOut_payload_170_3;
  reg        [7:0]    _zz_dataOut_payload_171;
  wire                _zz_dataOut_payload_172_4;
  wire       [7:0]    _zz_dataOut_payload_172_5;
  wire       [7:0]    _zz_dataOut_payload_174;
  wire                _zz_dataOut_payload_172_6;
  wire       [7:0]    _zz_dataOut_payload_172_7;
  wire       [7:0]    _zz_dataOut_payload_174_1;
  wire                _zz_dataOut_payload_172_8;
  wire                _zz_dataOut_payload_174_2;
  reg        [7:0]    _zz_dataOut_payload_172_9;
  reg        [7:0]    _zz_dataOut_payload_173;
  reg        [7:0]    _zz_dataOut_payload_174_3;
  reg        [7:0]    _zz_dataOut_payload_175;
  reg        [7:0]    _zz_dataOut_payload_168_22;
  reg        [7:0]    _zz_dataOut_payload_169_1;
  reg        [7:0]    _zz_dataOut_payload_170_4;
  reg        [7:0]    _zz_dataOut_payload_171_1;
  reg        [7:0]    _zz_dataOut_payload_172_10;
  reg        [7:0]    _zz_dataOut_payload_173_1;
  reg        [7:0]    _zz_dataOut_payload_174_4;
  reg        [7:0]    _zz_dataOut_payload_175_1;
  reg        [7:0]    _zz_dataOut_payload_160_95;
  reg        [7:0]    _zz_dataOut_payload_161_2;
  reg        [7:0]    _zz_dataOut_payload_162_5;
  reg        [7:0]    _zz_dataOut_payload_163_2;
  reg        [7:0]    _zz_dataOut_payload_164_11;
  reg        [7:0]    _zz_dataOut_payload_165_2;
  reg        [7:0]    _zz_dataOut_payload_166_5;
  reg        [7:0]    _zz_dataOut_payload_167_2;
  reg        [7:0]    _zz_dataOut_payload_168_23;
  reg        [7:0]    _zz_dataOut_payload_169_2;
  reg        [7:0]    _zz_dataOut_payload_170_5;
  reg        [7:0]    _zz_dataOut_payload_171_2;
  reg        [7:0]    _zz_dataOut_payload_172_11;
  reg        [7:0]    _zz_dataOut_payload_173_2;
  reg        [7:0]    _zz_dataOut_payload_174_5;
  reg        [7:0]    _zz_dataOut_payload_175_2;
  wire                _zz_dataOut_payload_176_16;
  wire       [7:0]    _zz_dataOut_payload_176_17;
  wire       [7:0]    _zz_dataOut_payload_184;
  wire                _zz_dataOut_payload_176_18;
  wire       [7:0]    _zz_dataOut_payload_176_19;
  wire       [7:0]    _zz_dataOut_payload_184_1;
  wire                _zz_dataOut_payload_176_20;
  wire       [7:0]    _zz_dataOut_payload_176_21;
  wire       [7:0]    _zz_dataOut_payload_184_2;
  wire                _zz_dataOut_payload_176_22;
  wire       [7:0]    _zz_dataOut_payload_176_23;
  wire       [7:0]    _zz_dataOut_payload_184_3;
  wire                _zz_dataOut_payload_176_24;
  wire       [7:0]    _zz_dataOut_payload_176_25;
  wire       [7:0]    _zz_dataOut_payload_184_4;
  wire                _zz_dataOut_payload_176_26;
  wire       [7:0]    _zz_dataOut_payload_176_27;
  wire       [7:0]    _zz_dataOut_payload_184_5;
  wire                _zz_dataOut_payload_176_28;
  wire       [7:0]    _zz_dataOut_payload_176_29;
  wire       [7:0]    _zz_dataOut_payload_184_6;
  wire                _zz_dataOut_payload_176_30;
  wire       [7:0]    _zz_dataOut_payload_176_31;
  wire       [7:0]    _zz_dataOut_payload_184_7;
  wire                _zz_dataOut_payload_176_32;
  wire       [7:0]    _zz_dataOut_payload_176_33;
  wire       [7:0]    _zz_dataOut_payload_180;
  wire                _zz_dataOut_payload_176_34;
  wire       [7:0]    _zz_dataOut_payload_176_35;
  wire       [7:0]    _zz_dataOut_payload_180_1;
  wire                _zz_dataOut_payload_176_36;
  wire       [7:0]    _zz_dataOut_payload_176_37;
  wire       [7:0]    _zz_dataOut_payload_180_2;
  wire                _zz_dataOut_payload_176_38;
  wire       [7:0]    _zz_dataOut_payload_176_39;
  wire       [7:0]    _zz_dataOut_payload_180_3;
  wire                _zz_dataOut_payload_176_40;
  wire       [7:0]    _zz_dataOut_payload_176_41;
  wire       [7:0]    _zz_dataOut_payload_178;
  wire                _zz_dataOut_payload_176_42;
  wire       [7:0]    _zz_dataOut_payload_176_43;
  wire       [7:0]    _zz_dataOut_payload_178_1;
  wire                _zz_dataOut_payload_176_44;
  wire                _zz_dataOut_payload_178_2;
  reg        [7:0]    _zz_dataOut_payload_176_45;
  reg        [7:0]    _zz_dataOut_payload_177;
  reg        [7:0]    _zz_dataOut_payload_178_3;
  reg        [7:0]    _zz_dataOut_payload_179;
  wire                _zz_dataOut_payload_180_4;
  wire       [7:0]    _zz_dataOut_payload_180_5;
  wire       [7:0]    _zz_dataOut_payload_182;
  wire                _zz_dataOut_payload_180_6;
  wire       [7:0]    _zz_dataOut_payload_180_7;
  wire       [7:0]    _zz_dataOut_payload_182_1;
  wire                _zz_dataOut_payload_180_8;
  wire                _zz_dataOut_payload_182_2;
  reg        [7:0]    _zz_dataOut_payload_180_9;
  reg        [7:0]    _zz_dataOut_payload_181;
  reg        [7:0]    _zz_dataOut_payload_182_3;
  reg        [7:0]    _zz_dataOut_payload_183;
  reg        [7:0]    _zz_dataOut_payload_176_46;
  reg        [7:0]    _zz_dataOut_payload_177_1;
  reg        [7:0]    _zz_dataOut_payload_178_4;
  reg        [7:0]    _zz_dataOut_payload_179_1;
  reg        [7:0]    _zz_dataOut_payload_180_10;
  reg        [7:0]    _zz_dataOut_payload_181_1;
  reg        [7:0]    _zz_dataOut_payload_182_4;
  reg        [7:0]    _zz_dataOut_payload_183_1;
  wire                _zz_dataOut_payload_184_8;
  wire       [7:0]    _zz_dataOut_payload_184_9;
  wire       [7:0]    _zz_dataOut_payload_188;
  wire                _zz_dataOut_payload_184_10;
  wire       [7:0]    _zz_dataOut_payload_184_11;
  wire       [7:0]    _zz_dataOut_payload_188_1;
  wire                _zz_dataOut_payload_184_12;
  wire       [7:0]    _zz_dataOut_payload_184_13;
  wire       [7:0]    _zz_dataOut_payload_188_2;
  wire                _zz_dataOut_payload_184_14;
  wire       [7:0]    _zz_dataOut_payload_184_15;
  wire       [7:0]    _zz_dataOut_payload_188_3;
  wire                _zz_dataOut_payload_184_16;
  wire       [7:0]    _zz_dataOut_payload_184_17;
  wire       [7:0]    _zz_dataOut_payload_186;
  wire                _zz_dataOut_payload_184_18;
  wire       [7:0]    _zz_dataOut_payload_184_19;
  wire       [7:0]    _zz_dataOut_payload_186_1;
  wire                _zz_dataOut_payload_184_20;
  wire                _zz_dataOut_payload_186_2;
  reg        [7:0]    _zz_dataOut_payload_184_21;
  reg        [7:0]    _zz_dataOut_payload_185;
  reg        [7:0]    _zz_dataOut_payload_186_3;
  reg        [7:0]    _zz_dataOut_payload_187;
  wire                _zz_dataOut_payload_188_4;
  wire       [7:0]    _zz_dataOut_payload_188_5;
  wire       [7:0]    _zz_dataOut_payload_190;
  wire                _zz_dataOut_payload_188_6;
  wire       [7:0]    _zz_dataOut_payload_188_7;
  wire       [7:0]    _zz_dataOut_payload_190_1;
  wire                _zz_dataOut_payload_188_8;
  wire                _zz_dataOut_payload_190_2;
  reg        [7:0]    _zz_dataOut_payload_188_9;
  reg        [7:0]    _zz_dataOut_payload_189;
  reg        [7:0]    _zz_dataOut_payload_190_3;
  reg        [7:0]    _zz_dataOut_payload_191;
  reg        [7:0]    _zz_dataOut_payload_184_22;
  reg        [7:0]    _zz_dataOut_payload_185_1;
  reg        [7:0]    _zz_dataOut_payload_186_4;
  reg        [7:0]    _zz_dataOut_payload_187_1;
  reg        [7:0]    _zz_dataOut_payload_188_10;
  reg        [7:0]    _zz_dataOut_payload_189_1;
  reg        [7:0]    _zz_dataOut_payload_190_4;
  reg        [7:0]    _zz_dataOut_payload_191_1;
  reg        [7:0]    _zz_dataOut_payload_176_47;
  reg        [7:0]    _zz_dataOut_payload_177_2;
  reg        [7:0]    _zz_dataOut_payload_178_5;
  reg        [7:0]    _zz_dataOut_payload_179_2;
  reg        [7:0]    _zz_dataOut_payload_180_11;
  reg        [7:0]    _zz_dataOut_payload_181_2;
  reg        [7:0]    _zz_dataOut_payload_182_5;
  reg        [7:0]    _zz_dataOut_payload_183_2;
  reg        [7:0]    _zz_dataOut_payload_184_23;
  reg        [7:0]    _zz_dataOut_payload_185_2;
  reg        [7:0]    _zz_dataOut_payload_186_5;
  reg        [7:0]    _zz_dataOut_payload_187_2;
  reg        [7:0]    _zz_dataOut_payload_188_11;
  reg        [7:0]    _zz_dataOut_payload_189_2;
  reg        [7:0]    _zz_dataOut_payload_190_5;
  reg        [7:0]    _zz_dataOut_payload_191_2;
  reg        [7:0]    _zz_dataOut_payload_160_96;
  reg        [7:0]    _zz_dataOut_payload_161_3;
  reg        [7:0]    _zz_dataOut_payload_162_6;
  reg        [7:0]    _zz_dataOut_payload_163_3;
  reg        [7:0]    _zz_dataOut_payload_164_12;
  reg        [7:0]    _zz_dataOut_payload_165_3;
  reg        [7:0]    _zz_dataOut_payload_166_6;
  reg        [7:0]    _zz_dataOut_payload_167_3;
  reg        [7:0]    _zz_dataOut_payload_168_24;
  reg        [7:0]    _zz_dataOut_payload_169_3;
  reg        [7:0]    _zz_dataOut_payload_170_6;
  reg        [7:0]    _zz_dataOut_payload_171_3;
  reg        [7:0]    _zz_dataOut_payload_172_12;
  reg        [7:0]    _zz_dataOut_payload_173_3;
  reg        [7:0]    _zz_dataOut_payload_174_6;
  reg        [7:0]    _zz_dataOut_payload_175_3;
  reg        [7:0]    _zz_dataOut_payload_176_48;
  reg        [7:0]    _zz_dataOut_payload_177_3;
  reg        [7:0]    _zz_dataOut_payload_178_6;
  reg        [7:0]    _zz_dataOut_payload_179_3;
  reg        [7:0]    _zz_dataOut_payload_180_12;
  reg        [7:0]    _zz_dataOut_payload_181_3;
  reg        [7:0]    _zz_dataOut_payload_182_6;
  reg        [7:0]    _zz_dataOut_payload_183_3;
  reg        [7:0]    _zz_dataOut_payload_184_24;
  reg        [7:0]    _zz_dataOut_payload_185_3;
  reg        [7:0]    _zz_dataOut_payload_186_6;
  reg        [7:0]    _zz_dataOut_payload_187_3;
  reg        [7:0]    _zz_dataOut_payload_188_12;
  reg        [7:0]    _zz_dataOut_payload_189_3;
  reg        [7:0]    _zz_dataOut_payload_190_6;
  reg        [7:0]    _zz_dataOut_payload_191_3;
  reg        [7:0]    _zz_dataOut_payload_128_385;
  reg        [7:0]    _zz_dataOut_payload_129_4;
  reg        [7:0]    _zz_dataOut_payload_130_7;
  reg        [7:0]    _zz_dataOut_payload_131_4;
  reg        [7:0]    _zz_dataOut_payload_132_13;
  reg        [7:0]    _zz_dataOut_payload_133_4;
  reg        [7:0]    _zz_dataOut_payload_134_7;
  reg        [7:0]    _zz_dataOut_payload_135_4;
  reg        [7:0]    _zz_dataOut_payload_136_25;
  reg        [7:0]    _zz_dataOut_payload_137_4;
  reg        [7:0]    _zz_dataOut_payload_138_7;
  reg        [7:0]    _zz_dataOut_payload_139_4;
  reg        [7:0]    _zz_dataOut_payload_140_13;
  reg        [7:0]    _zz_dataOut_payload_141_4;
  reg        [7:0]    _zz_dataOut_payload_142_7;
  reg        [7:0]    _zz_dataOut_payload_143_4;
  reg        [7:0]    _zz_dataOut_payload_144_49;
  reg        [7:0]    _zz_dataOut_payload_145_4;
  reg        [7:0]    _zz_dataOut_payload_146_7;
  reg        [7:0]    _zz_dataOut_payload_147_4;
  reg        [7:0]    _zz_dataOut_payload_148_13;
  reg        [7:0]    _zz_dataOut_payload_149_4;
  reg        [7:0]    _zz_dataOut_payload_150_7;
  reg        [7:0]    _zz_dataOut_payload_151_4;
  reg        [7:0]    _zz_dataOut_payload_152_25;
  reg        [7:0]    _zz_dataOut_payload_153_4;
  reg        [7:0]    _zz_dataOut_payload_154_7;
  reg        [7:0]    _zz_dataOut_payload_155_4;
  reg        [7:0]    _zz_dataOut_payload_156_13;
  reg        [7:0]    _zz_dataOut_payload_157_4;
  reg        [7:0]    _zz_dataOut_payload_158_7;
  reg        [7:0]    _zz_dataOut_payload_159_4;
  reg        [7:0]    _zz_dataOut_payload_160_97;
  reg        [7:0]    _zz_dataOut_payload_161_4;
  reg        [7:0]    _zz_dataOut_payload_162_7;
  reg        [7:0]    _zz_dataOut_payload_163_4;
  reg        [7:0]    _zz_dataOut_payload_164_13;
  reg        [7:0]    _zz_dataOut_payload_165_4;
  reg        [7:0]    _zz_dataOut_payload_166_7;
  reg        [7:0]    _zz_dataOut_payload_167_4;
  reg        [7:0]    _zz_dataOut_payload_168_25;
  reg        [7:0]    _zz_dataOut_payload_169_4;
  reg        [7:0]    _zz_dataOut_payload_170_7;
  reg        [7:0]    _zz_dataOut_payload_171_4;
  reg        [7:0]    _zz_dataOut_payload_172_13;
  reg        [7:0]    _zz_dataOut_payload_173_4;
  reg        [7:0]    _zz_dataOut_payload_174_7;
  reg        [7:0]    _zz_dataOut_payload_175_4;
  reg        [7:0]    _zz_dataOut_payload_176_49;
  reg        [7:0]    _zz_dataOut_payload_177_4;
  reg        [7:0]    _zz_dataOut_payload_178_7;
  reg        [7:0]    _zz_dataOut_payload_179_4;
  reg        [7:0]    _zz_dataOut_payload_180_13;
  reg        [7:0]    _zz_dataOut_payload_181_4;
  reg        [7:0]    _zz_dataOut_payload_182_7;
  reg        [7:0]    _zz_dataOut_payload_183_4;
  reg        [7:0]    _zz_dataOut_payload_184_25;
  reg        [7:0]    _zz_dataOut_payload_185_4;
  reg        [7:0]    _zz_dataOut_payload_186_7;
  reg        [7:0]    _zz_dataOut_payload_187_4;
  reg        [7:0]    _zz_dataOut_payload_188_13;
  reg        [7:0]    _zz_dataOut_payload_189_4;
  reg        [7:0]    _zz_dataOut_payload_190_7;
  reg        [7:0]    _zz_dataOut_payload_191_4;
  wire                _zz_dataOut_payload_192_64;
  wire       [7:0]    _zz_dataOut_payload_192_65;
  wire       [7:0]    _zz_dataOut_payload_224;
  wire                _zz_dataOut_payload_192_66;
  wire       [7:0]    _zz_dataOut_payload_192_67;
  wire       [7:0]    _zz_dataOut_payload_224_1;
  wire                _zz_dataOut_payload_192_68;
  wire       [7:0]    _zz_dataOut_payload_192_69;
  wire       [7:0]    _zz_dataOut_payload_224_2;
  wire                _zz_dataOut_payload_192_70;
  wire       [7:0]    _zz_dataOut_payload_192_71;
  wire       [7:0]    _zz_dataOut_payload_224_3;
  wire                _zz_dataOut_payload_192_72;
  wire       [7:0]    _zz_dataOut_payload_192_73;
  wire       [7:0]    _zz_dataOut_payload_224_4;
  wire                _zz_dataOut_payload_192_74;
  wire       [7:0]    _zz_dataOut_payload_192_75;
  wire       [7:0]    _zz_dataOut_payload_224_5;
  wire                _zz_dataOut_payload_192_76;
  wire       [7:0]    _zz_dataOut_payload_192_77;
  wire       [7:0]    _zz_dataOut_payload_224_6;
  wire                _zz_dataOut_payload_192_78;
  wire       [7:0]    _zz_dataOut_payload_192_79;
  wire       [7:0]    _zz_dataOut_payload_224_7;
  wire                _zz_dataOut_payload_192_80;
  wire       [7:0]    _zz_dataOut_payload_192_81;
  wire       [7:0]    _zz_dataOut_payload_224_8;
  wire                _zz_dataOut_payload_192_82;
  wire       [7:0]    _zz_dataOut_payload_192_83;
  wire       [7:0]    _zz_dataOut_payload_224_9;
  wire                _zz_dataOut_payload_192_84;
  wire       [7:0]    _zz_dataOut_payload_192_85;
  wire       [7:0]    _zz_dataOut_payload_224_10;
  wire                _zz_dataOut_payload_192_86;
  wire       [7:0]    _zz_dataOut_payload_192_87;
  wire       [7:0]    _zz_dataOut_payload_224_11;
  wire                _zz_dataOut_payload_192_88;
  wire       [7:0]    _zz_dataOut_payload_192_89;
  wire       [7:0]    _zz_dataOut_payload_224_12;
  wire                _zz_dataOut_payload_192_90;
  wire       [7:0]    _zz_dataOut_payload_192_91;
  wire       [7:0]    _zz_dataOut_payload_224_13;
  wire                _zz_dataOut_payload_192_92;
  wire       [7:0]    _zz_dataOut_payload_192_93;
  wire       [7:0]    _zz_dataOut_payload_224_14;
  wire                _zz_dataOut_payload_192_94;
  wire       [7:0]    _zz_dataOut_payload_192_95;
  wire       [7:0]    _zz_dataOut_payload_224_15;
  wire                _zz_dataOut_payload_192_96;
  wire       [7:0]    _zz_dataOut_payload_192_97;
  wire       [7:0]    _zz_dataOut_payload_224_16;
  wire                _zz_dataOut_payload_192_98;
  wire       [7:0]    _zz_dataOut_payload_192_99;
  wire       [7:0]    _zz_dataOut_payload_224_17;
  wire                _zz_dataOut_payload_192_100;
  wire       [7:0]    _zz_dataOut_payload_192_101;
  wire       [7:0]    _zz_dataOut_payload_224_18;
  wire                _zz_dataOut_payload_192_102;
  wire       [7:0]    _zz_dataOut_payload_192_103;
  wire       [7:0]    _zz_dataOut_payload_224_19;
  wire                _zz_dataOut_payload_192_104;
  wire       [7:0]    _zz_dataOut_payload_192_105;
  wire       [7:0]    _zz_dataOut_payload_224_20;
  wire                _zz_dataOut_payload_192_106;
  wire       [7:0]    _zz_dataOut_payload_192_107;
  wire       [7:0]    _zz_dataOut_payload_224_21;
  wire                _zz_dataOut_payload_192_108;
  wire       [7:0]    _zz_dataOut_payload_192_109;
  wire       [7:0]    _zz_dataOut_payload_224_22;
  wire                _zz_dataOut_payload_192_110;
  wire       [7:0]    _zz_dataOut_payload_192_111;
  wire       [7:0]    _zz_dataOut_payload_224_23;
  wire                _zz_dataOut_payload_192_112;
  wire       [7:0]    _zz_dataOut_payload_192_113;
  wire       [7:0]    _zz_dataOut_payload_224_24;
  wire                _zz_dataOut_payload_192_114;
  wire       [7:0]    _zz_dataOut_payload_192_115;
  wire       [7:0]    _zz_dataOut_payload_224_25;
  wire                _zz_dataOut_payload_192_116;
  wire       [7:0]    _zz_dataOut_payload_192_117;
  wire       [7:0]    _zz_dataOut_payload_224_26;
  wire                _zz_dataOut_payload_192_118;
  wire       [7:0]    _zz_dataOut_payload_192_119;
  wire       [7:0]    _zz_dataOut_payload_224_27;
  wire                _zz_dataOut_payload_192_120;
  wire       [7:0]    _zz_dataOut_payload_192_121;
  wire       [7:0]    _zz_dataOut_payload_224_28;
  wire                _zz_dataOut_payload_192_122;
  wire       [7:0]    _zz_dataOut_payload_192_123;
  wire       [7:0]    _zz_dataOut_payload_224_29;
  wire                _zz_dataOut_payload_192_124;
  wire       [7:0]    _zz_dataOut_payload_192_125;
  wire       [7:0]    _zz_dataOut_payload_224_30;
  wire                _zz_dataOut_payload_192_126;
  wire       [7:0]    _zz_dataOut_payload_192_127;
  wire       [7:0]    _zz_dataOut_payload_224_31;
  wire                _zz_dataOut_payload_192_128;
  wire       [7:0]    _zz_dataOut_payload_192_129;
  wire       [7:0]    _zz_dataOut_payload_208;
  wire                _zz_dataOut_payload_192_130;
  wire       [7:0]    _zz_dataOut_payload_192_131;
  wire       [7:0]    _zz_dataOut_payload_208_1;
  wire                _zz_dataOut_payload_192_132;
  wire       [7:0]    _zz_dataOut_payload_192_133;
  wire       [7:0]    _zz_dataOut_payload_208_2;
  wire                _zz_dataOut_payload_192_134;
  wire       [7:0]    _zz_dataOut_payload_192_135;
  wire       [7:0]    _zz_dataOut_payload_208_3;
  wire                _zz_dataOut_payload_192_136;
  wire       [7:0]    _zz_dataOut_payload_192_137;
  wire       [7:0]    _zz_dataOut_payload_208_4;
  wire                _zz_dataOut_payload_192_138;
  wire       [7:0]    _zz_dataOut_payload_192_139;
  wire       [7:0]    _zz_dataOut_payload_208_5;
  wire                _zz_dataOut_payload_192_140;
  wire       [7:0]    _zz_dataOut_payload_192_141;
  wire       [7:0]    _zz_dataOut_payload_208_6;
  wire                _zz_dataOut_payload_192_142;
  wire       [7:0]    _zz_dataOut_payload_192_143;
  wire       [7:0]    _zz_dataOut_payload_208_7;
  wire                _zz_dataOut_payload_192_144;
  wire       [7:0]    _zz_dataOut_payload_192_145;
  wire       [7:0]    _zz_dataOut_payload_208_8;
  wire                _zz_dataOut_payload_192_146;
  wire       [7:0]    _zz_dataOut_payload_192_147;
  wire       [7:0]    _zz_dataOut_payload_208_9;
  wire                _zz_dataOut_payload_192_148;
  wire       [7:0]    _zz_dataOut_payload_192_149;
  wire       [7:0]    _zz_dataOut_payload_208_10;
  wire                _zz_dataOut_payload_192_150;
  wire       [7:0]    _zz_dataOut_payload_192_151;
  wire       [7:0]    _zz_dataOut_payload_208_11;
  wire                _zz_dataOut_payload_192_152;
  wire       [7:0]    _zz_dataOut_payload_192_153;
  wire       [7:0]    _zz_dataOut_payload_208_12;
  wire                _zz_dataOut_payload_192_154;
  wire       [7:0]    _zz_dataOut_payload_192_155;
  wire       [7:0]    _zz_dataOut_payload_208_13;
  wire                _zz_dataOut_payload_192_156;
  wire       [7:0]    _zz_dataOut_payload_192_157;
  wire       [7:0]    _zz_dataOut_payload_208_14;
  wire                _zz_dataOut_payload_192_158;
  wire       [7:0]    _zz_dataOut_payload_192_159;
  wire       [7:0]    _zz_dataOut_payload_208_15;
  wire                _zz_dataOut_payload_192_160;
  wire       [7:0]    _zz_dataOut_payload_192_161;
  wire       [7:0]    _zz_dataOut_payload_200;
  wire                _zz_dataOut_payload_192_162;
  wire       [7:0]    _zz_dataOut_payload_192_163;
  wire       [7:0]    _zz_dataOut_payload_200_1;
  wire                _zz_dataOut_payload_192_164;
  wire       [7:0]    _zz_dataOut_payload_192_165;
  wire       [7:0]    _zz_dataOut_payload_200_2;
  wire                _zz_dataOut_payload_192_166;
  wire       [7:0]    _zz_dataOut_payload_192_167;
  wire       [7:0]    _zz_dataOut_payload_200_3;
  wire                _zz_dataOut_payload_192_168;
  wire       [7:0]    _zz_dataOut_payload_192_169;
  wire       [7:0]    _zz_dataOut_payload_200_4;
  wire                _zz_dataOut_payload_192_170;
  wire       [7:0]    _zz_dataOut_payload_192_171;
  wire       [7:0]    _zz_dataOut_payload_200_5;
  wire                _zz_dataOut_payload_192_172;
  wire       [7:0]    _zz_dataOut_payload_192_173;
  wire       [7:0]    _zz_dataOut_payload_200_6;
  wire                _zz_dataOut_payload_192_174;
  wire       [7:0]    _zz_dataOut_payload_192_175;
  wire       [7:0]    _zz_dataOut_payload_200_7;
  wire                _zz_dataOut_payload_192_176;
  wire       [7:0]    _zz_dataOut_payload_192_177;
  wire       [7:0]    _zz_dataOut_payload_196;
  wire                _zz_dataOut_payload_192_178;
  wire       [7:0]    _zz_dataOut_payload_192_179;
  wire       [7:0]    _zz_dataOut_payload_196_1;
  wire                _zz_dataOut_payload_192_180;
  wire       [7:0]    _zz_dataOut_payload_192_181;
  wire       [7:0]    _zz_dataOut_payload_196_2;
  wire                _zz_dataOut_payload_192_182;
  wire       [7:0]    _zz_dataOut_payload_192_183;
  wire       [7:0]    _zz_dataOut_payload_196_3;
  wire                _zz_dataOut_payload_192_184;
  wire       [7:0]    _zz_dataOut_payload_192_185;
  wire       [7:0]    _zz_dataOut_payload_194;
  wire                _zz_dataOut_payload_192_186;
  wire       [7:0]    _zz_dataOut_payload_192_187;
  wire       [7:0]    _zz_dataOut_payload_194_1;
  wire                _zz_dataOut_payload_192_188;
  wire                _zz_dataOut_payload_194_2;
  reg        [7:0]    _zz_dataOut_payload_192_189;
  reg        [7:0]    _zz_dataOut_payload_193;
  reg        [7:0]    _zz_dataOut_payload_194_3;
  reg        [7:0]    _zz_dataOut_payload_195;
  wire                _zz_dataOut_payload_196_4;
  wire       [7:0]    _zz_dataOut_payload_196_5;
  wire       [7:0]    _zz_dataOut_payload_198;
  wire                _zz_dataOut_payload_196_6;
  wire       [7:0]    _zz_dataOut_payload_196_7;
  wire       [7:0]    _zz_dataOut_payload_198_1;
  wire                _zz_dataOut_payload_196_8;
  wire                _zz_dataOut_payload_198_2;
  reg        [7:0]    _zz_dataOut_payload_196_9;
  reg        [7:0]    _zz_dataOut_payload_197;
  reg        [7:0]    _zz_dataOut_payload_198_3;
  reg        [7:0]    _zz_dataOut_payload_199;
  reg        [7:0]    _zz_dataOut_payload_192_190;
  reg        [7:0]    _zz_dataOut_payload_193_1;
  reg        [7:0]    _zz_dataOut_payload_194_4;
  reg        [7:0]    _zz_dataOut_payload_195_1;
  reg        [7:0]    _zz_dataOut_payload_196_10;
  reg        [7:0]    _zz_dataOut_payload_197_1;
  reg        [7:0]    _zz_dataOut_payload_198_4;
  reg        [7:0]    _zz_dataOut_payload_199_1;
  wire                _zz_dataOut_payload_200_8;
  wire       [7:0]    _zz_dataOut_payload_200_9;
  wire       [7:0]    _zz_dataOut_payload_204;
  wire                _zz_dataOut_payload_200_10;
  wire       [7:0]    _zz_dataOut_payload_200_11;
  wire       [7:0]    _zz_dataOut_payload_204_1;
  wire                _zz_dataOut_payload_200_12;
  wire       [7:0]    _zz_dataOut_payload_200_13;
  wire       [7:0]    _zz_dataOut_payload_204_2;
  wire                _zz_dataOut_payload_200_14;
  wire       [7:0]    _zz_dataOut_payload_200_15;
  wire       [7:0]    _zz_dataOut_payload_204_3;
  wire                _zz_dataOut_payload_200_16;
  wire       [7:0]    _zz_dataOut_payload_200_17;
  wire       [7:0]    _zz_dataOut_payload_202;
  wire                _zz_dataOut_payload_200_18;
  wire       [7:0]    _zz_dataOut_payload_200_19;
  wire       [7:0]    _zz_dataOut_payload_202_1;
  wire                _zz_dataOut_payload_200_20;
  wire                _zz_dataOut_payload_202_2;
  reg        [7:0]    _zz_dataOut_payload_200_21;
  reg        [7:0]    _zz_dataOut_payload_201;
  reg        [7:0]    _zz_dataOut_payload_202_3;
  reg        [7:0]    _zz_dataOut_payload_203;
  wire                _zz_dataOut_payload_204_4;
  wire       [7:0]    _zz_dataOut_payload_204_5;
  wire       [7:0]    _zz_dataOut_payload_206;
  wire                _zz_dataOut_payload_204_6;
  wire       [7:0]    _zz_dataOut_payload_204_7;
  wire       [7:0]    _zz_dataOut_payload_206_1;
  wire                _zz_dataOut_payload_204_8;
  wire                _zz_dataOut_payload_206_2;
  reg        [7:0]    _zz_dataOut_payload_204_9;
  reg        [7:0]    _zz_dataOut_payload_205;
  reg        [7:0]    _zz_dataOut_payload_206_3;
  reg        [7:0]    _zz_dataOut_payload_207;
  reg        [7:0]    _zz_dataOut_payload_200_22;
  reg        [7:0]    _zz_dataOut_payload_201_1;
  reg        [7:0]    _zz_dataOut_payload_202_4;
  reg        [7:0]    _zz_dataOut_payload_203_1;
  reg        [7:0]    _zz_dataOut_payload_204_10;
  reg        [7:0]    _zz_dataOut_payload_205_1;
  reg        [7:0]    _zz_dataOut_payload_206_4;
  reg        [7:0]    _zz_dataOut_payload_207_1;
  reg        [7:0]    _zz_dataOut_payload_192_191;
  reg        [7:0]    _zz_dataOut_payload_193_2;
  reg        [7:0]    _zz_dataOut_payload_194_5;
  reg        [7:0]    _zz_dataOut_payload_195_2;
  reg        [7:0]    _zz_dataOut_payload_196_11;
  reg        [7:0]    _zz_dataOut_payload_197_2;
  reg        [7:0]    _zz_dataOut_payload_198_5;
  reg        [7:0]    _zz_dataOut_payload_199_2;
  reg        [7:0]    _zz_dataOut_payload_200_23;
  reg        [7:0]    _zz_dataOut_payload_201_2;
  reg        [7:0]    _zz_dataOut_payload_202_5;
  reg        [7:0]    _zz_dataOut_payload_203_2;
  reg        [7:0]    _zz_dataOut_payload_204_11;
  reg        [7:0]    _zz_dataOut_payload_205_2;
  reg        [7:0]    _zz_dataOut_payload_206_5;
  reg        [7:0]    _zz_dataOut_payload_207_2;
  wire                _zz_dataOut_payload_208_16;
  wire       [7:0]    _zz_dataOut_payload_208_17;
  wire       [7:0]    _zz_dataOut_payload_216;
  wire                _zz_dataOut_payload_208_18;
  wire       [7:0]    _zz_dataOut_payload_208_19;
  wire       [7:0]    _zz_dataOut_payload_216_1;
  wire                _zz_dataOut_payload_208_20;
  wire       [7:0]    _zz_dataOut_payload_208_21;
  wire       [7:0]    _zz_dataOut_payload_216_2;
  wire                _zz_dataOut_payload_208_22;
  wire       [7:0]    _zz_dataOut_payload_208_23;
  wire       [7:0]    _zz_dataOut_payload_216_3;
  wire                _zz_dataOut_payload_208_24;
  wire       [7:0]    _zz_dataOut_payload_208_25;
  wire       [7:0]    _zz_dataOut_payload_216_4;
  wire                _zz_dataOut_payload_208_26;
  wire       [7:0]    _zz_dataOut_payload_208_27;
  wire       [7:0]    _zz_dataOut_payload_216_5;
  wire                _zz_dataOut_payload_208_28;
  wire       [7:0]    _zz_dataOut_payload_208_29;
  wire       [7:0]    _zz_dataOut_payload_216_6;
  wire                _zz_dataOut_payload_208_30;
  wire       [7:0]    _zz_dataOut_payload_208_31;
  wire       [7:0]    _zz_dataOut_payload_216_7;
  wire                _zz_dataOut_payload_208_32;
  wire       [7:0]    _zz_dataOut_payload_208_33;
  wire       [7:0]    _zz_dataOut_payload_212;
  wire                _zz_dataOut_payload_208_34;
  wire       [7:0]    _zz_dataOut_payload_208_35;
  wire       [7:0]    _zz_dataOut_payload_212_1;
  wire                _zz_dataOut_payload_208_36;
  wire       [7:0]    _zz_dataOut_payload_208_37;
  wire       [7:0]    _zz_dataOut_payload_212_2;
  wire                _zz_dataOut_payload_208_38;
  wire       [7:0]    _zz_dataOut_payload_208_39;
  wire       [7:0]    _zz_dataOut_payload_212_3;
  wire                _zz_dataOut_payload_208_40;
  wire       [7:0]    _zz_dataOut_payload_208_41;
  wire       [7:0]    _zz_dataOut_payload_210;
  wire                _zz_dataOut_payload_208_42;
  wire       [7:0]    _zz_dataOut_payload_208_43;
  wire       [7:0]    _zz_dataOut_payload_210_1;
  wire                _zz_dataOut_payload_208_44;
  wire                _zz_dataOut_payload_210_2;
  reg        [7:0]    _zz_dataOut_payload_208_45;
  reg        [7:0]    _zz_dataOut_payload_209;
  reg        [7:0]    _zz_dataOut_payload_210_3;
  reg        [7:0]    _zz_dataOut_payload_211;
  wire                _zz_dataOut_payload_212_4;
  wire       [7:0]    _zz_dataOut_payload_212_5;
  wire       [7:0]    _zz_dataOut_payload_214;
  wire                _zz_dataOut_payload_212_6;
  wire       [7:0]    _zz_dataOut_payload_212_7;
  wire       [7:0]    _zz_dataOut_payload_214_1;
  wire                _zz_dataOut_payload_212_8;
  wire                _zz_dataOut_payload_214_2;
  reg        [7:0]    _zz_dataOut_payload_212_9;
  reg        [7:0]    _zz_dataOut_payload_213;
  reg        [7:0]    _zz_dataOut_payload_214_3;
  reg        [7:0]    _zz_dataOut_payload_215;
  reg        [7:0]    _zz_dataOut_payload_208_46;
  reg        [7:0]    _zz_dataOut_payload_209_1;
  reg        [7:0]    _zz_dataOut_payload_210_4;
  reg        [7:0]    _zz_dataOut_payload_211_1;
  reg        [7:0]    _zz_dataOut_payload_212_10;
  reg        [7:0]    _zz_dataOut_payload_213_1;
  reg        [7:0]    _zz_dataOut_payload_214_4;
  reg        [7:0]    _zz_dataOut_payload_215_1;
  wire                _zz_dataOut_payload_216_8;
  wire       [7:0]    _zz_dataOut_payload_216_9;
  wire       [7:0]    _zz_dataOut_payload_220;
  wire                _zz_dataOut_payload_216_10;
  wire       [7:0]    _zz_dataOut_payload_216_11;
  wire       [7:0]    _zz_dataOut_payload_220_1;
  wire                _zz_dataOut_payload_216_12;
  wire       [7:0]    _zz_dataOut_payload_216_13;
  wire       [7:0]    _zz_dataOut_payload_220_2;
  wire                _zz_dataOut_payload_216_14;
  wire       [7:0]    _zz_dataOut_payload_216_15;
  wire       [7:0]    _zz_dataOut_payload_220_3;
  wire                _zz_dataOut_payload_216_16;
  wire       [7:0]    _zz_dataOut_payload_216_17;
  wire       [7:0]    _zz_dataOut_payload_218;
  wire                _zz_dataOut_payload_216_18;
  wire       [7:0]    _zz_dataOut_payload_216_19;
  wire       [7:0]    _zz_dataOut_payload_218_1;
  wire                _zz_dataOut_payload_216_20;
  wire                _zz_dataOut_payload_218_2;
  reg        [7:0]    _zz_dataOut_payload_216_21;
  reg        [7:0]    _zz_dataOut_payload_217;
  reg        [7:0]    _zz_dataOut_payload_218_3;
  reg        [7:0]    _zz_dataOut_payload_219;
  wire                _zz_dataOut_payload_220_4;
  wire       [7:0]    _zz_dataOut_payload_220_5;
  wire       [7:0]    _zz_dataOut_payload_222;
  wire                _zz_dataOut_payload_220_6;
  wire       [7:0]    _zz_dataOut_payload_220_7;
  wire       [7:0]    _zz_dataOut_payload_222_1;
  wire                _zz_dataOut_payload_220_8;
  wire                _zz_dataOut_payload_222_2;
  reg        [7:0]    _zz_dataOut_payload_220_9;
  reg        [7:0]    _zz_dataOut_payload_221;
  reg        [7:0]    _zz_dataOut_payload_222_3;
  reg        [7:0]    _zz_dataOut_payload_223;
  reg        [7:0]    _zz_dataOut_payload_216_22;
  reg        [7:0]    _zz_dataOut_payload_217_1;
  reg        [7:0]    _zz_dataOut_payload_218_4;
  reg        [7:0]    _zz_dataOut_payload_219_1;
  reg        [7:0]    _zz_dataOut_payload_220_10;
  reg        [7:0]    _zz_dataOut_payload_221_1;
  reg        [7:0]    _zz_dataOut_payload_222_4;
  reg        [7:0]    _zz_dataOut_payload_223_1;
  reg        [7:0]    _zz_dataOut_payload_208_47;
  reg        [7:0]    _zz_dataOut_payload_209_2;
  reg        [7:0]    _zz_dataOut_payload_210_5;
  reg        [7:0]    _zz_dataOut_payload_211_2;
  reg        [7:0]    _zz_dataOut_payload_212_11;
  reg        [7:0]    _zz_dataOut_payload_213_2;
  reg        [7:0]    _zz_dataOut_payload_214_5;
  reg        [7:0]    _zz_dataOut_payload_215_2;
  reg        [7:0]    _zz_dataOut_payload_216_23;
  reg        [7:0]    _zz_dataOut_payload_217_2;
  reg        [7:0]    _zz_dataOut_payload_218_5;
  reg        [7:0]    _zz_dataOut_payload_219_2;
  reg        [7:0]    _zz_dataOut_payload_220_11;
  reg        [7:0]    _zz_dataOut_payload_221_2;
  reg        [7:0]    _zz_dataOut_payload_222_5;
  reg        [7:0]    _zz_dataOut_payload_223_2;
  reg        [7:0]    _zz_dataOut_payload_192_192;
  reg        [7:0]    _zz_dataOut_payload_193_3;
  reg        [7:0]    _zz_dataOut_payload_194_6;
  reg        [7:0]    _zz_dataOut_payload_195_3;
  reg        [7:0]    _zz_dataOut_payload_196_12;
  reg        [7:0]    _zz_dataOut_payload_197_3;
  reg        [7:0]    _zz_dataOut_payload_198_6;
  reg        [7:0]    _zz_dataOut_payload_199_3;
  reg        [7:0]    _zz_dataOut_payload_200_24;
  reg        [7:0]    _zz_dataOut_payload_201_3;
  reg        [7:0]    _zz_dataOut_payload_202_6;
  reg        [7:0]    _zz_dataOut_payload_203_3;
  reg        [7:0]    _zz_dataOut_payload_204_12;
  reg        [7:0]    _zz_dataOut_payload_205_3;
  reg        [7:0]    _zz_dataOut_payload_206_6;
  reg        [7:0]    _zz_dataOut_payload_207_3;
  reg        [7:0]    _zz_dataOut_payload_208_48;
  reg        [7:0]    _zz_dataOut_payload_209_3;
  reg        [7:0]    _zz_dataOut_payload_210_6;
  reg        [7:0]    _zz_dataOut_payload_211_3;
  reg        [7:0]    _zz_dataOut_payload_212_12;
  reg        [7:0]    _zz_dataOut_payload_213_3;
  reg        [7:0]    _zz_dataOut_payload_214_6;
  reg        [7:0]    _zz_dataOut_payload_215_3;
  reg        [7:0]    _zz_dataOut_payload_216_24;
  reg        [7:0]    _zz_dataOut_payload_217_3;
  reg        [7:0]    _zz_dataOut_payload_218_6;
  reg        [7:0]    _zz_dataOut_payload_219_3;
  reg        [7:0]    _zz_dataOut_payload_220_12;
  reg        [7:0]    _zz_dataOut_payload_221_3;
  reg        [7:0]    _zz_dataOut_payload_222_6;
  reg        [7:0]    _zz_dataOut_payload_223_3;
  wire                _zz_dataOut_payload_224_32;
  wire       [7:0]    _zz_dataOut_payload_224_33;
  wire       [7:0]    _zz_dataOut_payload_240;
  wire                _zz_dataOut_payload_224_34;
  wire       [7:0]    _zz_dataOut_payload_224_35;
  wire       [7:0]    _zz_dataOut_payload_240_1;
  wire                _zz_dataOut_payload_224_36;
  wire       [7:0]    _zz_dataOut_payload_224_37;
  wire       [7:0]    _zz_dataOut_payload_240_2;
  wire                _zz_dataOut_payload_224_38;
  wire       [7:0]    _zz_dataOut_payload_224_39;
  wire       [7:0]    _zz_dataOut_payload_240_3;
  wire                _zz_dataOut_payload_224_40;
  wire       [7:0]    _zz_dataOut_payload_224_41;
  wire       [7:0]    _zz_dataOut_payload_240_4;
  wire                _zz_dataOut_payload_224_42;
  wire       [7:0]    _zz_dataOut_payload_224_43;
  wire       [7:0]    _zz_dataOut_payload_240_5;
  wire                _zz_dataOut_payload_224_44;
  wire       [7:0]    _zz_dataOut_payload_224_45;
  wire       [7:0]    _zz_dataOut_payload_240_6;
  wire                _zz_dataOut_payload_224_46;
  wire       [7:0]    _zz_dataOut_payload_224_47;
  wire       [7:0]    _zz_dataOut_payload_240_7;
  wire                _zz_dataOut_payload_224_48;
  wire       [7:0]    _zz_dataOut_payload_224_49;
  wire       [7:0]    _zz_dataOut_payload_240_8;
  wire                _zz_dataOut_payload_224_50;
  wire       [7:0]    _zz_dataOut_payload_224_51;
  wire       [7:0]    _zz_dataOut_payload_240_9;
  wire                _zz_dataOut_payload_224_52;
  wire       [7:0]    _zz_dataOut_payload_224_53;
  wire       [7:0]    _zz_dataOut_payload_240_10;
  wire                _zz_dataOut_payload_224_54;
  wire       [7:0]    _zz_dataOut_payload_224_55;
  wire       [7:0]    _zz_dataOut_payload_240_11;
  wire                _zz_dataOut_payload_224_56;
  wire       [7:0]    _zz_dataOut_payload_224_57;
  wire       [7:0]    _zz_dataOut_payload_240_12;
  wire                _zz_dataOut_payload_224_58;
  wire       [7:0]    _zz_dataOut_payload_224_59;
  wire       [7:0]    _zz_dataOut_payload_240_13;
  wire                _zz_dataOut_payload_224_60;
  wire       [7:0]    _zz_dataOut_payload_224_61;
  wire       [7:0]    _zz_dataOut_payload_240_14;
  wire                _zz_dataOut_payload_224_62;
  wire       [7:0]    _zz_dataOut_payload_224_63;
  wire       [7:0]    _zz_dataOut_payload_240_15;
  wire                _zz_dataOut_payload_224_64;
  wire       [7:0]    _zz_dataOut_payload_224_65;
  wire       [7:0]    _zz_dataOut_payload_232;
  wire                _zz_dataOut_payload_224_66;
  wire       [7:0]    _zz_dataOut_payload_224_67;
  wire       [7:0]    _zz_dataOut_payload_232_1;
  wire                _zz_dataOut_payload_224_68;
  wire       [7:0]    _zz_dataOut_payload_224_69;
  wire       [7:0]    _zz_dataOut_payload_232_2;
  wire                _zz_dataOut_payload_224_70;
  wire       [7:0]    _zz_dataOut_payload_224_71;
  wire       [7:0]    _zz_dataOut_payload_232_3;
  wire                _zz_dataOut_payload_224_72;
  wire       [7:0]    _zz_dataOut_payload_224_73;
  wire       [7:0]    _zz_dataOut_payload_232_4;
  wire                _zz_dataOut_payload_224_74;
  wire       [7:0]    _zz_dataOut_payload_224_75;
  wire       [7:0]    _zz_dataOut_payload_232_5;
  wire                _zz_dataOut_payload_224_76;
  wire       [7:0]    _zz_dataOut_payload_224_77;
  wire       [7:0]    _zz_dataOut_payload_232_6;
  wire                _zz_dataOut_payload_224_78;
  wire       [7:0]    _zz_dataOut_payload_224_79;
  wire       [7:0]    _zz_dataOut_payload_232_7;
  wire                _zz_dataOut_payload_224_80;
  wire       [7:0]    _zz_dataOut_payload_224_81;
  wire       [7:0]    _zz_dataOut_payload_228;
  wire                _zz_dataOut_payload_224_82;
  wire       [7:0]    _zz_dataOut_payload_224_83;
  wire       [7:0]    _zz_dataOut_payload_228_1;
  wire                _zz_dataOut_payload_224_84;
  wire       [7:0]    _zz_dataOut_payload_224_85;
  wire       [7:0]    _zz_dataOut_payload_228_2;
  wire                _zz_dataOut_payload_224_86;
  wire       [7:0]    _zz_dataOut_payload_224_87;
  wire       [7:0]    _zz_dataOut_payload_228_3;
  wire                _zz_dataOut_payload_224_88;
  wire       [7:0]    _zz_dataOut_payload_224_89;
  wire       [7:0]    _zz_dataOut_payload_226;
  wire                _zz_dataOut_payload_224_90;
  wire       [7:0]    _zz_dataOut_payload_224_91;
  wire       [7:0]    _zz_dataOut_payload_226_1;
  wire                _zz_dataOut_payload_224_92;
  wire                _zz_dataOut_payload_226_2;
  reg        [7:0]    _zz_dataOut_payload_224_93;
  reg        [7:0]    _zz_dataOut_payload_225;
  reg        [7:0]    _zz_dataOut_payload_226_3;
  reg        [7:0]    _zz_dataOut_payload_227;
  wire                _zz_dataOut_payload_228_4;
  wire       [7:0]    _zz_dataOut_payload_228_5;
  wire       [7:0]    _zz_dataOut_payload_230;
  wire                _zz_dataOut_payload_228_6;
  wire       [7:0]    _zz_dataOut_payload_228_7;
  wire       [7:0]    _zz_dataOut_payload_230_1;
  wire                _zz_dataOut_payload_228_8;
  wire                _zz_dataOut_payload_230_2;
  reg        [7:0]    _zz_dataOut_payload_228_9;
  reg        [7:0]    _zz_dataOut_payload_229;
  reg        [7:0]    _zz_dataOut_payload_230_3;
  reg        [7:0]    _zz_dataOut_payload_231;
  reg        [7:0]    _zz_dataOut_payload_224_94;
  reg        [7:0]    _zz_dataOut_payload_225_1;
  reg        [7:0]    _zz_dataOut_payload_226_4;
  reg        [7:0]    _zz_dataOut_payload_227_1;
  reg        [7:0]    _zz_dataOut_payload_228_10;
  reg        [7:0]    _zz_dataOut_payload_229_1;
  reg        [7:0]    _zz_dataOut_payload_230_4;
  reg        [7:0]    _zz_dataOut_payload_231_1;
  wire                _zz_dataOut_payload_232_8;
  wire       [7:0]    _zz_dataOut_payload_232_9;
  wire       [7:0]    _zz_dataOut_payload_236;
  wire                _zz_dataOut_payload_232_10;
  wire       [7:0]    _zz_dataOut_payload_232_11;
  wire       [7:0]    _zz_dataOut_payload_236_1;
  wire                _zz_dataOut_payload_232_12;
  wire       [7:0]    _zz_dataOut_payload_232_13;
  wire       [7:0]    _zz_dataOut_payload_236_2;
  wire                _zz_dataOut_payload_232_14;
  wire       [7:0]    _zz_dataOut_payload_232_15;
  wire       [7:0]    _zz_dataOut_payload_236_3;
  wire                _zz_dataOut_payload_232_16;
  wire       [7:0]    _zz_dataOut_payload_232_17;
  wire       [7:0]    _zz_dataOut_payload_234;
  wire                _zz_dataOut_payload_232_18;
  wire       [7:0]    _zz_dataOut_payload_232_19;
  wire       [7:0]    _zz_dataOut_payload_234_1;
  wire                _zz_dataOut_payload_232_20;
  wire                _zz_dataOut_payload_234_2;
  reg        [7:0]    _zz_dataOut_payload_232_21;
  reg        [7:0]    _zz_dataOut_payload_233;
  reg        [7:0]    _zz_dataOut_payload_234_3;
  reg        [7:0]    _zz_dataOut_payload_235;
  wire                _zz_dataOut_payload_236_4;
  wire       [7:0]    _zz_dataOut_payload_236_5;
  wire       [7:0]    _zz_dataOut_payload_238;
  wire                _zz_dataOut_payload_236_6;
  wire       [7:0]    _zz_dataOut_payload_236_7;
  wire       [7:0]    _zz_dataOut_payload_238_1;
  wire                _zz_dataOut_payload_236_8;
  wire                _zz_dataOut_payload_238_2;
  reg        [7:0]    _zz_dataOut_payload_236_9;
  reg        [7:0]    _zz_dataOut_payload_237;
  reg        [7:0]    _zz_dataOut_payload_238_3;
  reg        [7:0]    _zz_dataOut_payload_239;
  reg        [7:0]    _zz_dataOut_payload_232_22;
  reg        [7:0]    _zz_dataOut_payload_233_1;
  reg        [7:0]    _zz_dataOut_payload_234_4;
  reg        [7:0]    _zz_dataOut_payload_235_1;
  reg        [7:0]    _zz_dataOut_payload_236_10;
  reg        [7:0]    _zz_dataOut_payload_237_1;
  reg        [7:0]    _zz_dataOut_payload_238_4;
  reg        [7:0]    _zz_dataOut_payload_239_1;
  reg        [7:0]    _zz_dataOut_payload_224_95;
  reg        [7:0]    _zz_dataOut_payload_225_2;
  reg        [7:0]    _zz_dataOut_payload_226_5;
  reg        [7:0]    _zz_dataOut_payload_227_2;
  reg        [7:0]    _zz_dataOut_payload_228_11;
  reg        [7:0]    _zz_dataOut_payload_229_2;
  reg        [7:0]    _zz_dataOut_payload_230_5;
  reg        [7:0]    _zz_dataOut_payload_231_2;
  reg        [7:0]    _zz_dataOut_payload_232_23;
  reg        [7:0]    _zz_dataOut_payload_233_2;
  reg        [7:0]    _zz_dataOut_payload_234_5;
  reg        [7:0]    _zz_dataOut_payload_235_2;
  reg        [7:0]    _zz_dataOut_payload_236_11;
  reg        [7:0]    _zz_dataOut_payload_237_2;
  reg        [7:0]    _zz_dataOut_payload_238_5;
  reg        [7:0]    _zz_dataOut_payload_239_2;
  wire                _zz_dataOut_payload_240_16;
  wire       [7:0]    _zz_dataOut_payload_240_17;
  wire       [7:0]    _zz_dataOut_payload_248;
  wire                _zz_dataOut_payload_240_18;
  wire       [7:0]    _zz_dataOut_payload_240_19;
  wire       [7:0]    _zz_dataOut_payload_248_1;
  wire                _zz_dataOut_payload_240_20;
  wire       [7:0]    _zz_dataOut_payload_240_21;
  wire       [7:0]    _zz_dataOut_payload_248_2;
  wire                _zz_dataOut_payload_240_22;
  wire       [7:0]    _zz_dataOut_payload_240_23;
  wire       [7:0]    _zz_dataOut_payload_248_3;
  wire                _zz_dataOut_payload_240_24;
  wire       [7:0]    _zz_dataOut_payload_240_25;
  wire       [7:0]    _zz_dataOut_payload_248_4;
  wire                _zz_dataOut_payload_240_26;
  wire       [7:0]    _zz_dataOut_payload_240_27;
  wire       [7:0]    _zz_dataOut_payload_248_5;
  wire                _zz_dataOut_payload_240_28;
  wire       [7:0]    _zz_dataOut_payload_240_29;
  wire       [7:0]    _zz_dataOut_payload_248_6;
  wire                _zz_dataOut_payload_240_30;
  wire       [7:0]    _zz_dataOut_payload_240_31;
  wire       [7:0]    _zz_dataOut_payload_248_7;
  wire                _zz_dataOut_payload_240_32;
  wire       [7:0]    _zz_dataOut_payload_240_33;
  wire       [7:0]    _zz_dataOut_payload_244;
  wire                _zz_dataOut_payload_240_34;
  wire       [7:0]    _zz_dataOut_payload_240_35;
  wire       [7:0]    _zz_dataOut_payload_244_1;
  wire                _zz_dataOut_payload_240_36;
  wire       [7:0]    _zz_dataOut_payload_240_37;
  wire       [7:0]    _zz_dataOut_payload_244_2;
  wire                _zz_dataOut_payload_240_38;
  wire       [7:0]    _zz_dataOut_payload_240_39;
  wire       [7:0]    _zz_dataOut_payload_244_3;
  wire                _zz_dataOut_payload_240_40;
  wire       [7:0]    _zz_dataOut_payload_240_41;
  wire       [7:0]    _zz_dataOut_payload_242;
  wire                _zz_dataOut_payload_240_42;
  wire       [7:0]    _zz_dataOut_payload_240_43;
  wire       [7:0]    _zz_dataOut_payload_242_1;
  wire                _zz_dataOut_payload_240_44;
  wire                _zz_dataOut_payload_242_2;
  reg        [7:0]    _zz_dataOut_payload_240_45;
  reg        [7:0]    _zz_dataOut_payload_241;
  reg        [7:0]    _zz_dataOut_payload_242_3;
  reg        [7:0]    _zz_dataOut_payload_243;
  wire                _zz_dataOut_payload_244_4;
  wire       [7:0]    _zz_dataOut_payload_244_5;
  wire       [7:0]    _zz_dataOut_payload_246;
  wire                _zz_dataOut_payload_244_6;
  wire       [7:0]    _zz_dataOut_payload_244_7;
  wire       [7:0]    _zz_dataOut_payload_246_1;
  wire                _zz_dataOut_payload_244_8;
  wire                _zz_dataOut_payload_246_2;
  reg        [7:0]    _zz_dataOut_payload_244_9;
  reg        [7:0]    _zz_dataOut_payload_245;
  reg        [7:0]    _zz_dataOut_payload_246_3;
  reg        [7:0]    _zz_dataOut_payload_247;
  reg        [7:0]    _zz_dataOut_payload_240_46;
  reg        [7:0]    _zz_dataOut_payload_241_1;
  reg        [7:0]    _zz_dataOut_payload_242_4;
  reg        [7:0]    _zz_dataOut_payload_243_1;
  reg        [7:0]    _zz_dataOut_payload_244_10;
  reg        [7:0]    _zz_dataOut_payload_245_1;
  reg        [7:0]    _zz_dataOut_payload_246_4;
  reg        [7:0]    _zz_dataOut_payload_247_1;
  wire                _zz_dataOut_payload_248_8;
  wire       [7:0]    _zz_dataOut_payload_248_9;
  wire       [7:0]    _zz_dataOut_payload_252;
  wire                _zz_dataOut_payload_248_10;
  wire       [7:0]    _zz_dataOut_payload_248_11;
  wire       [7:0]    _zz_dataOut_payload_252_1;
  wire                _zz_dataOut_payload_248_12;
  wire       [7:0]    _zz_dataOut_payload_248_13;
  wire       [7:0]    _zz_dataOut_payload_252_2;
  wire                _zz_dataOut_payload_248_14;
  wire       [7:0]    _zz_dataOut_payload_248_15;
  wire       [7:0]    _zz_dataOut_payload_252_3;
  wire                _zz_dataOut_payload_248_16;
  wire       [7:0]    _zz_dataOut_payload_248_17;
  wire       [7:0]    _zz_dataOut_payload_250;
  wire                _zz_dataOut_payload_248_18;
  wire       [7:0]    _zz_dataOut_payload_248_19;
  wire       [7:0]    _zz_dataOut_payload_250_1;
  wire                _zz_dataOut_payload_248_20;
  wire                _zz_dataOut_payload_250_2;
  reg        [7:0]    _zz_dataOut_payload_248_21;
  reg        [7:0]    _zz_dataOut_payload_249;
  reg        [7:0]    _zz_dataOut_payload_250_3;
  reg        [7:0]    _zz_dataOut_payload_251;
  wire                _zz_dataOut_payload_252_4;
  wire       [7:0]    _zz_dataOut_payload_252_5;
  wire       [7:0]    _zz_dataOut_payload_254;
  wire                _zz_dataOut_payload_252_6;
  wire       [7:0]    _zz_dataOut_payload_252_7;
  wire       [7:0]    _zz_dataOut_payload_254_1;
  wire                _zz_dataOut_payload_252_8;
  wire                _zz_dataOut_payload_254_2;
  reg        [7:0]    _zz_dataOut_payload_252_9;
  reg        [7:0]    _zz_dataOut_payload_253;
  reg        [7:0]    _zz_dataOut_payload_254_3;
  reg        [7:0]    _zz_dataOut_payload_255;
  reg        [7:0]    _zz_dataOut_payload_248_22;
  reg        [7:0]    _zz_dataOut_payload_249_1;
  reg        [7:0]    _zz_dataOut_payload_250_4;
  reg        [7:0]    _zz_dataOut_payload_251_1;
  reg        [7:0]    _zz_dataOut_payload_252_10;
  reg        [7:0]    _zz_dataOut_payload_253_1;
  reg        [7:0]    _zz_dataOut_payload_254_4;
  reg        [7:0]    _zz_dataOut_payload_255_1;
  reg        [7:0]    _zz_dataOut_payload_240_47;
  reg        [7:0]    _zz_dataOut_payload_241_2;
  reg        [7:0]    _zz_dataOut_payload_242_5;
  reg        [7:0]    _zz_dataOut_payload_243_2;
  reg        [7:0]    _zz_dataOut_payload_244_11;
  reg        [7:0]    _zz_dataOut_payload_245_2;
  reg        [7:0]    _zz_dataOut_payload_246_5;
  reg        [7:0]    _zz_dataOut_payload_247_2;
  reg        [7:0]    _zz_dataOut_payload_248_23;
  reg        [7:0]    _zz_dataOut_payload_249_2;
  reg        [7:0]    _zz_dataOut_payload_250_5;
  reg        [7:0]    _zz_dataOut_payload_251_2;
  reg        [7:0]    _zz_dataOut_payload_252_11;
  reg        [7:0]    _zz_dataOut_payload_253_2;
  reg        [7:0]    _zz_dataOut_payload_254_5;
  reg        [7:0]    _zz_dataOut_payload_255_2;
  reg        [7:0]    _zz_dataOut_payload_224_96;
  reg        [7:0]    _zz_dataOut_payload_225_3;
  reg        [7:0]    _zz_dataOut_payload_226_6;
  reg        [7:0]    _zz_dataOut_payload_227_3;
  reg        [7:0]    _zz_dataOut_payload_228_12;
  reg        [7:0]    _zz_dataOut_payload_229_3;
  reg        [7:0]    _zz_dataOut_payload_230_6;
  reg        [7:0]    _zz_dataOut_payload_231_3;
  reg        [7:0]    _zz_dataOut_payload_232_24;
  reg        [7:0]    _zz_dataOut_payload_233_3;
  reg        [7:0]    _zz_dataOut_payload_234_6;
  reg        [7:0]    _zz_dataOut_payload_235_3;
  reg        [7:0]    _zz_dataOut_payload_236_12;
  reg        [7:0]    _zz_dataOut_payload_237_3;
  reg        [7:0]    _zz_dataOut_payload_238_6;
  reg        [7:0]    _zz_dataOut_payload_239_3;
  reg        [7:0]    _zz_dataOut_payload_240_48;
  reg        [7:0]    _zz_dataOut_payload_241_3;
  reg        [7:0]    _zz_dataOut_payload_242_6;
  reg        [7:0]    _zz_dataOut_payload_243_3;
  reg        [7:0]    _zz_dataOut_payload_244_12;
  reg        [7:0]    _zz_dataOut_payload_245_3;
  reg        [7:0]    _zz_dataOut_payload_246_6;
  reg        [7:0]    _zz_dataOut_payload_247_3;
  reg        [7:0]    _zz_dataOut_payload_248_24;
  reg        [7:0]    _zz_dataOut_payload_249_3;
  reg        [7:0]    _zz_dataOut_payload_250_6;
  reg        [7:0]    _zz_dataOut_payload_251_3;
  reg        [7:0]    _zz_dataOut_payload_252_12;
  reg        [7:0]    _zz_dataOut_payload_253_3;
  reg        [7:0]    _zz_dataOut_payload_254_6;
  reg        [7:0]    _zz_dataOut_payload_255_3;
  reg        [7:0]    _zz_dataOut_payload_192_193;
  reg        [7:0]    _zz_dataOut_payload_193_4;
  reg        [7:0]    _zz_dataOut_payload_194_7;
  reg        [7:0]    _zz_dataOut_payload_195_4;
  reg        [7:0]    _zz_dataOut_payload_196_13;
  reg        [7:0]    _zz_dataOut_payload_197_4;
  reg        [7:0]    _zz_dataOut_payload_198_7;
  reg        [7:0]    _zz_dataOut_payload_199_4;
  reg        [7:0]    _zz_dataOut_payload_200_25;
  reg        [7:0]    _zz_dataOut_payload_201_4;
  reg        [7:0]    _zz_dataOut_payload_202_7;
  reg        [7:0]    _zz_dataOut_payload_203_4;
  reg        [7:0]    _zz_dataOut_payload_204_13;
  reg        [7:0]    _zz_dataOut_payload_205_4;
  reg        [7:0]    _zz_dataOut_payload_206_7;
  reg        [7:0]    _zz_dataOut_payload_207_4;
  reg        [7:0]    _zz_dataOut_payload_208_49;
  reg        [7:0]    _zz_dataOut_payload_209_4;
  reg        [7:0]    _zz_dataOut_payload_210_7;
  reg        [7:0]    _zz_dataOut_payload_211_4;
  reg        [7:0]    _zz_dataOut_payload_212_13;
  reg        [7:0]    _zz_dataOut_payload_213_4;
  reg        [7:0]    _zz_dataOut_payload_214_7;
  reg        [7:0]    _zz_dataOut_payload_215_4;
  reg        [7:0]    _zz_dataOut_payload_216_25;
  reg        [7:0]    _zz_dataOut_payload_217_4;
  reg        [7:0]    _zz_dataOut_payload_218_7;
  reg        [7:0]    _zz_dataOut_payload_219_4;
  reg        [7:0]    _zz_dataOut_payload_220_13;
  reg        [7:0]    _zz_dataOut_payload_221_4;
  reg        [7:0]    _zz_dataOut_payload_222_7;
  reg        [7:0]    _zz_dataOut_payload_223_4;
  reg        [7:0]    _zz_dataOut_payload_224_97;
  reg        [7:0]    _zz_dataOut_payload_225_4;
  reg        [7:0]    _zz_dataOut_payload_226_7;
  reg        [7:0]    _zz_dataOut_payload_227_4;
  reg        [7:0]    _zz_dataOut_payload_228_13;
  reg        [7:0]    _zz_dataOut_payload_229_4;
  reg        [7:0]    _zz_dataOut_payload_230_7;
  reg        [7:0]    _zz_dataOut_payload_231_4;
  reg        [7:0]    _zz_dataOut_payload_232_25;
  reg        [7:0]    _zz_dataOut_payload_233_4;
  reg        [7:0]    _zz_dataOut_payload_234_7;
  reg        [7:0]    _zz_dataOut_payload_235_4;
  reg        [7:0]    _zz_dataOut_payload_236_13;
  reg        [7:0]    _zz_dataOut_payload_237_4;
  reg        [7:0]    _zz_dataOut_payload_238_7;
  reg        [7:0]    _zz_dataOut_payload_239_4;
  reg        [7:0]    _zz_dataOut_payload_240_49;
  reg        [7:0]    _zz_dataOut_payload_241_4;
  reg        [7:0]    _zz_dataOut_payload_242_7;
  reg        [7:0]    _zz_dataOut_payload_243_4;
  reg        [7:0]    _zz_dataOut_payload_244_13;
  reg        [7:0]    _zz_dataOut_payload_245_4;
  reg        [7:0]    _zz_dataOut_payload_246_7;
  reg        [7:0]    _zz_dataOut_payload_247_4;
  reg        [7:0]    _zz_dataOut_payload_248_25;
  reg        [7:0]    _zz_dataOut_payload_249_4;
  reg        [7:0]    _zz_dataOut_payload_250_7;
  reg        [7:0]    _zz_dataOut_payload_251_4;
  reg        [7:0]    _zz_dataOut_payload_252_13;
  reg        [7:0]    _zz_dataOut_payload_253_4;
  reg        [7:0]    _zz_dataOut_payload_254_7;
  reg        [7:0]    _zz_dataOut_payload_255_4;
  reg        [7:0]    _zz_dataOut_payload_128_386;
  reg        [7:0]    _zz_dataOut_payload_129_5;
  reg        [7:0]    _zz_dataOut_payload_130_8;
  reg        [7:0]    _zz_dataOut_payload_131_5;
  reg        [7:0]    _zz_dataOut_payload_132_14;
  reg        [7:0]    _zz_dataOut_payload_133_5;
  reg        [7:0]    _zz_dataOut_payload_134_8;
  reg        [7:0]    _zz_dataOut_payload_135_5;
  reg        [7:0]    _zz_dataOut_payload_136_26;
  reg        [7:0]    _zz_dataOut_payload_137_5;
  reg        [7:0]    _zz_dataOut_payload_138_8;
  reg        [7:0]    _zz_dataOut_payload_139_5;
  reg        [7:0]    _zz_dataOut_payload_140_14;
  reg        [7:0]    _zz_dataOut_payload_141_5;
  reg        [7:0]    _zz_dataOut_payload_142_8;
  reg        [7:0]    _zz_dataOut_payload_143_5;
  reg        [7:0]    _zz_dataOut_payload_144_50;
  reg        [7:0]    _zz_dataOut_payload_145_5;
  reg        [7:0]    _zz_dataOut_payload_146_8;
  reg        [7:0]    _zz_dataOut_payload_147_5;
  reg        [7:0]    _zz_dataOut_payload_148_14;
  reg        [7:0]    _zz_dataOut_payload_149_5;
  reg        [7:0]    _zz_dataOut_payload_150_8;
  reg        [7:0]    _zz_dataOut_payload_151_5;
  reg        [7:0]    _zz_dataOut_payload_152_26;
  reg        [7:0]    _zz_dataOut_payload_153_5;
  reg        [7:0]    _zz_dataOut_payload_154_8;
  reg        [7:0]    _zz_dataOut_payload_155_5;
  reg        [7:0]    _zz_dataOut_payload_156_14;
  reg        [7:0]    _zz_dataOut_payload_157_5;
  reg        [7:0]    _zz_dataOut_payload_158_8;
  reg        [7:0]    _zz_dataOut_payload_159_5;
  reg        [7:0]    _zz_dataOut_payload_160_98;
  reg        [7:0]    _zz_dataOut_payload_161_5;
  reg        [7:0]    _zz_dataOut_payload_162_8;
  reg        [7:0]    _zz_dataOut_payload_163_5;
  reg        [7:0]    _zz_dataOut_payload_164_14;
  reg        [7:0]    _zz_dataOut_payload_165_5;
  reg        [7:0]    _zz_dataOut_payload_166_8;
  reg        [7:0]    _zz_dataOut_payload_167_5;
  reg        [7:0]    _zz_dataOut_payload_168_26;
  reg        [7:0]    _zz_dataOut_payload_169_5;
  reg        [7:0]    _zz_dataOut_payload_170_8;
  reg        [7:0]    _zz_dataOut_payload_171_5;
  reg        [7:0]    _zz_dataOut_payload_172_14;
  reg        [7:0]    _zz_dataOut_payload_173_5;
  reg        [7:0]    _zz_dataOut_payload_174_8;
  reg        [7:0]    _zz_dataOut_payload_175_5;
  reg        [7:0]    _zz_dataOut_payload_176_50;
  reg        [7:0]    _zz_dataOut_payload_177_5;
  reg        [7:0]    _zz_dataOut_payload_178_8;
  reg        [7:0]    _zz_dataOut_payload_179_5;
  reg        [7:0]    _zz_dataOut_payload_180_14;
  reg        [7:0]    _zz_dataOut_payload_181_5;
  reg        [7:0]    _zz_dataOut_payload_182_8;
  reg        [7:0]    _zz_dataOut_payload_183_5;
  reg        [7:0]    _zz_dataOut_payload_184_26;
  reg        [7:0]    _zz_dataOut_payload_185_5;
  reg        [7:0]    _zz_dataOut_payload_186_8;
  reg        [7:0]    _zz_dataOut_payload_187_5;
  reg        [7:0]    _zz_dataOut_payload_188_14;
  reg        [7:0]    _zz_dataOut_payload_189_5;
  reg        [7:0]    _zz_dataOut_payload_190_8;
  reg        [7:0]    _zz_dataOut_payload_191_5;
  reg        [7:0]    _zz_dataOut_payload_192_194;
  reg        [7:0]    _zz_dataOut_payload_193_5;
  reg        [7:0]    _zz_dataOut_payload_194_8;
  reg        [7:0]    _zz_dataOut_payload_195_5;
  reg        [7:0]    _zz_dataOut_payload_196_14;
  reg        [7:0]    _zz_dataOut_payload_197_5;
  reg        [7:0]    _zz_dataOut_payload_198_8;
  reg        [7:0]    _zz_dataOut_payload_199_5;
  reg        [7:0]    _zz_dataOut_payload_200_26;
  reg        [7:0]    _zz_dataOut_payload_201_5;
  reg        [7:0]    _zz_dataOut_payload_202_8;
  reg        [7:0]    _zz_dataOut_payload_203_5;
  reg        [7:0]    _zz_dataOut_payload_204_14;
  reg        [7:0]    _zz_dataOut_payload_205_5;
  reg        [7:0]    _zz_dataOut_payload_206_8;
  reg        [7:0]    _zz_dataOut_payload_207_5;
  reg        [7:0]    _zz_dataOut_payload_208_50;
  reg        [7:0]    _zz_dataOut_payload_209_5;
  reg        [7:0]    _zz_dataOut_payload_210_8;
  reg        [7:0]    _zz_dataOut_payload_211_5;
  reg        [7:0]    _zz_dataOut_payload_212_14;
  reg        [7:0]    _zz_dataOut_payload_213_5;
  reg        [7:0]    _zz_dataOut_payload_214_8;
  reg        [7:0]    _zz_dataOut_payload_215_5;
  reg        [7:0]    _zz_dataOut_payload_216_26;
  reg        [7:0]    _zz_dataOut_payload_217_5;
  reg        [7:0]    _zz_dataOut_payload_218_8;
  reg        [7:0]    _zz_dataOut_payload_219_5;
  reg        [7:0]    _zz_dataOut_payload_220_14;
  reg        [7:0]    _zz_dataOut_payload_221_5;
  reg        [7:0]    _zz_dataOut_payload_222_8;
  reg        [7:0]    _zz_dataOut_payload_223_5;
  reg        [7:0]    _zz_dataOut_payload_224_98;
  reg        [7:0]    _zz_dataOut_payload_225_5;
  reg        [7:0]    _zz_dataOut_payload_226_8;
  reg        [7:0]    _zz_dataOut_payload_227_5;
  reg        [7:0]    _zz_dataOut_payload_228_14;
  reg        [7:0]    _zz_dataOut_payload_229_5;
  reg        [7:0]    _zz_dataOut_payload_230_8;
  reg        [7:0]    _zz_dataOut_payload_231_5;
  reg        [7:0]    _zz_dataOut_payload_232_26;
  reg        [7:0]    _zz_dataOut_payload_233_5;
  reg        [7:0]    _zz_dataOut_payload_234_8;
  reg        [7:0]    _zz_dataOut_payload_235_5;
  reg        [7:0]    _zz_dataOut_payload_236_14;
  reg        [7:0]    _zz_dataOut_payload_237_5;
  reg        [7:0]    _zz_dataOut_payload_238_8;
  reg        [7:0]    _zz_dataOut_payload_239_5;
  reg        [7:0]    _zz_dataOut_payload_240_50;
  reg        [7:0]    _zz_dataOut_payload_241_5;
  reg        [7:0]    _zz_dataOut_payload_242_8;
  reg        [7:0]    _zz_dataOut_payload_243_5;
  reg        [7:0]    _zz_dataOut_payload_244_14;
  reg        [7:0]    _zz_dataOut_payload_245_5;
  reg        [7:0]    _zz_dataOut_payload_246_8;
  reg        [7:0]    _zz_dataOut_payload_247_5;
  reg        [7:0]    _zz_dataOut_payload_248_26;
  reg        [7:0]    _zz_dataOut_payload_249_5;
  reg        [7:0]    _zz_dataOut_payload_250_8;
  reg        [7:0]    _zz_dataOut_payload_251_5;
  reg        [7:0]    _zz_dataOut_payload_252_14;
  reg        [7:0]    _zz_dataOut_payload_253_5;
  reg        [7:0]    _zz_dataOut_payload_254_8;
  reg        [7:0]    _zz_dataOut_payload_255_5;
  reg        [7:0]    _zz_dataOut_payload_0_16643;
  reg        [7:0]    _zz_dataOut_payload_1_6;
  reg        [7:0]    _zz_dataOut_payload_2_9;
  reg        [7:0]    _zz_dataOut_payload_3_6;
  reg        [7:0]    _zz_dataOut_payload_4_15;
  reg        [7:0]    _zz_dataOut_payload_5_6;
  reg        [7:0]    _zz_dataOut_payload_6_9;
  reg        [7:0]    _zz_dataOut_payload_7_6;
  reg        [7:0]    _zz_dataOut_payload_8_27;
  reg        [7:0]    _zz_dataOut_payload_9_6;
  reg        [7:0]    _zz_dataOut_payload_10_9;
  reg        [7:0]    _zz_dataOut_payload_11_6;
  reg        [7:0]    _zz_dataOut_payload_12_15;
  reg        [7:0]    _zz_dataOut_payload_13_6;
  reg        [7:0]    _zz_dataOut_payload_14_9;
  reg        [7:0]    _zz_dataOut_payload_15_6;
  reg        [7:0]    _zz_dataOut_payload_16_51;
  reg        [7:0]    _zz_dataOut_payload_17_6;
  reg        [7:0]    _zz_dataOut_payload_18_9;
  reg        [7:0]    _zz_dataOut_payload_19_6;
  reg        [7:0]    _zz_dataOut_payload_20_15;
  reg        [7:0]    _zz_dataOut_payload_21_6;
  reg        [7:0]    _zz_dataOut_payload_22_9;
  reg        [7:0]    _zz_dataOut_payload_23_6;
  reg        [7:0]    _zz_dataOut_payload_24_27;
  reg        [7:0]    _zz_dataOut_payload_25_6;
  reg        [7:0]    _zz_dataOut_payload_26_9;
  reg        [7:0]    _zz_dataOut_payload_27_6;
  reg        [7:0]    _zz_dataOut_payload_28_15;
  reg        [7:0]    _zz_dataOut_payload_29_6;
  reg        [7:0]    _zz_dataOut_payload_30_9;
  reg        [7:0]    _zz_dataOut_payload_31_6;
  reg        [7:0]    _zz_dataOut_payload_32_99;
  reg        [7:0]    _zz_dataOut_payload_33_6;
  reg        [7:0]    _zz_dataOut_payload_34_9;
  reg        [7:0]    _zz_dataOut_payload_35_6;
  reg        [7:0]    _zz_dataOut_payload_36_15;
  reg        [7:0]    _zz_dataOut_payload_37_6;
  reg        [7:0]    _zz_dataOut_payload_38_9;
  reg        [7:0]    _zz_dataOut_payload_39_6;
  reg        [7:0]    _zz_dataOut_payload_40_27;
  reg        [7:0]    _zz_dataOut_payload_41_6;
  reg        [7:0]    _zz_dataOut_payload_42_9;
  reg        [7:0]    _zz_dataOut_payload_43_6;
  reg        [7:0]    _zz_dataOut_payload_44_15;
  reg        [7:0]    _zz_dataOut_payload_45_6;
  reg        [7:0]    _zz_dataOut_payload_46_9;
  reg        [7:0]    _zz_dataOut_payload_47_6;
  reg        [7:0]    _zz_dataOut_payload_48_51;
  reg        [7:0]    _zz_dataOut_payload_49_6;
  reg        [7:0]    _zz_dataOut_payload_50_9;
  reg        [7:0]    _zz_dataOut_payload_51_6;
  reg        [7:0]    _zz_dataOut_payload_52_15;
  reg        [7:0]    _zz_dataOut_payload_53_6;
  reg        [7:0]    _zz_dataOut_payload_54_9;
  reg        [7:0]    _zz_dataOut_payload_55_6;
  reg        [7:0]    _zz_dataOut_payload_56_27;
  reg        [7:0]    _zz_dataOut_payload_57_6;
  reg        [7:0]    _zz_dataOut_payload_58_9;
  reg        [7:0]    _zz_dataOut_payload_59_6;
  reg        [7:0]    _zz_dataOut_payload_60_15;
  reg        [7:0]    _zz_dataOut_payload_61_6;
  reg        [7:0]    _zz_dataOut_payload_62_9;
  reg        [7:0]    _zz_dataOut_payload_63_6;
  reg        [7:0]    _zz_dataOut_payload_64_195;
  reg        [7:0]    _zz_dataOut_payload_65_6;
  reg        [7:0]    _zz_dataOut_payload_66_9;
  reg        [7:0]    _zz_dataOut_payload_67_6;
  reg        [7:0]    _zz_dataOut_payload_68_15;
  reg        [7:0]    _zz_dataOut_payload_69_6;
  reg        [7:0]    _zz_dataOut_payload_70_9;
  reg        [7:0]    _zz_dataOut_payload_71_6;
  reg        [7:0]    _zz_dataOut_payload_72_27;
  reg        [7:0]    _zz_dataOut_payload_73_6;
  reg        [7:0]    _zz_dataOut_payload_74_9;
  reg        [7:0]    _zz_dataOut_payload_75_6;
  reg        [7:0]    _zz_dataOut_payload_76_15;
  reg        [7:0]    _zz_dataOut_payload_77_6;
  reg        [7:0]    _zz_dataOut_payload_78_9;
  reg        [7:0]    _zz_dataOut_payload_79_6;
  reg        [7:0]    _zz_dataOut_payload_80_51;
  reg        [7:0]    _zz_dataOut_payload_81_6;
  reg        [7:0]    _zz_dataOut_payload_82_9;
  reg        [7:0]    _zz_dataOut_payload_83_6;
  reg        [7:0]    _zz_dataOut_payload_84_15;
  reg        [7:0]    _zz_dataOut_payload_85_6;
  reg        [7:0]    _zz_dataOut_payload_86_9;
  reg        [7:0]    _zz_dataOut_payload_87_6;
  reg        [7:0]    _zz_dataOut_payload_88_27;
  reg        [7:0]    _zz_dataOut_payload_89_6;
  reg        [7:0]    _zz_dataOut_payload_90_9;
  reg        [7:0]    _zz_dataOut_payload_91_6;
  reg        [7:0]    _zz_dataOut_payload_92_15;
  reg        [7:0]    _zz_dataOut_payload_93_6;
  reg        [7:0]    _zz_dataOut_payload_94_9;
  reg        [7:0]    _zz_dataOut_payload_95_6;
  reg        [7:0]    _zz_dataOut_payload_96_99;
  reg        [7:0]    _zz_dataOut_payload_97_6;
  reg        [7:0]    _zz_dataOut_payload_98_9;
  reg        [7:0]    _zz_dataOut_payload_99_6;
  reg        [7:0]    _zz_dataOut_payload_100_15;
  reg        [7:0]    _zz_dataOut_payload_101_6;
  reg        [7:0]    _zz_dataOut_payload_102_9;
  reg        [7:0]    _zz_dataOut_payload_103_6;
  reg        [7:0]    _zz_dataOut_payload_104_27;
  reg        [7:0]    _zz_dataOut_payload_105_6;
  reg        [7:0]    _zz_dataOut_payload_106_9;
  reg        [7:0]    _zz_dataOut_payload_107_6;
  reg        [7:0]    _zz_dataOut_payload_108_15;
  reg        [7:0]    _zz_dataOut_payload_109_6;
  reg        [7:0]    _zz_dataOut_payload_110_9;
  reg        [7:0]    _zz_dataOut_payload_111_6;
  reg        [7:0]    _zz_dataOut_payload_112_51;
  reg        [7:0]    _zz_dataOut_payload_113_6;
  reg        [7:0]    _zz_dataOut_payload_114_9;
  reg        [7:0]    _zz_dataOut_payload_115_6;
  reg        [7:0]    _zz_dataOut_payload_116_15;
  reg        [7:0]    _zz_dataOut_payload_117_6;
  reg        [7:0]    _zz_dataOut_payload_118_9;
  reg        [7:0]    _zz_dataOut_payload_119_6;
  reg        [7:0]    _zz_dataOut_payload_120_27;
  reg        [7:0]    _zz_dataOut_payload_121_6;
  reg        [7:0]    _zz_dataOut_payload_122_9;
  reg        [7:0]    _zz_dataOut_payload_123_6;
  reg        [7:0]    _zz_dataOut_payload_124_15;
  reg        [7:0]    _zz_dataOut_payload_125_6;
  reg        [7:0]    _zz_dataOut_payload_126_9;
  reg        [7:0]    _zz_dataOut_payload_127_6;
  reg        [7:0]    _zz_dataOut_payload_128_387;
  reg        [7:0]    _zz_dataOut_payload_129_6;
  reg        [7:0]    _zz_dataOut_payload_130_9;
  reg        [7:0]    _zz_dataOut_payload_131_6;
  reg        [7:0]    _zz_dataOut_payload_132_15;
  reg        [7:0]    _zz_dataOut_payload_133_6;
  reg        [7:0]    _zz_dataOut_payload_134_9;
  reg        [7:0]    _zz_dataOut_payload_135_6;
  reg        [7:0]    _zz_dataOut_payload_136_27;
  reg        [7:0]    _zz_dataOut_payload_137_6;
  reg        [7:0]    _zz_dataOut_payload_138_9;
  reg        [7:0]    _zz_dataOut_payload_139_6;
  reg        [7:0]    _zz_dataOut_payload_140_15;
  reg        [7:0]    _zz_dataOut_payload_141_6;
  reg        [7:0]    _zz_dataOut_payload_142_9;
  reg        [7:0]    _zz_dataOut_payload_143_6;
  reg        [7:0]    _zz_dataOut_payload_144_51;
  reg        [7:0]    _zz_dataOut_payload_145_6;
  reg        [7:0]    _zz_dataOut_payload_146_9;
  reg        [7:0]    _zz_dataOut_payload_147_6;
  reg        [7:0]    _zz_dataOut_payload_148_15;
  reg        [7:0]    _zz_dataOut_payload_149_6;
  reg        [7:0]    _zz_dataOut_payload_150_9;
  reg        [7:0]    _zz_dataOut_payload_151_6;
  reg        [7:0]    _zz_dataOut_payload_152_27;
  reg        [7:0]    _zz_dataOut_payload_153_6;
  reg        [7:0]    _zz_dataOut_payload_154_9;
  reg        [7:0]    _zz_dataOut_payload_155_6;
  reg        [7:0]    _zz_dataOut_payload_156_15;
  reg        [7:0]    _zz_dataOut_payload_157_6;
  reg        [7:0]    _zz_dataOut_payload_158_9;
  reg        [7:0]    _zz_dataOut_payload_159_6;
  reg        [7:0]    _zz_dataOut_payload_160_99;
  reg        [7:0]    _zz_dataOut_payload_161_6;
  reg        [7:0]    _zz_dataOut_payload_162_9;
  reg        [7:0]    _zz_dataOut_payload_163_6;
  reg        [7:0]    _zz_dataOut_payload_164_15;
  reg        [7:0]    _zz_dataOut_payload_165_6;
  reg        [7:0]    _zz_dataOut_payload_166_9;
  reg        [7:0]    _zz_dataOut_payload_167_6;
  reg        [7:0]    _zz_dataOut_payload_168_27;
  reg        [7:0]    _zz_dataOut_payload_169_6;
  reg        [7:0]    _zz_dataOut_payload_170_9;
  reg        [7:0]    _zz_dataOut_payload_171_6;
  reg        [7:0]    _zz_dataOut_payload_172_15;
  reg        [7:0]    _zz_dataOut_payload_173_6;
  reg        [7:0]    _zz_dataOut_payload_174_9;
  reg        [7:0]    _zz_dataOut_payload_175_6;
  reg        [7:0]    _zz_dataOut_payload_176_51;
  reg        [7:0]    _zz_dataOut_payload_177_6;
  reg        [7:0]    _zz_dataOut_payload_178_9;
  reg        [7:0]    _zz_dataOut_payload_179_6;
  reg        [7:0]    _zz_dataOut_payload_180_15;
  reg        [7:0]    _zz_dataOut_payload_181_6;
  reg        [7:0]    _zz_dataOut_payload_182_9;
  reg        [7:0]    _zz_dataOut_payload_183_6;
  reg        [7:0]    _zz_dataOut_payload_184_27;
  reg        [7:0]    _zz_dataOut_payload_185_6;
  reg        [7:0]    _zz_dataOut_payload_186_9;
  reg        [7:0]    _zz_dataOut_payload_187_6;
  reg        [7:0]    _zz_dataOut_payload_188_15;
  reg        [7:0]    _zz_dataOut_payload_189_6;
  reg        [7:0]    _zz_dataOut_payload_190_9;
  reg        [7:0]    _zz_dataOut_payload_191_6;
  reg        [7:0]    _zz_dataOut_payload_192_195;
  reg        [7:0]    _zz_dataOut_payload_193_6;
  reg        [7:0]    _zz_dataOut_payload_194_9;
  reg        [7:0]    _zz_dataOut_payload_195_6;
  reg        [7:0]    _zz_dataOut_payload_196_15;
  reg        [7:0]    _zz_dataOut_payload_197_6;
  reg        [7:0]    _zz_dataOut_payload_198_9;
  reg        [7:0]    _zz_dataOut_payload_199_6;
  reg        [7:0]    _zz_dataOut_payload_200_27;
  reg        [7:0]    _zz_dataOut_payload_201_6;
  reg        [7:0]    _zz_dataOut_payload_202_9;
  reg        [7:0]    _zz_dataOut_payload_203_6;
  reg        [7:0]    _zz_dataOut_payload_204_15;
  reg        [7:0]    _zz_dataOut_payload_205_6;
  reg        [7:0]    _zz_dataOut_payload_206_9;
  reg        [7:0]    _zz_dataOut_payload_207_6;
  reg        [7:0]    _zz_dataOut_payload_208_51;
  reg        [7:0]    _zz_dataOut_payload_209_6;
  reg        [7:0]    _zz_dataOut_payload_210_9;
  reg        [7:0]    _zz_dataOut_payload_211_6;
  reg        [7:0]    _zz_dataOut_payload_212_15;
  reg        [7:0]    _zz_dataOut_payload_213_6;
  reg        [7:0]    _zz_dataOut_payload_214_9;
  reg        [7:0]    _zz_dataOut_payload_215_6;
  reg        [7:0]    _zz_dataOut_payload_216_27;
  reg        [7:0]    _zz_dataOut_payload_217_6;
  reg        [7:0]    _zz_dataOut_payload_218_9;
  reg        [7:0]    _zz_dataOut_payload_219_6;
  reg        [7:0]    _zz_dataOut_payload_220_15;
  reg        [7:0]    _zz_dataOut_payload_221_6;
  reg        [7:0]    _zz_dataOut_payload_222_9;
  reg        [7:0]    _zz_dataOut_payload_223_6;
  reg        [7:0]    _zz_dataOut_payload_224_99;
  reg        [7:0]    _zz_dataOut_payload_225_6;
  reg        [7:0]    _zz_dataOut_payload_226_9;
  reg        [7:0]    _zz_dataOut_payload_227_6;
  reg        [7:0]    _zz_dataOut_payload_228_15;
  reg        [7:0]    _zz_dataOut_payload_229_6;
  reg        [7:0]    _zz_dataOut_payload_230_9;
  reg        [7:0]    _zz_dataOut_payload_231_6;
  reg        [7:0]    _zz_dataOut_payload_232_27;
  reg        [7:0]    _zz_dataOut_payload_233_6;
  reg        [7:0]    _zz_dataOut_payload_234_9;
  reg        [7:0]    _zz_dataOut_payload_235_6;
  reg        [7:0]    _zz_dataOut_payload_236_15;
  reg        [7:0]    _zz_dataOut_payload_237_6;
  reg        [7:0]    _zz_dataOut_payload_238_9;
  reg        [7:0]    _zz_dataOut_payload_239_6;
  reg        [7:0]    _zz_dataOut_payload_240_51;
  reg        [7:0]    _zz_dataOut_payload_241_6;
  reg        [7:0]    _zz_dataOut_payload_242_9;
  reg        [7:0]    _zz_dataOut_payload_243_6;
  reg        [7:0]    _zz_dataOut_payload_244_15;
  reg        [7:0]    _zz_dataOut_payload_245_6;
  reg        [7:0]    _zz_dataOut_payload_246_9;
  reg        [7:0]    _zz_dataOut_payload_247_6;
  reg        [7:0]    _zz_dataOut_payload_248_27;
  reg        [7:0]    _zz_dataOut_payload_249_6;
  reg        [7:0]    _zz_dataOut_payload_250_9;
  reg        [7:0]    _zz_dataOut_payload_251_6;
  reg        [7:0]    _zz_dataOut_payload_252_15;
  reg        [7:0]    _zz_dataOut_payload_253_6;
  reg        [7:0]    _zz_dataOut_payload_254_9;
  reg        [7:0]    _zz_dataOut_payload_255_6;
  reg        [7:0]    _zz_dataOut_payload_0_16644;
  reg        [7:0]    _zz_dataOut_payload_1_7;
  reg        [7:0]    _zz_dataOut_payload_2_10;
  reg        [7:0]    _zz_dataOut_payload_3_7;
  reg        [7:0]    _zz_dataOut_payload_4_16;
  reg        [7:0]    _zz_dataOut_payload_5_7;
  reg        [7:0]    _zz_dataOut_payload_6_10;
  reg        [7:0]    _zz_dataOut_payload_7_7;
  reg        [7:0]    _zz_dataOut_payload_8_28;
  reg        [7:0]    _zz_dataOut_payload_9_7;
  reg        [7:0]    _zz_dataOut_payload_10_10;
  reg        [7:0]    _zz_dataOut_payload_11_7;
  reg        [7:0]    _zz_dataOut_payload_12_16;
  reg        [7:0]    _zz_dataOut_payload_13_7;
  reg        [7:0]    _zz_dataOut_payload_14_10;
  reg        [7:0]    _zz_dataOut_payload_15_7;
  reg        [7:0]    _zz_dataOut_payload_16_52;
  reg        [7:0]    _zz_dataOut_payload_17_7;
  reg        [7:0]    _zz_dataOut_payload_18_10;
  reg        [7:0]    _zz_dataOut_payload_19_7;
  reg        [7:0]    _zz_dataOut_payload_20_16;
  reg        [7:0]    _zz_dataOut_payload_21_7;
  reg        [7:0]    _zz_dataOut_payload_22_10;
  reg        [7:0]    _zz_dataOut_payload_23_7;
  reg        [7:0]    _zz_dataOut_payload_24_28;
  reg        [7:0]    _zz_dataOut_payload_25_7;
  reg        [7:0]    _zz_dataOut_payload_26_10;
  reg        [7:0]    _zz_dataOut_payload_27_7;
  reg        [7:0]    _zz_dataOut_payload_28_16;
  reg        [7:0]    _zz_dataOut_payload_29_7;
  reg        [7:0]    _zz_dataOut_payload_30_10;
  reg        [7:0]    _zz_dataOut_payload_31_7;
  reg        [7:0]    _zz_dataOut_payload_32_100;
  reg        [7:0]    _zz_dataOut_payload_33_7;
  reg        [7:0]    _zz_dataOut_payload_34_10;
  reg        [7:0]    _zz_dataOut_payload_35_7;
  reg        [7:0]    _zz_dataOut_payload_36_16;
  reg        [7:0]    _zz_dataOut_payload_37_7;
  reg        [7:0]    _zz_dataOut_payload_38_10;
  reg        [7:0]    _zz_dataOut_payload_39_7;
  reg        [7:0]    _zz_dataOut_payload_40_28;
  reg        [7:0]    _zz_dataOut_payload_41_7;
  reg        [7:0]    _zz_dataOut_payload_42_10;
  reg        [7:0]    _zz_dataOut_payload_43_7;
  reg        [7:0]    _zz_dataOut_payload_44_16;
  reg        [7:0]    _zz_dataOut_payload_45_7;
  reg        [7:0]    _zz_dataOut_payload_46_10;
  reg        [7:0]    _zz_dataOut_payload_47_7;
  reg        [7:0]    _zz_dataOut_payload_48_52;
  reg        [7:0]    _zz_dataOut_payload_49_7;
  reg        [7:0]    _zz_dataOut_payload_50_10;
  reg        [7:0]    _zz_dataOut_payload_51_7;
  reg        [7:0]    _zz_dataOut_payload_52_16;
  reg        [7:0]    _zz_dataOut_payload_53_7;
  reg        [7:0]    _zz_dataOut_payload_54_10;
  reg        [7:0]    _zz_dataOut_payload_55_7;
  reg        [7:0]    _zz_dataOut_payload_56_28;
  reg        [7:0]    _zz_dataOut_payload_57_7;
  reg        [7:0]    _zz_dataOut_payload_58_10;
  reg        [7:0]    _zz_dataOut_payload_59_7;
  reg        [7:0]    _zz_dataOut_payload_60_16;
  reg        [7:0]    _zz_dataOut_payload_61_7;
  reg        [7:0]    _zz_dataOut_payload_62_10;
  reg        [7:0]    _zz_dataOut_payload_63_7;
  reg        [7:0]    _zz_dataOut_payload_64_196;
  reg        [7:0]    _zz_dataOut_payload_65_7;
  reg        [7:0]    _zz_dataOut_payload_66_10;
  reg        [7:0]    _zz_dataOut_payload_67_7;
  reg        [7:0]    _zz_dataOut_payload_68_16;
  reg        [7:0]    _zz_dataOut_payload_69_7;
  reg        [7:0]    _zz_dataOut_payload_70_10;
  reg        [7:0]    _zz_dataOut_payload_71_7;
  reg        [7:0]    _zz_dataOut_payload_72_28;
  reg        [7:0]    _zz_dataOut_payload_73_7;
  reg        [7:0]    _zz_dataOut_payload_74_10;
  reg        [7:0]    _zz_dataOut_payload_75_7;
  reg        [7:0]    _zz_dataOut_payload_76_16;
  reg        [7:0]    _zz_dataOut_payload_77_7;
  reg        [7:0]    _zz_dataOut_payload_78_10;
  reg        [7:0]    _zz_dataOut_payload_79_7;
  reg        [7:0]    _zz_dataOut_payload_80_52;
  reg        [7:0]    _zz_dataOut_payload_81_7;
  reg        [7:0]    _zz_dataOut_payload_82_10;
  reg        [7:0]    _zz_dataOut_payload_83_7;
  reg        [7:0]    _zz_dataOut_payload_84_16;
  reg        [7:0]    _zz_dataOut_payload_85_7;
  reg        [7:0]    _zz_dataOut_payload_86_10;
  reg        [7:0]    _zz_dataOut_payload_87_7;
  reg        [7:0]    _zz_dataOut_payload_88_28;
  reg        [7:0]    _zz_dataOut_payload_89_7;
  reg        [7:0]    _zz_dataOut_payload_90_10;
  reg        [7:0]    _zz_dataOut_payload_91_7;
  reg        [7:0]    _zz_dataOut_payload_92_16;
  reg        [7:0]    _zz_dataOut_payload_93_7;
  reg        [7:0]    _zz_dataOut_payload_94_10;
  reg        [7:0]    _zz_dataOut_payload_95_7;
  reg        [7:0]    _zz_dataOut_payload_96_100;
  reg        [7:0]    _zz_dataOut_payload_97_7;
  reg        [7:0]    _zz_dataOut_payload_98_10;
  reg        [7:0]    _zz_dataOut_payload_99_7;
  reg        [7:0]    _zz_dataOut_payload_100_16;
  reg        [7:0]    _zz_dataOut_payload_101_7;
  reg        [7:0]    _zz_dataOut_payload_102_10;
  reg        [7:0]    _zz_dataOut_payload_103_7;
  reg        [7:0]    _zz_dataOut_payload_104_28;
  reg        [7:0]    _zz_dataOut_payload_105_7;
  reg        [7:0]    _zz_dataOut_payload_106_10;
  reg        [7:0]    _zz_dataOut_payload_107_7;
  reg        [7:0]    _zz_dataOut_payload_108_16;
  reg        [7:0]    _zz_dataOut_payload_109_7;
  reg        [7:0]    _zz_dataOut_payload_110_10;
  reg        [7:0]    _zz_dataOut_payload_111_7;
  reg        [7:0]    _zz_dataOut_payload_112_52;
  reg        [7:0]    _zz_dataOut_payload_113_7;
  reg        [7:0]    _zz_dataOut_payload_114_10;
  reg        [7:0]    _zz_dataOut_payload_115_7;
  reg        [7:0]    _zz_dataOut_payload_116_16;
  reg        [7:0]    _zz_dataOut_payload_117_7;
  reg        [7:0]    _zz_dataOut_payload_118_10;
  reg        [7:0]    _zz_dataOut_payload_119_7;
  reg        [7:0]    _zz_dataOut_payload_120_28;
  reg        [7:0]    _zz_dataOut_payload_121_7;
  reg        [7:0]    _zz_dataOut_payload_122_10;
  reg        [7:0]    _zz_dataOut_payload_123_7;
  reg        [7:0]    _zz_dataOut_payload_124_16;
  reg        [7:0]    _zz_dataOut_payload_125_7;
  reg        [7:0]    _zz_dataOut_payload_126_10;
  reg        [7:0]    _zz_dataOut_payload_127_7;
  reg        [7:0]    _zz_dataOut_payload_128_388;
  reg        [7:0]    _zz_dataOut_payload_129_7;
  reg        [7:0]    _zz_dataOut_payload_130_10;
  reg        [7:0]    _zz_dataOut_payload_131_7;
  reg        [7:0]    _zz_dataOut_payload_132_16;
  reg        [7:0]    _zz_dataOut_payload_133_7;
  reg        [7:0]    _zz_dataOut_payload_134_10;
  reg        [7:0]    _zz_dataOut_payload_135_7;
  reg        [7:0]    _zz_dataOut_payload_136_28;
  reg        [7:0]    _zz_dataOut_payload_137_7;
  reg        [7:0]    _zz_dataOut_payload_138_10;
  reg        [7:0]    _zz_dataOut_payload_139_7;
  reg        [7:0]    _zz_dataOut_payload_140_16;
  reg        [7:0]    _zz_dataOut_payload_141_7;
  reg        [7:0]    _zz_dataOut_payload_142_10;
  reg        [7:0]    _zz_dataOut_payload_143_7;
  reg        [7:0]    _zz_dataOut_payload_144_52;
  reg        [7:0]    _zz_dataOut_payload_145_7;
  reg        [7:0]    _zz_dataOut_payload_146_10;
  reg        [7:0]    _zz_dataOut_payload_147_7;
  reg        [7:0]    _zz_dataOut_payload_148_16;
  reg        [7:0]    _zz_dataOut_payload_149_7;
  reg        [7:0]    _zz_dataOut_payload_150_10;
  reg        [7:0]    _zz_dataOut_payload_151_7;
  reg        [7:0]    _zz_dataOut_payload_152_28;
  reg        [7:0]    _zz_dataOut_payload_153_7;
  reg        [7:0]    _zz_dataOut_payload_154_10;
  reg        [7:0]    _zz_dataOut_payload_155_7;
  reg        [7:0]    _zz_dataOut_payload_156_16;
  reg        [7:0]    _zz_dataOut_payload_157_7;
  reg        [7:0]    _zz_dataOut_payload_158_10;
  reg        [7:0]    _zz_dataOut_payload_159_7;
  reg        [7:0]    _zz_dataOut_payload_160_100;
  reg        [7:0]    _zz_dataOut_payload_161_7;
  reg        [7:0]    _zz_dataOut_payload_162_10;
  reg        [7:0]    _zz_dataOut_payload_163_7;
  reg        [7:0]    _zz_dataOut_payload_164_16;
  reg        [7:0]    _zz_dataOut_payload_165_7;
  reg        [7:0]    _zz_dataOut_payload_166_10;
  reg        [7:0]    _zz_dataOut_payload_167_7;
  reg        [7:0]    _zz_dataOut_payload_168_28;
  reg        [7:0]    _zz_dataOut_payload_169_7;
  reg        [7:0]    _zz_dataOut_payload_170_10;
  reg        [7:0]    _zz_dataOut_payload_171_7;
  reg        [7:0]    _zz_dataOut_payload_172_16;
  reg        [7:0]    _zz_dataOut_payload_173_7;
  reg        [7:0]    _zz_dataOut_payload_174_10;
  reg        [7:0]    _zz_dataOut_payload_175_7;
  reg        [7:0]    _zz_dataOut_payload_176_52;
  reg        [7:0]    _zz_dataOut_payload_177_7;
  reg        [7:0]    _zz_dataOut_payload_178_10;
  reg        [7:0]    _zz_dataOut_payload_179_7;
  reg        [7:0]    _zz_dataOut_payload_180_16;
  reg        [7:0]    _zz_dataOut_payload_181_7;
  reg        [7:0]    _zz_dataOut_payload_182_10;
  reg        [7:0]    _zz_dataOut_payload_183_7;
  reg        [7:0]    _zz_dataOut_payload_184_28;
  reg        [7:0]    _zz_dataOut_payload_185_7;
  reg        [7:0]    _zz_dataOut_payload_186_10;
  reg        [7:0]    _zz_dataOut_payload_187_7;
  reg        [7:0]    _zz_dataOut_payload_188_16;
  reg        [7:0]    _zz_dataOut_payload_189_7;
  reg        [7:0]    _zz_dataOut_payload_190_10;
  reg        [7:0]    _zz_dataOut_payload_191_7;
  reg        [7:0]    _zz_dataOut_payload_192_196;
  reg        [7:0]    _zz_dataOut_payload_193_7;
  reg        [7:0]    _zz_dataOut_payload_194_10;
  reg        [7:0]    _zz_dataOut_payload_195_7;
  reg        [7:0]    _zz_dataOut_payload_196_16;
  reg        [7:0]    _zz_dataOut_payload_197_7;
  reg        [7:0]    _zz_dataOut_payload_198_10;
  reg        [7:0]    _zz_dataOut_payload_199_7;
  reg        [7:0]    _zz_dataOut_payload_200_28;
  reg        [7:0]    _zz_dataOut_payload_201_7;
  reg        [7:0]    _zz_dataOut_payload_202_10;
  reg        [7:0]    _zz_dataOut_payload_203_7;
  reg        [7:0]    _zz_dataOut_payload_204_16;
  reg        [7:0]    _zz_dataOut_payload_205_7;
  reg        [7:0]    _zz_dataOut_payload_206_10;
  reg        [7:0]    _zz_dataOut_payload_207_7;
  reg        [7:0]    _zz_dataOut_payload_208_52;
  reg        [7:0]    _zz_dataOut_payload_209_7;
  reg        [7:0]    _zz_dataOut_payload_210_10;
  reg        [7:0]    _zz_dataOut_payload_211_7;
  reg        [7:0]    _zz_dataOut_payload_212_16;
  reg        [7:0]    _zz_dataOut_payload_213_7;
  reg        [7:0]    _zz_dataOut_payload_214_10;
  reg        [7:0]    _zz_dataOut_payload_215_7;
  reg        [7:0]    _zz_dataOut_payload_216_28;
  reg        [7:0]    _zz_dataOut_payload_217_7;
  reg        [7:0]    _zz_dataOut_payload_218_10;
  reg        [7:0]    _zz_dataOut_payload_219_7;
  reg        [7:0]    _zz_dataOut_payload_220_16;
  reg        [7:0]    _zz_dataOut_payload_221_7;
  reg        [7:0]    _zz_dataOut_payload_222_10;
  reg        [7:0]    _zz_dataOut_payload_223_7;
  reg        [7:0]    _zz_dataOut_payload_224_100;
  reg        [7:0]    _zz_dataOut_payload_225_7;
  reg        [7:0]    _zz_dataOut_payload_226_10;
  reg        [7:0]    _zz_dataOut_payload_227_7;
  reg        [7:0]    _zz_dataOut_payload_228_16;
  reg        [7:0]    _zz_dataOut_payload_229_7;
  reg        [7:0]    _zz_dataOut_payload_230_10;
  reg        [7:0]    _zz_dataOut_payload_231_7;
  reg        [7:0]    _zz_dataOut_payload_232_28;
  reg        [7:0]    _zz_dataOut_payload_233_7;
  reg        [7:0]    _zz_dataOut_payload_234_10;
  reg        [7:0]    _zz_dataOut_payload_235_7;
  reg        [7:0]    _zz_dataOut_payload_236_16;
  reg        [7:0]    _zz_dataOut_payload_237_7;
  reg        [7:0]    _zz_dataOut_payload_238_10;
  reg        [7:0]    _zz_dataOut_payload_239_7;
  reg        [7:0]    _zz_dataOut_payload_240_52;
  reg        [7:0]    _zz_dataOut_payload_241_7;
  reg        [7:0]    _zz_dataOut_payload_242_10;
  reg        [7:0]    _zz_dataOut_payload_243_7;
  reg        [7:0]    _zz_dataOut_payload_244_16;
  reg        [7:0]    _zz_dataOut_payload_245_7;
  reg        [7:0]    _zz_dataOut_payload_246_10;
  reg        [7:0]    _zz_dataOut_payload_247_7;
  reg        [7:0]    _zz_dataOut_payload_248_28;
  reg        [7:0]    _zz_dataOut_payload_249_7;
  reg        [7:0]    _zz_dataOut_payload_250_10;
  reg        [7:0]    _zz_dataOut_payload_251_7;
  reg        [7:0]    _zz_dataOut_payload_252_16;
  reg        [7:0]    _zz_dataOut_payload_253_7;
  reg        [7:0]    _zz_dataOut_payload_254_10;
  reg        [7:0]    _zz_dataOut_payload_255_7;
  reg                 dataIn_valid_delay_1;
  reg                 dataIn_valid_delay_2;
  reg                 dataIn_valid_delay_3;
  reg                 dataIn_valid_delay_4;
  reg                 dataIn_valid_delay_5;
  reg                 dataIn_valid_delay_6;
  reg                 dataIn_valid_delay_7;
  reg                 dataIn_valid_delay_8;
  reg                 dataIn_valid_delay_9;
  reg                 dataIn_valid_delay_10;
  reg                 dataIn_valid_delay_11;
  reg                 dataIn_valid_delay_12;
  reg                 dataIn_valid_delay_13;
  reg                 dataIn_valid_delay_14;
  reg                 dataIn_valid_delay_15;
  reg                 dataIn_valid_delay_16;
  reg                 dataIn_valid_delay_17;
  reg                 dataIn_valid_delay_18;
  reg                 dataIn_valid_delay_19;
  reg                 dataIn_valid_delay_20;
  reg                 dataIn_valid_delay_21;
  reg                 dataIn_valid_delay_22;
  reg                 dataIn_valid_delay_23;
  reg                 dataIn_valid_delay_24;
  reg                 dataIn_valid_delay_25;
  reg                 dataIn_valid_delay_26;
  reg                 dataIn_valid_delay_27;
  reg                 dataIn_valid_delay_28;
  reg                 dataIn_valid_delay_29;
  reg                 dataIn_valid_delay_30;
  reg                 dataIn_valid_delay_31;
  reg                 dataIn_valid_delay_32;
  reg                 dataIn_valid_delay_33;
  reg                 dataIn_valid_delay_34;
  reg                 dataIn_valid_delay_35;
  reg                 dataIn_valid_delay_36;

  assign _zz_dataOut_payload_0 = (dataIn_payload_0 < dataIn_payload_1);
  assign _zz_dataOut_payload_0_1 = (dataIn_payload_2 < dataIn_payload_3);
  assign _zz_dataOut_payload_0_2 = (dataIn_payload_4 < dataIn_payload_5);
  assign _zz_dataOut_payload_0_3 = (dataIn_payload_6 < dataIn_payload_7);
  assign _zz_dataOut_payload_0_4 = (dataIn_payload_8 < dataIn_payload_9);
  assign _zz_dataOut_payload_0_5 = (dataIn_payload_10 < dataIn_payload_11);
  assign _zz_dataOut_payload_0_6 = (dataIn_payload_12 < dataIn_payload_13);
  assign _zz_dataOut_payload_0_7 = (dataIn_payload_14 < dataIn_payload_15);
  assign _zz_dataOut_payload_0_8 = (dataIn_payload_16 < dataIn_payload_17);
  assign _zz_dataOut_payload_0_9 = (dataIn_payload_18 < dataIn_payload_19);
  assign _zz_dataOut_payload_0_10 = (dataIn_payload_20 < dataIn_payload_21);
  assign _zz_dataOut_payload_0_11 = (dataIn_payload_22 < dataIn_payload_23);
  assign _zz_dataOut_payload_0_12 = (dataIn_payload_24 < dataIn_payload_25);
  assign _zz_dataOut_payload_0_13 = (dataIn_payload_26 < dataIn_payload_27);
  assign _zz_dataOut_payload_0_14 = (dataIn_payload_28 < dataIn_payload_29);
  assign _zz_dataOut_payload_0_15 = (dataIn_payload_30 < dataIn_payload_31);
  assign _zz_dataOut_payload_0_16 = (dataIn_payload_32 < dataIn_payload_33);
  assign _zz_dataOut_payload_0_17 = (dataIn_payload_34 < dataIn_payload_35);
  assign _zz_dataOut_payload_0_18 = (dataIn_payload_36 < dataIn_payload_37);
  assign _zz_dataOut_payload_0_19 = (dataIn_payload_38 < dataIn_payload_39);
  assign _zz_dataOut_payload_0_20 = (dataIn_payload_40 < dataIn_payload_41);
  assign _zz_dataOut_payload_0_21 = (dataIn_payload_42 < dataIn_payload_43);
  assign _zz_dataOut_payload_0_22 = (dataIn_payload_44 < dataIn_payload_45);
  assign _zz_dataOut_payload_0_23 = (dataIn_payload_46 < dataIn_payload_47);
  assign _zz_dataOut_payload_0_24 = (dataIn_payload_48 < dataIn_payload_49);
  assign _zz_dataOut_payload_0_25 = (dataIn_payload_50 < dataIn_payload_51);
  assign _zz_dataOut_payload_0_26 = (dataIn_payload_52 < dataIn_payload_53);
  assign _zz_dataOut_payload_0_27 = (dataIn_payload_54 < dataIn_payload_55);
  assign _zz_dataOut_payload_0_28 = (dataIn_payload_56 < dataIn_payload_57);
  assign _zz_dataOut_payload_0_29 = (dataIn_payload_58 < dataIn_payload_59);
  assign _zz_dataOut_payload_0_30 = (dataIn_payload_60 < dataIn_payload_61);
  assign _zz_dataOut_payload_0_31 = (dataIn_payload_62 < dataIn_payload_63);
  assign _zz_dataOut_payload_0_32 = (dataIn_payload_64 < dataIn_payload_65);
  assign _zz_dataOut_payload_0_33 = (dataIn_payload_66 < dataIn_payload_67);
  assign _zz_dataOut_payload_0_34 = (dataIn_payload_68 < dataIn_payload_69);
  assign _zz_dataOut_payload_0_35 = (dataIn_payload_70 < dataIn_payload_71);
  assign _zz_dataOut_payload_0_36 = (dataIn_payload_72 < dataIn_payload_73);
  assign _zz_dataOut_payload_0_37 = (dataIn_payload_74 < dataIn_payload_75);
  assign _zz_dataOut_payload_0_38 = (dataIn_payload_76 < dataIn_payload_77);
  assign _zz_dataOut_payload_0_39 = (dataIn_payload_78 < dataIn_payload_79);
  assign _zz_dataOut_payload_0_40 = (dataIn_payload_80 < dataIn_payload_81);
  assign _zz_dataOut_payload_0_41 = (dataIn_payload_82 < dataIn_payload_83);
  assign _zz_dataOut_payload_0_42 = (dataIn_payload_84 < dataIn_payload_85);
  assign _zz_dataOut_payload_0_43 = (dataIn_payload_86 < dataIn_payload_87);
  assign _zz_dataOut_payload_0_44 = (dataIn_payload_88 < dataIn_payload_89);
  assign _zz_dataOut_payload_0_45 = (dataIn_payload_90 < dataIn_payload_91);
  assign _zz_dataOut_payload_0_46 = (dataIn_payload_92 < dataIn_payload_93);
  assign _zz_dataOut_payload_0_47 = (dataIn_payload_94 < dataIn_payload_95);
  assign _zz_dataOut_payload_0_48 = (dataIn_payload_96 < dataIn_payload_97);
  assign _zz_dataOut_payload_0_49 = (dataIn_payload_98 < dataIn_payload_99);
  assign _zz_dataOut_payload_0_50 = (dataIn_payload_100 < dataIn_payload_101);
  assign _zz_dataOut_payload_0_51 = (dataIn_payload_102 < dataIn_payload_103);
  assign _zz_dataOut_payload_0_52 = (dataIn_payload_104 < dataIn_payload_105);
  assign _zz_dataOut_payload_0_53 = (dataIn_payload_106 < dataIn_payload_107);
  assign _zz_dataOut_payload_0_54 = (dataIn_payload_108 < dataIn_payload_109);
  assign _zz_dataOut_payload_0_55 = (dataIn_payload_110 < dataIn_payload_111);
  assign _zz_dataOut_payload_0_56 = (dataIn_payload_112 < dataIn_payload_113);
  assign _zz_dataOut_payload_0_57 = (dataIn_payload_114 < dataIn_payload_115);
  assign _zz_dataOut_payload_0_58 = (dataIn_payload_116 < dataIn_payload_117);
  assign _zz_dataOut_payload_0_59 = (dataIn_payload_118 < dataIn_payload_119);
  assign _zz_dataOut_payload_0_60 = (dataIn_payload_120 < dataIn_payload_121);
  assign _zz_dataOut_payload_0_61 = (dataIn_payload_122 < dataIn_payload_123);
  assign _zz_dataOut_payload_0_62 = (dataIn_payload_124 < dataIn_payload_125);
  assign _zz_dataOut_payload_0_63 = (dataIn_payload_126 < dataIn_payload_127);
  assign _zz_dataOut_payload_0_64 = (dataIn_payload_128 < dataIn_payload_129);
  assign _zz_dataOut_payload_0_65 = (dataIn_payload_130 < dataIn_payload_131);
  assign _zz_dataOut_payload_0_66 = (dataIn_payload_132 < dataIn_payload_133);
  assign _zz_dataOut_payload_0_67 = (dataIn_payload_134 < dataIn_payload_135);
  assign _zz_dataOut_payload_0_68 = (dataIn_payload_136 < dataIn_payload_137);
  assign _zz_dataOut_payload_0_69 = (dataIn_payload_138 < dataIn_payload_139);
  assign _zz_dataOut_payload_0_70 = (dataIn_payload_140 < dataIn_payload_141);
  assign _zz_dataOut_payload_0_71 = (dataIn_payload_142 < dataIn_payload_143);
  assign _zz_dataOut_payload_0_72 = (dataIn_payload_144 < dataIn_payload_145);
  assign _zz_dataOut_payload_0_73 = (dataIn_payload_146 < dataIn_payload_147);
  assign _zz_dataOut_payload_0_74 = (dataIn_payload_148 < dataIn_payload_149);
  assign _zz_dataOut_payload_0_75 = (dataIn_payload_150 < dataIn_payload_151);
  assign _zz_dataOut_payload_0_76 = (dataIn_payload_152 < dataIn_payload_153);
  assign _zz_dataOut_payload_0_77 = (dataIn_payload_154 < dataIn_payload_155);
  assign _zz_dataOut_payload_0_78 = (dataIn_payload_156 < dataIn_payload_157);
  assign _zz_dataOut_payload_0_79 = (dataIn_payload_158 < dataIn_payload_159);
  assign _zz_dataOut_payload_0_80 = (dataIn_payload_160 < dataIn_payload_161);
  assign _zz_dataOut_payload_0_81 = (dataIn_payload_162 < dataIn_payload_163);
  assign _zz_dataOut_payload_0_82 = (dataIn_payload_164 < dataIn_payload_165);
  assign _zz_dataOut_payload_0_83 = (dataIn_payload_166 < dataIn_payload_167);
  assign _zz_dataOut_payload_0_84 = (dataIn_payload_168 < dataIn_payload_169);
  assign _zz_dataOut_payload_0_85 = (dataIn_payload_170 < dataIn_payload_171);
  assign _zz_dataOut_payload_0_86 = (dataIn_payload_172 < dataIn_payload_173);
  assign _zz_dataOut_payload_0_87 = (dataIn_payload_174 < dataIn_payload_175);
  assign _zz_dataOut_payload_0_88 = (dataIn_payload_176 < dataIn_payload_177);
  assign _zz_dataOut_payload_0_89 = (dataIn_payload_178 < dataIn_payload_179);
  assign _zz_dataOut_payload_0_90 = (dataIn_payload_180 < dataIn_payload_181);
  assign _zz_dataOut_payload_0_91 = (dataIn_payload_182 < dataIn_payload_183);
  assign _zz_dataOut_payload_0_92 = (dataIn_payload_184 < dataIn_payload_185);
  assign _zz_dataOut_payload_0_93 = (dataIn_payload_186 < dataIn_payload_187);
  assign _zz_dataOut_payload_0_94 = (dataIn_payload_188 < dataIn_payload_189);
  assign _zz_dataOut_payload_0_95 = (dataIn_payload_190 < dataIn_payload_191);
  assign _zz_dataOut_payload_0_96 = (dataIn_payload_192 < dataIn_payload_193);
  assign _zz_dataOut_payload_0_97 = (dataIn_payload_194 < dataIn_payload_195);
  assign _zz_dataOut_payload_0_98 = (dataIn_payload_196 < dataIn_payload_197);
  assign _zz_dataOut_payload_0_99 = (dataIn_payload_198 < dataIn_payload_199);
  assign _zz_dataOut_payload_0_100 = (dataIn_payload_200 < dataIn_payload_201);
  assign _zz_dataOut_payload_0_101 = (dataIn_payload_202 < dataIn_payload_203);
  assign _zz_dataOut_payload_0_102 = (dataIn_payload_204 < dataIn_payload_205);
  assign _zz_dataOut_payload_0_103 = (dataIn_payload_206 < dataIn_payload_207);
  assign _zz_dataOut_payload_0_104 = (dataIn_payload_208 < dataIn_payload_209);
  assign _zz_dataOut_payload_0_105 = (dataIn_payload_210 < dataIn_payload_211);
  assign _zz_dataOut_payload_0_106 = (dataIn_payload_212 < dataIn_payload_213);
  assign _zz_dataOut_payload_0_107 = (dataIn_payload_214 < dataIn_payload_215);
  assign _zz_dataOut_payload_0_108 = (dataIn_payload_216 < dataIn_payload_217);
  assign _zz_dataOut_payload_0_109 = (dataIn_payload_218 < dataIn_payload_219);
  assign _zz_dataOut_payload_0_110 = (dataIn_payload_220 < dataIn_payload_221);
  assign _zz_dataOut_payload_0_111 = (dataIn_payload_222 < dataIn_payload_223);
  assign _zz_dataOut_payload_0_112 = (dataIn_payload_224 < dataIn_payload_225);
  assign _zz_dataOut_payload_0_113 = (dataIn_payload_226 < dataIn_payload_227);
  assign _zz_dataOut_payload_0_114 = (dataIn_payload_228 < dataIn_payload_229);
  assign _zz_dataOut_payload_0_115 = (dataIn_payload_230 < dataIn_payload_231);
  assign _zz_dataOut_payload_0_116 = (dataIn_payload_232 < dataIn_payload_233);
  assign _zz_dataOut_payload_0_117 = (dataIn_payload_234 < dataIn_payload_235);
  assign _zz_dataOut_payload_0_118 = (dataIn_payload_236 < dataIn_payload_237);
  assign _zz_dataOut_payload_0_119 = (dataIn_payload_238 < dataIn_payload_239);
  assign _zz_dataOut_payload_0_120 = (dataIn_payload_240 < dataIn_payload_241);
  assign _zz_dataOut_payload_0_121 = (dataIn_payload_242 < dataIn_payload_243);
  assign _zz_dataOut_payload_0_122 = (dataIn_payload_244 < dataIn_payload_245);
  assign _zz_dataOut_payload_0_123 = (dataIn_payload_246 < dataIn_payload_247);
  assign _zz_dataOut_payload_0_124 = (dataIn_payload_248 < dataIn_payload_249);
  assign _zz_dataOut_payload_0_125 = (dataIn_payload_250 < dataIn_payload_251);
  assign _zz_dataOut_payload_0_126 = (dataIn_payload_252 < dataIn_payload_253);
  assign _zz_dataOut_payload_0_127 = (dataIn_payload_254 < dataIn_payload_255);
  assign _zz_dataOut_payload_0_384 = (_zz_dataOut_payload_0_128 < _zz_dataOut_payload_0_131);
  assign _zz_dataOut_payload_0_385 = (_zz_dataOut_payload_0_384 ? _zz_dataOut_payload_0_128 : _zz_dataOut_payload_0_131);
  assign _zz_dataOut_payload_0_386 = (_zz_dataOut_payload_0_384 ? _zz_dataOut_payload_0_131 : _zz_dataOut_payload_0_128);
  assign _zz_dataOut_payload_0_387 = (_zz_dataOut_payload_0_129 < _zz_dataOut_payload_0_130);
  assign _zz_dataOut_payload_0_388 = (_zz_dataOut_payload_0_387 ? _zz_dataOut_payload_0_129 : _zz_dataOut_payload_0_130);
  assign _zz_dataOut_payload_0_389 = (_zz_dataOut_payload_0_387 ? _zz_dataOut_payload_0_130 : _zz_dataOut_payload_0_129);
  assign _zz_dataOut_payload_0_390 = (_zz_dataOut_payload_0_385 < _zz_dataOut_payload_0_388);
  assign _zz_dataOut_payload_0_391 = (_zz_dataOut_payload_0_389 < _zz_dataOut_payload_0_386);
  assign _zz_dataOut_payload_0_396 = (_zz_dataOut_payload_0_132 < _zz_dataOut_payload_0_135);
  assign _zz_dataOut_payload_0_397 = (_zz_dataOut_payload_0_396 ? _zz_dataOut_payload_0_132 : _zz_dataOut_payload_0_135);
  assign _zz_dataOut_payload_0_398 = (_zz_dataOut_payload_0_396 ? _zz_dataOut_payload_0_135 : _zz_dataOut_payload_0_132);
  assign _zz_dataOut_payload_0_399 = (_zz_dataOut_payload_0_133 < _zz_dataOut_payload_0_134);
  assign _zz_dataOut_payload_0_400 = (_zz_dataOut_payload_0_399 ? _zz_dataOut_payload_0_133 : _zz_dataOut_payload_0_134);
  assign _zz_dataOut_payload_0_401 = (_zz_dataOut_payload_0_399 ? _zz_dataOut_payload_0_134 : _zz_dataOut_payload_0_133);
  assign _zz_dataOut_payload_0_402 = (_zz_dataOut_payload_0_397 < _zz_dataOut_payload_0_400);
  assign _zz_dataOut_payload_0_403 = (_zz_dataOut_payload_0_401 < _zz_dataOut_payload_0_398);
  assign _zz_dataOut_payload_0_408 = (_zz_dataOut_payload_0_136 < _zz_dataOut_payload_0_139);
  assign _zz_dataOut_payload_0_409 = (_zz_dataOut_payload_0_408 ? _zz_dataOut_payload_0_136 : _zz_dataOut_payload_0_139);
  assign _zz_dataOut_payload_0_410 = (_zz_dataOut_payload_0_408 ? _zz_dataOut_payload_0_139 : _zz_dataOut_payload_0_136);
  assign _zz_dataOut_payload_0_411 = (_zz_dataOut_payload_0_137 < _zz_dataOut_payload_0_138);
  assign _zz_dataOut_payload_0_412 = (_zz_dataOut_payload_0_411 ? _zz_dataOut_payload_0_137 : _zz_dataOut_payload_0_138);
  assign _zz_dataOut_payload_0_413 = (_zz_dataOut_payload_0_411 ? _zz_dataOut_payload_0_138 : _zz_dataOut_payload_0_137);
  assign _zz_dataOut_payload_0_414 = (_zz_dataOut_payload_0_409 < _zz_dataOut_payload_0_412);
  assign _zz_dataOut_payload_0_415 = (_zz_dataOut_payload_0_413 < _zz_dataOut_payload_0_410);
  assign _zz_dataOut_payload_0_420 = (_zz_dataOut_payload_0_140 < _zz_dataOut_payload_0_143);
  assign _zz_dataOut_payload_0_421 = (_zz_dataOut_payload_0_420 ? _zz_dataOut_payload_0_140 : _zz_dataOut_payload_0_143);
  assign _zz_dataOut_payload_0_422 = (_zz_dataOut_payload_0_420 ? _zz_dataOut_payload_0_143 : _zz_dataOut_payload_0_140);
  assign _zz_dataOut_payload_0_423 = (_zz_dataOut_payload_0_141 < _zz_dataOut_payload_0_142);
  assign _zz_dataOut_payload_0_424 = (_zz_dataOut_payload_0_423 ? _zz_dataOut_payload_0_141 : _zz_dataOut_payload_0_142);
  assign _zz_dataOut_payload_0_425 = (_zz_dataOut_payload_0_423 ? _zz_dataOut_payload_0_142 : _zz_dataOut_payload_0_141);
  assign _zz_dataOut_payload_0_426 = (_zz_dataOut_payload_0_421 < _zz_dataOut_payload_0_424);
  assign _zz_dataOut_payload_0_427 = (_zz_dataOut_payload_0_425 < _zz_dataOut_payload_0_422);
  assign _zz_dataOut_payload_0_432 = (_zz_dataOut_payload_0_144 < _zz_dataOut_payload_0_147);
  assign _zz_dataOut_payload_0_433 = (_zz_dataOut_payload_0_432 ? _zz_dataOut_payload_0_144 : _zz_dataOut_payload_0_147);
  assign _zz_dataOut_payload_0_434 = (_zz_dataOut_payload_0_432 ? _zz_dataOut_payload_0_147 : _zz_dataOut_payload_0_144);
  assign _zz_dataOut_payload_0_435 = (_zz_dataOut_payload_0_145 < _zz_dataOut_payload_0_146);
  assign _zz_dataOut_payload_0_436 = (_zz_dataOut_payload_0_435 ? _zz_dataOut_payload_0_145 : _zz_dataOut_payload_0_146);
  assign _zz_dataOut_payload_0_437 = (_zz_dataOut_payload_0_435 ? _zz_dataOut_payload_0_146 : _zz_dataOut_payload_0_145);
  assign _zz_dataOut_payload_0_438 = (_zz_dataOut_payload_0_433 < _zz_dataOut_payload_0_436);
  assign _zz_dataOut_payload_0_439 = (_zz_dataOut_payload_0_437 < _zz_dataOut_payload_0_434);
  assign _zz_dataOut_payload_0_444 = (_zz_dataOut_payload_0_148 < _zz_dataOut_payload_0_151);
  assign _zz_dataOut_payload_0_445 = (_zz_dataOut_payload_0_444 ? _zz_dataOut_payload_0_148 : _zz_dataOut_payload_0_151);
  assign _zz_dataOut_payload_0_446 = (_zz_dataOut_payload_0_444 ? _zz_dataOut_payload_0_151 : _zz_dataOut_payload_0_148);
  assign _zz_dataOut_payload_0_447 = (_zz_dataOut_payload_0_149 < _zz_dataOut_payload_0_150);
  assign _zz_dataOut_payload_0_448 = (_zz_dataOut_payload_0_447 ? _zz_dataOut_payload_0_149 : _zz_dataOut_payload_0_150);
  assign _zz_dataOut_payload_0_449 = (_zz_dataOut_payload_0_447 ? _zz_dataOut_payload_0_150 : _zz_dataOut_payload_0_149);
  assign _zz_dataOut_payload_0_450 = (_zz_dataOut_payload_0_445 < _zz_dataOut_payload_0_448);
  assign _zz_dataOut_payload_0_451 = (_zz_dataOut_payload_0_449 < _zz_dataOut_payload_0_446);
  assign _zz_dataOut_payload_0_456 = (_zz_dataOut_payload_0_152 < _zz_dataOut_payload_0_155);
  assign _zz_dataOut_payload_0_457 = (_zz_dataOut_payload_0_456 ? _zz_dataOut_payload_0_152 : _zz_dataOut_payload_0_155);
  assign _zz_dataOut_payload_0_458 = (_zz_dataOut_payload_0_456 ? _zz_dataOut_payload_0_155 : _zz_dataOut_payload_0_152);
  assign _zz_dataOut_payload_0_459 = (_zz_dataOut_payload_0_153 < _zz_dataOut_payload_0_154);
  assign _zz_dataOut_payload_0_460 = (_zz_dataOut_payload_0_459 ? _zz_dataOut_payload_0_153 : _zz_dataOut_payload_0_154);
  assign _zz_dataOut_payload_0_461 = (_zz_dataOut_payload_0_459 ? _zz_dataOut_payload_0_154 : _zz_dataOut_payload_0_153);
  assign _zz_dataOut_payload_0_462 = (_zz_dataOut_payload_0_457 < _zz_dataOut_payload_0_460);
  assign _zz_dataOut_payload_0_463 = (_zz_dataOut_payload_0_461 < _zz_dataOut_payload_0_458);
  assign _zz_dataOut_payload_0_468 = (_zz_dataOut_payload_0_156 < _zz_dataOut_payload_0_159);
  assign _zz_dataOut_payload_0_469 = (_zz_dataOut_payload_0_468 ? _zz_dataOut_payload_0_156 : _zz_dataOut_payload_0_159);
  assign _zz_dataOut_payload_0_470 = (_zz_dataOut_payload_0_468 ? _zz_dataOut_payload_0_159 : _zz_dataOut_payload_0_156);
  assign _zz_dataOut_payload_0_471 = (_zz_dataOut_payload_0_157 < _zz_dataOut_payload_0_158);
  assign _zz_dataOut_payload_0_472 = (_zz_dataOut_payload_0_471 ? _zz_dataOut_payload_0_157 : _zz_dataOut_payload_0_158);
  assign _zz_dataOut_payload_0_473 = (_zz_dataOut_payload_0_471 ? _zz_dataOut_payload_0_158 : _zz_dataOut_payload_0_157);
  assign _zz_dataOut_payload_0_474 = (_zz_dataOut_payload_0_469 < _zz_dataOut_payload_0_472);
  assign _zz_dataOut_payload_0_475 = (_zz_dataOut_payload_0_473 < _zz_dataOut_payload_0_470);
  assign _zz_dataOut_payload_0_480 = (_zz_dataOut_payload_0_160 < _zz_dataOut_payload_0_163);
  assign _zz_dataOut_payload_0_481 = (_zz_dataOut_payload_0_480 ? _zz_dataOut_payload_0_160 : _zz_dataOut_payload_0_163);
  assign _zz_dataOut_payload_0_482 = (_zz_dataOut_payload_0_480 ? _zz_dataOut_payload_0_163 : _zz_dataOut_payload_0_160);
  assign _zz_dataOut_payload_0_483 = (_zz_dataOut_payload_0_161 < _zz_dataOut_payload_0_162);
  assign _zz_dataOut_payload_0_484 = (_zz_dataOut_payload_0_483 ? _zz_dataOut_payload_0_161 : _zz_dataOut_payload_0_162);
  assign _zz_dataOut_payload_0_485 = (_zz_dataOut_payload_0_483 ? _zz_dataOut_payload_0_162 : _zz_dataOut_payload_0_161);
  assign _zz_dataOut_payload_0_486 = (_zz_dataOut_payload_0_481 < _zz_dataOut_payload_0_484);
  assign _zz_dataOut_payload_0_487 = (_zz_dataOut_payload_0_485 < _zz_dataOut_payload_0_482);
  assign _zz_dataOut_payload_0_492 = (_zz_dataOut_payload_0_164 < _zz_dataOut_payload_0_167);
  assign _zz_dataOut_payload_0_493 = (_zz_dataOut_payload_0_492 ? _zz_dataOut_payload_0_164 : _zz_dataOut_payload_0_167);
  assign _zz_dataOut_payload_0_494 = (_zz_dataOut_payload_0_492 ? _zz_dataOut_payload_0_167 : _zz_dataOut_payload_0_164);
  assign _zz_dataOut_payload_0_495 = (_zz_dataOut_payload_0_165 < _zz_dataOut_payload_0_166);
  assign _zz_dataOut_payload_0_496 = (_zz_dataOut_payload_0_495 ? _zz_dataOut_payload_0_165 : _zz_dataOut_payload_0_166);
  assign _zz_dataOut_payload_0_497 = (_zz_dataOut_payload_0_495 ? _zz_dataOut_payload_0_166 : _zz_dataOut_payload_0_165);
  assign _zz_dataOut_payload_0_498 = (_zz_dataOut_payload_0_493 < _zz_dataOut_payload_0_496);
  assign _zz_dataOut_payload_0_499 = (_zz_dataOut_payload_0_497 < _zz_dataOut_payload_0_494);
  assign _zz_dataOut_payload_0_504 = (_zz_dataOut_payload_0_168 < _zz_dataOut_payload_0_171);
  assign _zz_dataOut_payload_0_505 = (_zz_dataOut_payload_0_504 ? _zz_dataOut_payload_0_168 : _zz_dataOut_payload_0_171);
  assign _zz_dataOut_payload_0_506 = (_zz_dataOut_payload_0_504 ? _zz_dataOut_payload_0_171 : _zz_dataOut_payload_0_168);
  assign _zz_dataOut_payload_0_507 = (_zz_dataOut_payload_0_169 < _zz_dataOut_payload_0_170);
  assign _zz_dataOut_payload_0_508 = (_zz_dataOut_payload_0_507 ? _zz_dataOut_payload_0_169 : _zz_dataOut_payload_0_170);
  assign _zz_dataOut_payload_0_509 = (_zz_dataOut_payload_0_507 ? _zz_dataOut_payload_0_170 : _zz_dataOut_payload_0_169);
  assign _zz_dataOut_payload_0_510 = (_zz_dataOut_payload_0_505 < _zz_dataOut_payload_0_508);
  assign _zz_dataOut_payload_0_511 = (_zz_dataOut_payload_0_509 < _zz_dataOut_payload_0_506);
  assign _zz_dataOut_payload_0_516 = (_zz_dataOut_payload_0_172 < _zz_dataOut_payload_0_175);
  assign _zz_dataOut_payload_0_517 = (_zz_dataOut_payload_0_516 ? _zz_dataOut_payload_0_172 : _zz_dataOut_payload_0_175);
  assign _zz_dataOut_payload_0_518 = (_zz_dataOut_payload_0_516 ? _zz_dataOut_payload_0_175 : _zz_dataOut_payload_0_172);
  assign _zz_dataOut_payload_0_519 = (_zz_dataOut_payload_0_173 < _zz_dataOut_payload_0_174);
  assign _zz_dataOut_payload_0_520 = (_zz_dataOut_payload_0_519 ? _zz_dataOut_payload_0_173 : _zz_dataOut_payload_0_174);
  assign _zz_dataOut_payload_0_521 = (_zz_dataOut_payload_0_519 ? _zz_dataOut_payload_0_174 : _zz_dataOut_payload_0_173);
  assign _zz_dataOut_payload_0_522 = (_zz_dataOut_payload_0_517 < _zz_dataOut_payload_0_520);
  assign _zz_dataOut_payload_0_523 = (_zz_dataOut_payload_0_521 < _zz_dataOut_payload_0_518);
  assign _zz_dataOut_payload_0_528 = (_zz_dataOut_payload_0_176 < _zz_dataOut_payload_0_179);
  assign _zz_dataOut_payload_0_529 = (_zz_dataOut_payload_0_528 ? _zz_dataOut_payload_0_176 : _zz_dataOut_payload_0_179);
  assign _zz_dataOut_payload_0_530 = (_zz_dataOut_payload_0_528 ? _zz_dataOut_payload_0_179 : _zz_dataOut_payload_0_176);
  assign _zz_dataOut_payload_0_531 = (_zz_dataOut_payload_0_177 < _zz_dataOut_payload_0_178);
  assign _zz_dataOut_payload_0_532 = (_zz_dataOut_payload_0_531 ? _zz_dataOut_payload_0_177 : _zz_dataOut_payload_0_178);
  assign _zz_dataOut_payload_0_533 = (_zz_dataOut_payload_0_531 ? _zz_dataOut_payload_0_178 : _zz_dataOut_payload_0_177);
  assign _zz_dataOut_payload_0_534 = (_zz_dataOut_payload_0_529 < _zz_dataOut_payload_0_532);
  assign _zz_dataOut_payload_0_535 = (_zz_dataOut_payload_0_533 < _zz_dataOut_payload_0_530);
  assign _zz_dataOut_payload_0_540 = (_zz_dataOut_payload_0_180 < _zz_dataOut_payload_0_183);
  assign _zz_dataOut_payload_0_541 = (_zz_dataOut_payload_0_540 ? _zz_dataOut_payload_0_180 : _zz_dataOut_payload_0_183);
  assign _zz_dataOut_payload_0_542 = (_zz_dataOut_payload_0_540 ? _zz_dataOut_payload_0_183 : _zz_dataOut_payload_0_180);
  assign _zz_dataOut_payload_0_543 = (_zz_dataOut_payload_0_181 < _zz_dataOut_payload_0_182);
  assign _zz_dataOut_payload_0_544 = (_zz_dataOut_payload_0_543 ? _zz_dataOut_payload_0_181 : _zz_dataOut_payload_0_182);
  assign _zz_dataOut_payload_0_545 = (_zz_dataOut_payload_0_543 ? _zz_dataOut_payload_0_182 : _zz_dataOut_payload_0_181);
  assign _zz_dataOut_payload_0_546 = (_zz_dataOut_payload_0_541 < _zz_dataOut_payload_0_544);
  assign _zz_dataOut_payload_0_547 = (_zz_dataOut_payload_0_545 < _zz_dataOut_payload_0_542);
  assign _zz_dataOut_payload_0_552 = (_zz_dataOut_payload_0_184 < _zz_dataOut_payload_0_187);
  assign _zz_dataOut_payload_0_553 = (_zz_dataOut_payload_0_552 ? _zz_dataOut_payload_0_184 : _zz_dataOut_payload_0_187);
  assign _zz_dataOut_payload_0_554 = (_zz_dataOut_payload_0_552 ? _zz_dataOut_payload_0_187 : _zz_dataOut_payload_0_184);
  assign _zz_dataOut_payload_0_555 = (_zz_dataOut_payload_0_185 < _zz_dataOut_payload_0_186);
  assign _zz_dataOut_payload_0_556 = (_zz_dataOut_payload_0_555 ? _zz_dataOut_payload_0_185 : _zz_dataOut_payload_0_186);
  assign _zz_dataOut_payload_0_557 = (_zz_dataOut_payload_0_555 ? _zz_dataOut_payload_0_186 : _zz_dataOut_payload_0_185);
  assign _zz_dataOut_payload_0_558 = (_zz_dataOut_payload_0_553 < _zz_dataOut_payload_0_556);
  assign _zz_dataOut_payload_0_559 = (_zz_dataOut_payload_0_557 < _zz_dataOut_payload_0_554);
  assign _zz_dataOut_payload_0_564 = (_zz_dataOut_payload_0_188 < _zz_dataOut_payload_0_191);
  assign _zz_dataOut_payload_0_565 = (_zz_dataOut_payload_0_564 ? _zz_dataOut_payload_0_188 : _zz_dataOut_payload_0_191);
  assign _zz_dataOut_payload_0_566 = (_zz_dataOut_payload_0_564 ? _zz_dataOut_payload_0_191 : _zz_dataOut_payload_0_188);
  assign _zz_dataOut_payload_0_567 = (_zz_dataOut_payload_0_189 < _zz_dataOut_payload_0_190);
  assign _zz_dataOut_payload_0_568 = (_zz_dataOut_payload_0_567 ? _zz_dataOut_payload_0_189 : _zz_dataOut_payload_0_190);
  assign _zz_dataOut_payload_0_569 = (_zz_dataOut_payload_0_567 ? _zz_dataOut_payload_0_190 : _zz_dataOut_payload_0_189);
  assign _zz_dataOut_payload_0_570 = (_zz_dataOut_payload_0_565 < _zz_dataOut_payload_0_568);
  assign _zz_dataOut_payload_0_571 = (_zz_dataOut_payload_0_569 < _zz_dataOut_payload_0_566);
  assign _zz_dataOut_payload_0_576 = (_zz_dataOut_payload_0_192 < _zz_dataOut_payload_0_195);
  assign _zz_dataOut_payload_0_577 = (_zz_dataOut_payload_0_576 ? _zz_dataOut_payload_0_192 : _zz_dataOut_payload_0_195);
  assign _zz_dataOut_payload_0_578 = (_zz_dataOut_payload_0_576 ? _zz_dataOut_payload_0_195 : _zz_dataOut_payload_0_192);
  assign _zz_dataOut_payload_0_579 = (_zz_dataOut_payload_0_193 < _zz_dataOut_payload_0_194);
  assign _zz_dataOut_payload_0_580 = (_zz_dataOut_payload_0_579 ? _zz_dataOut_payload_0_193 : _zz_dataOut_payload_0_194);
  assign _zz_dataOut_payload_0_581 = (_zz_dataOut_payload_0_579 ? _zz_dataOut_payload_0_194 : _zz_dataOut_payload_0_193);
  assign _zz_dataOut_payload_0_582 = (_zz_dataOut_payload_0_577 < _zz_dataOut_payload_0_580);
  assign _zz_dataOut_payload_0_583 = (_zz_dataOut_payload_0_581 < _zz_dataOut_payload_0_578);
  assign _zz_dataOut_payload_0_588 = (_zz_dataOut_payload_0_196 < _zz_dataOut_payload_0_199);
  assign _zz_dataOut_payload_0_589 = (_zz_dataOut_payload_0_588 ? _zz_dataOut_payload_0_196 : _zz_dataOut_payload_0_199);
  assign _zz_dataOut_payload_0_590 = (_zz_dataOut_payload_0_588 ? _zz_dataOut_payload_0_199 : _zz_dataOut_payload_0_196);
  assign _zz_dataOut_payload_0_591 = (_zz_dataOut_payload_0_197 < _zz_dataOut_payload_0_198);
  assign _zz_dataOut_payload_0_592 = (_zz_dataOut_payload_0_591 ? _zz_dataOut_payload_0_197 : _zz_dataOut_payload_0_198);
  assign _zz_dataOut_payload_0_593 = (_zz_dataOut_payload_0_591 ? _zz_dataOut_payload_0_198 : _zz_dataOut_payload_0_197);
  assign _zz_dataOut_payload_0_594 = (_zz_dataOut_payload_0_589 < _zz_dataOut_payload_0_592);
  assign _zz_dataOut_payload_0_595 = (_zz_dataOut_payload_0_593 < _zz_dataOut_payload_0_590);
  assign _zz_dataOut_payload_0_600 = (_zz_dataOut_payload_0_200 < _zz_dataOut_payload_0_203);
  assign _zz_dataOut_payload_0_601 = (_zz_dataOut_payload_0_600 ? _zz_dataOut_payload_0_200 : _zz_dataOut_payload_0_203);
  assign _zz_dataOut_payload_0_602 = (_zz_dataOut_payload_0_600 ? _zz_dataOut_payload_0_203 : _zz_dataOut_payload_0_200);
  assign _zz_dataOut_payload_0_603 = (_zz_dataOut_payload_0_201 < _zz_dataOut_payload_0_202);
  assign _zz_dataOut_payload_0_604 = (_zz_dataOut_payload_0_603 ? _zz_dataOut_payload_0_201 : _zz_dataOut_payload_0_202);
  assign _zz_dataOut_payload_0_605 = (_zz_dataOut_payload_0_603 ? _zz_dataOut_payload_0_202 : _zz_dataOut_payload_0_201);
  assign _zz_dataOut_payload_0_606 = (_zz_dataOut_payload_0_601 < _zz_dataOut_payload_0_604);
  assign _zz_dataOut_payload_0_607 = (_zz_dataOut_payload_0_605 < _zz_dataOut_payload_0_602);
  assign _zz_dataOut_payload_0_612 = (_zz_dataOut_payload_0_204 < _zz_dataOut_payload_0_207);
  assign _zz_dataOut_payload_0_613 = (_zz_dataOut_payload_0_612 ? _zz_dataOut_payload_0_204 : _zz_dataOut_payload_0_207);
  assign _zz_dataOut_payload_0_614 = (_zz_dataOut_payload_0_612 ? _zz_dataOut_payload_0_207 : _zz_dataOut_payload_0_204);
  assign _zz_dataOut_payload_0_615 = (_zz_dataOut_payload_0_205 < _zz_dataOut_payload_0_206);
  assign _zz_dataOut_payload_0_616 = (_zz_dataOut_payload_0_615 ? _zz_dataOut_payload_0_205 : _zz_dataOut_payload_0_206);
  assign _zz_dataOut_payload_0_617 = (_zz_dataOut_payload_0_615 ? _zz_dataOut_payload_0_206 : _zz_dataOut_payload_0_205);
  assign _zz_dataOut_payload_0_618 = (_zz_dataOut_payload_0_613 < _zz_dataOut_payload_0_616);
  assign _zz_dataOut_payload_0_619 = (_zz_dataOut_payload_0_617 < _zz_dataOut_payload_0_614);
  assign _zz_dataOut_payload_0_624 = (_zz_dataOut_payload_0_208 < _zz_dataOut_payload_0_211);
  assign _zz_dataOut_payload_0_625 = (_zz_dataOut_payload_0_624 ? _zz_dataOut_payload_0_208 : _zz_dataOut_payload_0_211);
  assign _zz_dataOut_payload_0_626 = (_zz_dataOut_payload_0_624 ? _zz_dataOut_payload_0_211 : _zz_dataOut_payload_0_208);
  assign _zz_dataOut_payload_0_627 = (_zz_dataOut_payload_0_209 < _zz_dataOut_payload_0_210);
  assign _zz_dataOut_payload_0_628 = (_zz_dataOut_payload_0_627 ? _zz_dataOut_payload_0_209 : _zz_dataOut_payload_0_210);
  assign _zz_dataOut_payload_0_629 = (_zz_dataOut_payload_0_627 ? _zz_dataOut_payload_0_210 : _zz_dataOut_payload_0_209);
  assign _zz_dataOut_payload_0_630 = (_zz_dataOut_payload_0_625 < _zz_dataOut_payload_0_628);
  assign _zz_dataOut_payload_0_631 = (_zz_dataOut_payload_0_629 < _zz_dataOut_payload_0_626);
  assign _zz_dataOut_payload_0_636 = (_zz_dataOut_payload_0_212 < _zz_dataOut_payload_0_215);
  assign _zz_dataOut_payload_0_637 = (_zz_dataOut_payload_0_636 ? _zz_dataOut_payload_0_212 : _zz_dataOut_payload_0_215);
  assign _zz_dataOut_payload_0_638 = (_zz_dataOut_payload_0_636 ? _zz_dataOut_payload_0_215 : _zz_dataOut_payload_0_212);
  assign _zz_dataOut_payload_0_639 = (_zz_dataOut_payload_0_213 < _zz_dataOut_payload_0_214);
  assign _zz_dataOut_payload_0_640 = (_zz_dataOut_payload_0_639 ? _zz_dataOut_payload_0_213 : _zz_dataOut_payload_0_214);
  assign _zz_dataOut_payload_0_641 = (_zz_dataOut_payload_0_639 ? _zz_dataOut_payload_0_214 : _zz_dataOut_payload_0_213);
  assign _zz_dataOut_payload_0_642 = (_zz_dataOut_payload_0_637 < _zz_dataOut_payload_0_640);
  assign _zz_dataOut_payload_0_643 = (_zz_dataOut_payload_0_641 < _zz_dataOut_payload_0_638);
  assign _zz_dataOut_payload_0_648 = (_zz_dataOut_payload_0_216 < _zz_dataOut_payload_0_219);
  assign _zz_dataOut_payload_0_649 = (_zz_dataOut_payload_0_648 ? _zz_dataOut_payload_0_216 : _zz_dataOut_payload_0_219);
  assign _zz_dataOut_payload_0_650 = (_zz_dataOut_payload_0_648 ? _zz_dataOut_payload_0_219 : _zz_dataOut_payload_0_216);
  assign _zz_dataOut_payload_0_651 = (_zz_dataOut_payload_0_217 < _zz_dataOut_payload_0_218);
  assign _zz_dataOut_payload_0_652 = (_zz_dataOut_payload_0_651 ? _zz_dataOut_payload_0_217 : _zz_dataOut_payload_0_218);
  assign _zz_dataOut_payload_0_653 = (_zz_dataOut_payload_0_651 ? _zz_dataOut_payload_0_218 : _zz_dataOut_payload_0_217);
  assign _zz_dataOut_payload_0_654 = (_zz_dataOut_payload_0_649 < _zz_dataOut_payload_0_652);
  assign _zz_dataOut_payload_0_655 = (_zz_dataOut_payload_0_653 < _zz_dataOut_payload_0_650);
  assign _zz_dataOut_payload_0_660 = (_zz_dataOut_payload_0_220 < _zz_dataOut_payload_0_223);
  assign _zz_dataOut_payload_0_661 = (_zz_dataOut_payload_0_660 ? _zz_dataOut_payload_0_220 : _zz_dataOut_payload_0_223);
  assign _zz_dataOut_payload_0_662 = (_zz_dataOut_payload_0_660 ? _zz_dataOut_payload_0_223 : _zz_dataOut_payload_0_220);
  assign _zz_dataOut_payload_0_663 = (_zz_dataOut_payload_0_221 < _zz_dataOut_payload_0_222);
  assign _zz_dataOut_payload_0_664 = (_zz_dataOut_payload_0_663 ? _zz_dataOut_payload_0_221 : _zz_dataOut_payload_0_222);
  assign _zz_dataOut_payload_0_665 = (_zz_dataOut_payload_0_663 ? _zz_dataOut_payload_0_222 : _zz_dataOut_payload_0_221);
  assign _zz_dataOut_payload_0_666 = (_zz_dataOut_payload_0_661 < _zz_dataOut_payload_0_664);
  assign _zz_dataOut_payload_0_667 = (_zz_dataOut_payload_0_665 < _zz_dataOut_payload_0_662);
  assign _zz_dataOut_payload_0_672 = (_zz_dataOut_payload_0_224 < _zz_dataOut_payload_0_227);
  assign _zz_dataOut_payload_0_673 = (_zz_dataOut_payload_0_672 ? _zz_dataOut_payload_0_224 : _zz_dataOut_payload_0_227);
  assign _zz_dataOut_payload_0_674 = (_zz_dataOut_payload_0_672 ? _zz_dataOut_payload_0_227 : _zz_dataOut_payload_0_224);
  assign _zz_dataOut_payload_0_675 = (_zz_dataOut_payload_0_225 < _zz_dataOut_payload_0_226);
  assign _zz_dataOut_payload_0_676 = (_zz_dataOut_payload_0_675 ? _zz_dataOut_payload_0_225 : _zz_dataOut_payload_0_226);
  assign _zz_dataOut_payload_0_677 = (_zz_dataOut_payload_0_675 ? _zz_dataOut_payload_0_226 : _zz_dataOut_payload_0_225);
  assign _zz_dataOut_payload_0_678 = (_zz_dataOut_payload_0_673 < _zz_dataOut_payload_0_676);
  assign _zz_dataOut_payload_0_679 = (_zz_dataOut_payload_0_677 < _zz_dataOut_payload_0_674);
  assign _zz_dataOut_payload_0_684 = (_zz_dataOut_payload_0_228 < _zz_dataOut_payload_0_231);
  assign _zz_dataOut_payload_0_685 = (_zz_dataOut_payload_0_684 ? _zz_dataOut_payload_0_228 : _zz_dataOut_payload_0_231);
  assign _zz_dataOut_payload_0_686 = (_zz_dataOut_payload_0_684 ? _zz_dataOut_payload_0_231 : _zz_dataOut_payload_0_228);
  assign _zz_dataOut_payload_0_687 = (_zz_dataOut_payload_0_229 < _zz_dataOut_payload_0_230);
  assign _zz_dataOut_payload_0_688 = (_zz_dataOut_payload_0_687 ? _zz_dataOut_payload_0_229 : _zz_dataOut_payload_0_230);
  assign _zz_dataOut_payload_0_689 = (_zz_dataOut_payload_0_687 ? _zz_dataOut_payload_0_230 : _zz_dataOut_payload_0_229);
  assign _zz_dataOut_payload_0_690 = (_zz_dataOut_payload_0_685 < _zz_dataOut_payload_0_688);
  assign _zz_dataOut_payload_0_691 = (_zz_dataOut_payload_0_689 < _zz_dataOut_payload_0_686);
  assign _zz_dataOut_payload_0_696 = (_zz_dataOut_payload_0_232 < _zz_dataOut_payload_0_235);
  assign _zz_dataOut_payload_0_697 = (_zz_dataOut_payload_0_696 ? _zz_dataOut_payload_0_232 : _zz_dataOut_payload_0_235);
  assign _zz_dataOut_payload_0_698 = (_zz_dataOut_payload_0_696 ? _zz_dataOut_payload_0_235 : _zz_dataOut_payload_0_232);
  assign _zz_dataOut_payload_0_699 = (_zz_dataOut_payload_0_233 < _zz_dataOut_payload_0_234);
  assign _zz_dataOut_payload_0_700 = (_zz_dataOut_payload_0_699 ? _zz_dataOut_payload_0_233 : _zz_dataOut_payload_0_234);
  assign _zz_dataOut_payload_0_701 = (_zz_dataOut_payload_0_699 ? _zz_dataOut_payload_0_234 : _zz_dataOut_payload_0_233);
  assign _zz_dataOut_payload_0_702 = (_zz_dataOut_payload_0_697 < _zz_dataOut_payload_0_700);
  assign _zz_dataOut_payload_0_703 = (_zz_dataOut_payload_0_701 < _zz_dataOut_payload_0_698);
  assign _zz_dataOut_payload_0_708 = (_zz_dataOut_payload_0_236 < _zz_dataOut_payload_0_239);
  assign _zz_dataOut_payload_0_709 = (_zz_dataOut_payload_0_708 ? _zz_dataOut_payload_0_236 : _zz_dataOut_payload_0_239);
  assign _zz_dataOut_payload_0_710 = (_zz_dataOut_payload_0_708 ? _zz_dataOut_payload_0_239 : _zz_dataOut_payload_0_236);
  assign _zz_dataOut_payload_0_711 = (_zz_dataOut_payload_0_237 < _zz_dataOut_payload_0_238);
  assign _zz_dataOut_payload_0_712 = (_zz_dataOut_payload_0_711 ? _zz_dataOut_payload_0_237 : _zz_dataOut_payload_0_238);
  assign _zz_dataOut_payload_0_713 = (_zz_dataOut_payload_0_711 ? _zz_dataOut_payload_0_238 : _zz_dataOut_payload_0_237);
  assign _zz_dataOut_payload_0_714 = (_zz_dataOut_payload_0_709 < _zz_dataOut_payload_0_712);
  assign _zz_dataOut_payload_0_715 = (_zz_dataOut_payload_0_713 < _zz_dataOut_payload_0_710);
  assign _zz_dataOut_payload_0_720 = (_zz_dataOut_payload_0_240 < _zz_dataOut_payload_0_243);
  assign _zz_dataOut_payload_0_721 = (_zz_dataOut_payload_0_720 ? _zz_dataOut_payload_0_240 : _zz_dataOut_payload_0_243);
  assign _zz_dataOut_payload_0_722 = (_zz_dataOut_payload_0_720 ? _zz_dataOut_payload_0_243 : _zz_dataOut_payload_0_240);
  assign _zz_dataOut_payload_0_723 = (_zz_dataOut_payload_0_241 < _zz_dataOut_payload_0_242);
  assign _zz_dataOut_payload_0_724 = (_zz_dataOut_payload_0_723 ? _zz_dataOut_payload_0_241 : _zz_dataOut_payload_0_242);
  assign _zz_dataOut_payload_0_725 = (_zz_dataOut_payload_0_723 ? _zz_dataOut_payload_0_242 : _zz_dataOut_payload_0_241);
  assign _zz_dataOut_payload_0_726 = (_zz_dataOut_payload_0_721 < _zz_dataOut_payload_0_724);
  assign _zz_dataOut_payload_0_727 = (_zz_dataOut_payload_0_725 < _zz_dataOut_payload_0_722);
  assign _zz_dataOut_payload_0_732 = (_zz_dataOut_payload_0_244 < _zz_dataOut_payload_0_247);
  assign _zz_dataOut_payload_0_733 = (_zz_dataOut_payload_0_732 ? _zz_dataOut_payload_0_244 : _zz_dataOut_payload_0_247);
  assign _zz_dataOut_payload_0_734 = (_zz_dataOut_payload_0_732 ? _zz_dataOut_payload_0_247 : _zz_dataOut_payload_0_244);
  assign _zz_dataOut_payload_0_735 = (_zz_dataOut_payload_0_245 < _zz_dataOut_payload_0_246);
  assign _zz_dataOut_payload_0_736 = (_zz_dataOut_payload_0_735 ? _zz_dataOut_payload_0_245 : _zz_dataOut_payload_0_246);
  assign _zz_dataOut_payload_0_737 = (_zz_dataOut_payload_0_735 ? _zz_dataOut_payload_0_246 : _zz_dataOut_payload_0_245);
  assign _zz_dataOut_payload_0_738 = (_zz_dataOut_payload_0_733 < _zz_dataOut_payload_0_736);
  assign _zz_dataOut_payload_0_739 = (_zz_dataOut_payload_0_737 < _zz_dataOut_payload_0_734);
  assign _zz_dataOut_payload_0_744 = (_zz_dataOut_payload_0_248 < _zz_dataOut_payload_0_251);
  assign _zz_dataOut_payload_0_745 = (_zz_dataOut_payload_0_744 ? _zz_dataOut_payload_0_248 : _zz_dataOut_payload_0_251);
  assign _zz_dataOut_payload_0_746 = (_zz_dataOut_payload_0_744 ? _zz_dataOut_payload_0_251 : _zz_dataOut_payload_0_248);
  assign _zz_dataOut_payload_0_747 = (_zz_dataOut_payload_0_249 < _zz_dataOut_payload_0_250);
  assign _zz_dataOut_payload_0_748 = (_zz_dataOut_payload_0_747 ? _zz_dataOut_payload_0_249 : _zz_dataOut_payload_0_250);
  assign _zz_dataOut_payload_0_749 = (_zz_dataOut_payload_0_747 ? _zz_dataOut_payload_0_250 : _zz_dataOut_payload_0_249);
  assign _zz_dataOut_payload_0_750 = (_zz_dataOut_payload_0_745 < _zz_dataOut_payload_0_748);
  assign _zz_dataOut_payload_0_751 = (_zz_dataOut_payload_0_749 < _zz_dataOut_payload_0_746);
  assign _zz_dataOut_payload_0_756 = (_zz_dataOut_payload_0_252 < _zz_dataOut_payload_0_255);
  assign _zz_dataOut_payload_0_757 = (_zz_dataOut_payload_0_756 ? _zz_dataOut_payload_0_252 : _zz_dataOut_payload_0_255);
  assign _zz_dataOut_payload_0_758 = (_zz_dataOut_payload_0_756 ? _zz_dataOut_payload_0_255 : _zz_dataOut_payload_0_252);
  assign _zz_dataOut_payload_0_759 = (_zz_dataOut_payload_0_253 < _zz_dataOut_payload_0_254);
  assign _zz_dataOut_payload_0_760 = (_zz_dataOut_payload_0_759 ? _zz_dataOut_payload_0_253 : _zz_dataOut_payload_0_254);
  assign _zz_dataOut_payload_0_761 = (_zz_dataOut_payload_0_759 ? _zz_dataOut_payload_0_254 : _zz_dataOut_payload_0_253);
  assign _zz_dataOut_payload_0_762 = (_zz_dataOut_payload_0_757 < _zz_dataOut_payload_0_760);
  assign _zz_dataOut_payload_0_763 = (_zz_dataOut_payload_0_761 < _zz_dataOut_payload_0_758);
  assign _zz_dataOut_payload_0_768 = (_zz_dataOut_payload_0_256 < _zz_dataOut_payload_0_259);
  assign _zz_dataOut_payload_0_769 = (_zz_dataOut_payload_0_768 ? _zz_dataOut_payload_0_256 : _zz_dataOut_payload_0_259);
  assign _zz_dataOut_payload_0_770 = (_zz_dataOut_payload_0_768 ? _zz_dataOut_payload_0_259 : _zz_dataOut_payload_0_256);
  assign _zz_dataOut_payload_0_771 = (_zz_dataOut_payload_0_257 < _zz_dataOut_payload_0_258);
  assign _zz_dataOut_payload_0_772 = (_zz_dataOut_payload_0_771 ? _zz_dataOut_payload_0_257 : _zz_dataOut_payload_0_258);
  assign _zz_dataOut_payload_0_773 = (_zz_dataOut_payload_0_771 ? _zz_dataOut_payload_0_258 : _zz_dataOut_payload_0_257);
  assign _zz_dataOut_payload_0_774 = (_zz_dataOut_payload_0_769 < _zz_dataOut_payload_0_772);
  assign _zz_dataOut_payload_0_775 = (_zz_dataOut_payload_0_773 < _zz_dataOut_payload_0_770);
  assign _zz_dataOut_payload_0_780 = (_zz_dataOut_payload_0_260 < _zz_dataOut_payload_0_263);
  assign _zz_dataOut_payload_0_781 = (_zz_dataOut_payload_0_780 ? _zz_dataOut_payload_0_260 : _zz_dataOut_payload_0_263);
  assign _zz_dataOut_payload_0_782 = (_zz_dataOut_payload_0_780 ? _zz_dataOut_payload_0_263 : _zz_dataOut_payload_0_260);
  assign _zz_dataOut_payload_0_783 = (_zz_dataOut_payload_0_261 < _zz_dataOut_payload_0_262);
  assign _zz_dataOut_payload_0_784 = (_zz_dataOut_payload_0_783 ? _zz_dataOut_payload_0_261 : _zz_dataOut_payload_0_262);
  assign _zz_dataOut_payload_0_785 = (_zz_dataOut_payload_0_783 ? _zz_dataOut_payload_0_262 : _zz_dataOut_payload_0_261);
  assign _zz_dataOut_payload_0_786 = (_zz_dataOut_payload_0_781 < _zz_dataOut_payload_0_784);
  assign _zz_dataOut_payload_0_787 = (_zz_dataOut_payload_0_785 < _zz_dataOut_payload_0_782);
  assign _zz_dataOut_payload_0_792 = (_zz_dataOut_payload_0_264 < _zz_dataOut_payload_0_267);
  assign _zz_dataOut_payload_0_793 = (_zz_dataOut_payload_0_792 ? _zz_dataOut_payload_0_264 : _zz_dataOut_payload_0_267);
  assign _zz_dataOut_payload_0_794 = (_zz_dataOut_payload_0_792 ? _zz_dataOut_payload_0_267 : _zz_dataOut_payload_0_264);
  assign _zz_dataOut_payload_0_795 = (_zz_dataOut_payload_0_265 < _zz_dataOut_payload_0_266);
  assign _zz_dataOut_payload_0_796 = (_zz_dataOut_payload_0_795 ? _zz_dataOut_payload_0_265 : _zz_dataOut_payload_0_266);
  assign _zz_dataOut_payload_0_797 = (_zz_dataOut_payload_0_795 ? _zz_dataOut_payload_0_266 : _zz_dataOut_payload_0_265);
  assign _zz_dataOut_payload_0_798 = (_zz_dataOut_payload_0_793 < _zz_dataOut_payload_0_796);
  assign _zz_dataOut_payload_0_799 = (_zz_dataOut_payload_0_797 < _zz_dataOut_payload_0_794);
  assign _zz_dataOut_payload_0_804 = (_zz_dataOut_payload_0_268 < _zz_dataOut_payload_0_271);
  assign _zz_dataOut_payload_0_805 = (_zz_dataOut_payload_0_804 ? _zz_dataOut_payload_0_268 : _zz_dataOut_payload_0_271);
  assign _zz_dataOut_payload_0_806 = (_zz_dataOut_payload_0_804 ? _zz_dataOut_payload_0_271 : _zz_dataOut_payload_0_268);
  assign _zz_dataOut_payload_0_807 = (_zz_dataOut_payload_0_269 < _zz_dataOut_payload_0_270);
  assign _zz_dataOut_payload_0_808 = (_zz_dataOut_payload_0_807 ? _zz_dataOut_payload_0_269 : _zz_dataOut_payload_0_270);
  assign _zz_dataOut_payload_0_809 = (_zz_dataOut_payload_0_807 ? _zz_dataOut_payload_0_270 : _zz_dataOut_payload_0_269);
  assign _zz_dataOut_payload_0_810 = (_zz_dataOut_payload_0_805 < _zz_dataOut_payload_0_808);
  assign _zz_dataOut_payload_0_811 = (_zz_dataOut_payload_0_809 < _zz_dataOut_payload_0_806);
  assign _zz_dataOut_payload_0_816 = (_zz_dataOut_payload_0_272 < _zz_dataOut_payload_0_275);
  assign _zz_dataOut_payload_0_817 = (_zz_dataOut_payload_0_816 ? _zz_dataOut_payload_0_272 : _zz_dataOut_payload_0_275);
  assign _zz_dataOut_payload_0_818 = (_zz_dataOut_payload_0_816 ? _zz_dataOut_payload_0_275 : _zz_dataOut_payload_0_272);
  assign _zz_dataOut_payload_0_819 = (_zz_dataOut_payload_0_273 < _zz_dataOut_payload_0_274);
  assign _zz_dataOut_payload_0_820 = (_zz_dataOut_payload_0_819 ? _zz_dataOut_payload_0_273 : _zz_dataOut_payload_0_274);
  assign _zz_dataOut_payload_0_821 = (_zz_dataOut_payload_0_819 ? _zz_dataOut_payload_0_274 : _zz_dataOut_payload_0_273);
  assign _zz_dataOut_payload_0_822 = (_zz_dataOut_payload_0_817 < _zz_dataOut_payload_0_820);
  assign _zz_dataOut_payload_0_823 = (_zz_dataOut_payload_0_821 < _zz_dataOut_payload_0_818);
  assign _zz_dataOut_payload_0_828 = (_zz_dataOut_payload_0_276 < _zz_dataOut_payload_0_279);
  assign _zz_dataOut_payload_0_829 = (_zz_dataOut_payload_0_828 ? _zz_dataOut_payload_0_276 : _zz_dataOut_payload_0_279);
  assign _zz_dataOut_payload_0_830 = (_zz_dataOut_payload_0_828 ? _zz_dataOut_payload_0_279 : _zz_dataOut_payload_0_276);
  assign _zz_dataOut_payload_0_831 = (_zz_dataOut_payload_0_277 < _zz_dataOut_payload_0_278);
  assign _zz_dataOut_payload_0_832 = (_zz_dataOut_payload_0_831 ? _zz_dataOut_payload_0_277 : _zz_dataOut_payload_0_278);
  assign _zz_dataOut_payload_0_833 = (_zz_dataOut_payload_0_831 ? _zz_dataOut_payload_0_278 : _zz_dataOut_payload_0_277);
  assign _zz_dataOut_payload_0_834 = (_zz_dataOut_payload_0_829 < _zz_dataOut_payload_0_832);
  assign _zz_dataOut_payload_0_835 = (_zz_dataOut_payload_0_833 < _zz_dataOut_payload_0_830);
  assign _zz_dataOut_payload_0_840 = (_zz_dataOut_payload_0_280 < _zz_dataOut_payload_0_283);
  assign _zz_dataOut_payload_0_841 = (_zz_dataOut_payload_0_840 ? _zz_dataOut_payload_0_280 : _zz_dataOut_payload_0_283);
  assign _zz_dataOut_payload_0_842 = (_zz_dataOut_payload_0_840 ? _zz_dataOut_payload_0_283 : _zz_dataOut_payload_0_280);
  assign _zz_dataOut_payload_0_843 = (_zz_dataOut_payload_0_281 < _zz_dataOut_payload_0_282);
  assign _zz_dataOut_payload_0_844 = (_zz_dataOut_payload_0_843 ? _zz_dataOut_payload_0_281 : _zz_dataOut_payload_0_282);
  assign _zz_dataOut_payload_0_845 = (_zz_dataOut_payload_0_843 ? _zz_dataOut_payload_0_282 : _zz_dataOut_payload_0_281);
  assign _zz_dataOut_payload_0_846 = (_zz_dataOut_payload_0_841 < _zz_dataOut_payload_0_844);
  assign _zz_dataOut_payload_0_847 = (_zz_dataOut_payload_0_845 < _zz_dataOut_payload_0_842);
  assign _zz_dataOut_payload_0_852 = (_zz_dataOut_payload_0_284 < _zz_dataOut_payload_0_287);
  assign _zz_dataOut_payload_0_853 = (_zz_dataOut_payload_0_852 ? _zz_dataOut_payload_0_284 : _zz_dataOut_payload_0_287);
  assign _zz_dataOut_payload_0_854 = (_zz_dataOut_payload_0_852 ? _zz_dataOut_payload_0_287 : _zz_dataOut_payload_0_284);
  assign _zz_dataOut_payload_0_855 = (_zz_dataOut_payload_0_285 < _zz_dataOut_payload_0_286);
  assign _zz_dataOut_payload_0_856 = (_zz_dataOut_payload_0_855 ? _zz_dataOut_payload_0_285 : _zz_dataOut_payload_0_286);
  assign _zz_dataOut_payload_0_857 = (_zz_dataOut_payload_0_855 ? _zz_dataOut_payload_0_286 : _zz_dataOut_payload_0_285);
  assign _zz_dataOut_payload_0_858 = (_zz_dataOut_payload_0_853 < _zz_dataOut_payload_0_856);
  assign _zz_dataOut_payload_0_859 = (_zz_dataOut_payload_0_857 < _zz_dataOut_payload_0_854);
  assign _zz_dataOut_payload_0_864 = (_zz_dataOut_payload_0_288 < _zz_dataOut_payload_0_291);
  assign _zz_dataOut_payload_0_865 = (_zz_dataOut_payload_0_864 ? _zz_dataOut_payload_0_288 : _zz_dataOut_payload_0_291);
  assign _zz_dataOut_payload_0_866 = (_zz_dataOut_payload_0_864 ? _zz_dataOut_payload_0_291 : _zz_dataOut_payload_0_288);
  assign _zz_dataOut_payload_0_867 = (_zz_dataOut_payload_0_289 < _zz_dataOut_payload_0_290);
  assign _zz_dataOut_payload_0_868 = (_zz_dataOut_payload_0_867 ? _zz_dataOut_payload_0_289 : _zz_dataOut_payload_0_290);
  assign _zz_dataOut_payload_0_869 = (_zz_dataOut_payload_0_867 ? _zz_dataOut_payload_0_290 : _zz_dataOut_payload_0_289);
  assign _zz_dataOut_payload_0_870 = (_zz_dataOut_payload_0_865 < _zz_dataOut_payload_0_868);
  assign _zz_dataOut_payload_0_871 = (_zz_dataOut_payload_0_869 < _zz_dataOut_payload_0_866);
  assign _zz_dataOut_payload_0_876 = (_zz_dataOut_payload_0_292 < _zz_dataOut_payload_0_295);
  assign _zz_dataOut_payload_0_877 = (_zz_dataOut_payload_0_876 ? _zz_dataOut_payload_0_292 : _zz_dataOut_payload_0_295);
  assign _zz_dataOut_payload_0_878 = (_zz_dataOut_payload_0_876 ? _zz_dataOut_payload_0_295 : _zz_dataOut_payload_0_292);
  assign _zz_dataOut_payload_0_879 = (_zz_dataOut_payload_0_293 < _zz_dataOut_payload_0_294);
  assign _zz_dataOut_payload_0_880 = (_zz_dataOut_payload_0_879 ? _zz_dataOut_payload_0_293 : _zz_dataOut_payload_0_294);
  assign _zz_dataOut_payload_0_881 = (_zz_dataOut_payload_0_879 ? _zz_dataOut_payload_0_294 : _zz_dataOut_payload_0_293);
  assign _zz_dataOut_payload_0_882 = (_zz_dataOut_payload_0_877 < _zz_dataOut_payload_0_880);
  assign _zz_dataOut_payload_0_883 = (_zz_dataOut_payload_0_881 < _zz_dataOut_payload_0_878);
  assign _zz_dataOut_payload_0_888 = (_zz_dataOut_payload_0_296 < _zz_dataOut_payload_0_299);
  assign _zz_dataOut_payload_0_889 = (_zz_dataOut_payload_0_888 ? _zz_dataOut_payload_0_296 : _zz_dataOut_payload_0_299);
  assign _zz_dataOut_payload_0_890 = (_zz_dataOut_payload_0_888 ? _zz_dataOut_payload_0_299 : _zz_dataOut_payload_0_296);
  assign _zz_dataOut_payload_0_891 = (_zz_dataOut_payload_0_297 < _zz_dataOut_payload_0_298);
  assign _zz_dataOut_payload_0_892 = (_zz_dataOut_payload_0_891 ? _zz_dataOut_payload_0_297 : _zz_dataOut_payload_0_298);
  assign _zz_dataOut_payload_0_893 = (_zz_dataOut_payload_0_891 ? _zz_dataOut_payload_0_298 : _zz_dataOut_payload_0_297);
  assign _zz_dataOut_payload_0_894 = (_zz_dataOut_payload_0_889 < _zz_dataOut_payload_0_892);
  assign _zz_dataOut_payload_0_895 = (_zz_dataOut_payload_0_893 < _zz_dataOut_payload_0_890);
  assign _zz_dataOut_payload_0_900 = (_zz_dataOut_payload_0_300 < _zz_dataOut_payload_0_303);
  assign _zz_dataOut_payload_0_901 = (_zz_dataOut_payload_0_900 ? _zz_dataOut_payload_0_300 : _zz_dataOut_payload_0_303);
  assign _zz_dataOut_payload_0_902 = (_zz_dataOut_payload_0_900 ? _zz_dataOut_payload_0_303 : _zz_dataOut_payload_0_300);
  assign _zz_dataOut_payload_0_903 = (_zz_dataOut_payload_0_301 < _zz_dataOut_payload_0_302);
  assign _zz_dataOut_payload_0_904 = (_zz_dataOut_payload_0_903 ? _zz_dataOut_payload_0_301 : _zz_dataOut_payload_0_302);
  assign _zz_dataOut_payload_0_905 = (_zz_dataOut_payload_0_903 ? _zz_dataOut_payload_0_302 : _zz_dataOut_payload_0_301);
  assign _zz_dataOut_payload_0_906 = (_zz_dataOut_payload_0_901 < _zz_dataOut_payload_0_904);
  assign _zz_dataOut_payload_0_907 = (_zz_dataOut_payload_0_905 < _zz_dataOut_payload_0_902);
  assign _zz_dataOut_payload_0_912 = (_zz_dataOut_payload_0_304 < _zz_dataOut_payload_0_307);
  assign _zz_dataOut_payload_0_913 = (_zz_dataOut_payload_0_912 ? _zz_dataOut_payload_0_304 : _zz_dataOut_payload_0_307);
  assign _zz_dataOut_payload_0_914 = (_zz_dataOut_payload_0_912 ? _zz_dataOut_payload_0_307 : _zz_dataOut_payload_0_304);
  assign _zz_dataOut_payload_0_915 = (_zz_dataOut_payload_0_305 < _zz_dataOut_payload_0_306);
  assign _zz_dataOut_payload_0_916 = (_zz_dataOut_payload_0_915 ? _zz_dataOut_payload_0_305 : _zz_dataOut_payload_0_306);
  assign _zz_dataOut_payload_0_917 = (_zz_dataOut_payload_0_915 ? _zz_dataOut_payload_0_306 : _zz_dataOut_payload_0_305);
  assign _zz_dataOut_payload_0_918 = (_zz_dataOut_payload_0_913 < _zz_dataOut_payload_0_916);
  assign _zz_dataOut_payload_0_919 = (_zz_dataOut_payload_0_917 < _zz_dataOut_payload_0_914);
  assign _zz_dataOut_payload_0_924 = (_zz_dataOut_payload_0_308 < _zz_dataOut_payload_0_311);
  assign _zz_dataOut_payload_0_925 = (_zz_dataOut_payload_0_924 ? _zz_dataOut_payload_0_308 : _zz_dataOut_payload_0_311);
  assign _zz_dataOut_payload_0_926 = (_zz_dataOut_payload_0_924 ? _zz_dataOut_payload_0_311 : _zz_dataOut_payload_0_308);
  assign _zz_dataOut_payload_0_927 = (_zz_dataOut_payload_0_309 < _zz_dataOut_payload_0_310);
  assign _zz_dataOut_payload_0_928 = (_zz_dataOut_payload_0_927 ? _zz_dataOut_payload_0_309 : _zz_dataOut_payload_0_310);
  assign _zz_dataOut_payload_0_929 = (_zz_dataOut_payload_0_927 ? _zz_dataOut_payload_0_310 : _zz_dataOut_payload_0_309);
  assign _zz_dataOut_payload_0_930 = (_zz_dataOut_payload_0_925 < _zz_dataOut_payload_0_928);
  assign _zz_dataOut_payload_0_931 = (_zz_dataOut_payload_0_929 < _zz_dataOut_payload_0_926);
  assign _zz_dataOut_payload_0_936 = (_zz_dataOut_payload_0_312 < _zz_dataOut_payload_0_315);
  assign _zz_dataOut_payload_0_937 = (_zz_dataOut_payload_0_936 ? _zz_dataOut_payload_0_312 : _zz_dataOut_payload_0_315);
  assign _zz_dataOut_payload_0_938 = (_zz_dataOut_payload_0_936 ? _zz_dataOut_payload_0_315 : _zz_dataOut_payload_0_312);
  assign _zz_dataOut_payload_0_939 = (_zz_dataOut_payload_0_313 < _zz_dataOut_payload_0_314);
  assign _zz_dataOut_payload_0_940 = (_zz_dataOut_payload_0_939 ? _zz_dataOut_payload_0_313 : _zz_dataOut_payload_0_314);
  assign _zz_dataOut_payload_0_941 = (_zz_dataOut_payload_0_939 ? _zz_dataOut_payload_0_314 : _zz_dataOut_payload_0_313);
  assign _zz_dataOut_payload_0_942 = (_zz_dataOut_payload_0_937 < _zz_dataOut_payload_0_940);
  assign _zz_dataOut_payload_0_943 = (_zz_dataOut_payload_0_941 < _zz_dataOut_payload_0_938);
  assign _zz_dataOut_payload_0_948 = (_zz_dataOut_payload_0_316 < _zz_dataOut_payload_0_319);
  assign _zz_dataOut_payload_0_949 = (_zz_dataOut_payload_0_948 ? _zz_dataOut_payload_0_316 : _zz_dataOut_payload_0_319);
  assign _zz_dataOut_payload_0_950 = (_zz_dataOut_payload_0_948 ? _zz_dataOut_payload_0_319 : _zz_dataOut_payload_0_316);
  assign _zz_dataOut_payload_0_951 = (_zz_dataOut_payload_0_317 < _zz_dataOut_payload_0_318);
  assign _zz_dataOut_payload_0_952 = (_zz_dataOut_payload_0_951 ? _zz_dataOut_payload_0_317 : _zz_dataOut_payload_0_318);
  assign _zz_dataOut_payload_0_953 = (_zz_dataOut_payload_0_951 ? _zz_dataOut_payload_0_318 : _zz_dataOut_payload_0_317);
  assign _zz_dataOut_payload_0_954 = (_zz_dataOut_payload_0_949 < _zz_dataOut_payload_0_952);
  assign _zz_dataOut_payload_0_955 = (_zz_dataOut_payload_0_953 < _zz_dataOut_payload_0_950);
  assign _zz_dataOut_payload_0_960 = (_zz_dataOut_payload_0_320 < _zz_dataOut_payload_0_323);
  assign _zz_dataOut_payload_0_961 = (_zz_dataOut_payload_0_960 ? _zz_dataOut_payload_0_320 : _zz_dataOut_payload_0_323);
  assign _zz_dataOut_payload_0_962 = (_zz_dataOut_payload_0_960 ? _zz_dataOut_payload_0_323 : _zz_dataOut_payload_0_320);
  assign _zz_dataOut_payload_0_963 = (_zz_dataOut_payload_0_321 < _zz_dataOut_payload_0_322);
  assign _zz_dataOut_payload_0_964 = (_zz_dataOut_payload_0_963 ? _zz_dataOut_payload_0_321 : _zz_dataOut_payload_0_322);
  assign _zz_dataOut_payload_0_965 = (_zz_dataOut_payload_0_963 ? _zz_dataOut_payload_0_322 : _zz_dataOut_payload_0_321);
  assign _zz_dataOut_payload_0_966 = (_zz_dataOut_payload_0_961 < _zz_dataOut_payload_0_964);
  assign _zz_dataOut_payload_0_967 = (_zz_dataOut_payload_0_965 < _zz_dataOut_payload_0_962);
  assign _zz_dataOut_payload_0_972 = (_zz_dataOut_payload_0_324 < _zz_dataOut_payload_0_327);
  assign _zz_dataOut_payload_0_973 = (_zz_dataOut_payload_0_972 ? _zz_dataOut_payload_0_324 : _zz_dataOut_payload_0_327);
  assign _zz_dataOut_payload_0_974 = (_zz_dataOut_payload_0_972 ? _zz_dataOut_payload_0_327 : _zz_dataOut_payload_0_324);
  assign _zz_dataOut_payload_0_975 = (_zz_dataOut_payload_0_325 < _zz_dataOut_payload_0_326);
  assign _zz_dataOut_payload_0_976 = (_zz_dataOut_payload_0_975 ? _zz_dataOut_payload_0_325 : _zz_dataOut_payload_0_326);
  assign _zz_dataOut_payload_0_977 = (_zz_dataOut_payload_0_975 ? _zz_dataOut_payload_0_326 : _zz_dataOut_payload_0_325);
  assign _zz_dataOut_payload_0_978 = (_zz_dataOut_payload_0_973 < _zz_dataOut_payload_0_976);
  assign _zz_dataOut_payload_0_979 = (_zz_dataOut_payload_0_977 < _zz_dataOut_payload_0_974);
  assign _zz_dataOut_payload_0_984 = (_zz_dataOut_payload_0_328 < _zz_dataOut_payload_0_331);
  assign _zz_dataOut_payload_0_985 = (_zz_dataOut_payload_0_984 ? _zz_dataOut_payload_0_328 : _zz_dataOut_payload_0_331);
  assign _zz_dataOut_payload_0_986 = (_zz_dataOut_payload_0_984 ? _zz_dataOut_payload_0_331 : _zz_dataOut_payload_0_328);
  assign _zz_dataOut_payload_0_987 = (_zz_dataOut_payload_0_329 < _zz_dataOut_payload_0_330);
  assign _zz_dataOut_payload_0_988 = (_zz_dataOut_payload_0_987 ? _zz_dataOut_payload_0_329 : _zz_dataOut_payload_0_330);
  assign _zz_dataOut_payload_0_989 = (_zz_dataOut_payload_0_987 ? _zz_dataOut_payload_0_330 : _zz_dataOut_payload_0_329);
  assign _zz_dataOut_payload_0_990 = (_zz_dataOut_payload_0_985 < _zz_dataOut_payload_0_988);
  assign _zz_dataOut_payload_0_991 = (_zz_dataOut_payload_0_989 < _zz_dataOut_payload_0_986);
  assign _zz_dataOut_payload_0_996 = (_zz_dataOut_payload_0_332 < _zz_dataOut_payload_0_335);
  assign _zz_dataOut_payload_0_997 = (_zz_dataOut_payload_0_996 ? _zz_dataOut_payload_0_332 : _zz_dataOut_payload_0_335);
  assign _zz_dataOut_payload_0_998 = (_zz_dataOut_payload_0_996 ? _zz_dataOut_payload_0_335 : _zz_dataOut_payload_0_332);
  assign _zz_dataOut_payload_0_999 = (_zz_dataOut_payload_0_333 < _zz_dataOut_payload_0_334);
  assign _zz_dataOut_payload_0_1000 = (_zz_dataOut_payload_0_999 ? _zz_dataOut_payload_0_333 : _zz_dataOut_payload_0_334);
  assign _zz_dataOut_payload_0_1001 = (_zz_dataOut_payload_0_999 ? _zz_dataOut_payload_0_334 : _zz_dataOut_payload_0_333);
  assign _zz_dataOut_payload_0_1002 = (_zz_dataOut_payload_0_997 < _zz_dataOut_payload_0_1000);
  assign _zz_dataOut_payload_0_1003 = (_zz_dataOut_payload_0_1001 < _zz_dataOut_payload_0_998);
  assign _zz_dataOut_payload_0_1008 = (_zz_dataOut_payload_0_336 < _zz_dataOut_payload_0_339);
  assign _zz_dataOut_payload_0_1009 = (_zz_dataOut_payload_0_1008 ? _zz_dataOut_payload_0_336 : _zz_dataOut_payload_0_339);
  assign _zz_dataOut_payload_0_1010 = (_zz_dataOut_payload_0_1008 ? _zz_dataOut_payload_0_339 : _zz_dataOut_payload_0_336);
  assign _zz_dataOut_payload_0_1011 = (_zz_dataOut_payload_0_337 < _zz_dataOut_payload_0_338);
  assign _zz_dataOut_payload_0_1012 = (_zz_dataOut_payload_0_1011 ? _zz_dataOut_payload_0_337 : _zz_dataOut_payload_0_338);
  assign _zz_dataOut_payload_0_1013 = (_zz_dataOut_payload_0_1011 ? _zz_dataOut_payload_0_338 : _zz_dataOut_payload_0_337);
  assign _zz_dataOut_payload_0_1014 = (_zz_dataOut_payload_0_1009 < _zz_dataOut_payload_0_1012);
  assign _zz_dataOut_payload_0_1015 = (_zz_dataOut_payload_0_1013 < _zz_dataOut_payload_0_1010);
  assign _zz_dataOut_payload_0_1020 = (_zz_dataOut_payload_0_340 < _zz_dataOut_payload_0_343);
  assign _zz_dataOut_payload_0_1021 = (_zz_dataOut_payload_0_1020 ? _zz_dataOut_payload_0_340 : _zz_dataOut_payload_0_343);
  assign _zz_dataOut_payload_0_1022 = (_zz_dataOut_payload_0_1020 ? _zz_dataOut_payload_0_343 : _zz_dataOut_payload_0_340);
  assign _zz_dataOut_payload_0_1023 = (_zz_dataOut_payload_0_341 < _zz_dataOut_payload_0_342);
  assign _zz_dataOut_payload_0_1024 = (_zz_dataOut_payload_0_1023 ? _zz_dataOut_payload_0_341 : _zz_dataOut_payload_0_342);
  assign _zz_dataOut_payload_0_1025 = (_zz_dataOut_payload_0_1023 ? _zz_dataOut_payload_0_342 : _zz_dataOut_payload_0_341);
  assign _zz_dataOut_payload_0_1026 = (_zz_dataOut_payload_0_1021 < _zz_dataOut_payload_0_1024);
  assign _zz_dataOut_payload_0_1027 = (_zz_dataOut_payload_0_1025 < _zz_dataOut_payload_0_1022);
  assign _zz_dataOut_payload_0_1032 = (_zz_dataOut_payload_0_344 < _zz_dataOut_payload_0_347);
  assign _zz_dataOut_payload_0_1033 = (_zz_dataOut_payload_0_1032 ? _zz_dataOut_payload_0_344 : _zz_dataOut_payload_0_347);
  assign _zz_dataOut_payload_0_1034 = (_zz_dataOut_payload_0_1032 ? _zz_dataOut_payload_0_347 : _zz_dataOut_payload_0_344);
  assign _zz_dataOut_payload_0_1035 = (_zz_dataOut_payload_0_345 < _zz_dataOut_payload_0_346);
  assign _zz_dataOut_payload_0_1036 = (_zz_dataOut_payload_0_1035 ? _zz_dataOut_payload_0_345 : _zz_dataOut_payload_0_346);
  assign _zz_dataOut_payload_0_1037 = (_zz_dataOut_payload_0_1035 ? _zz_dataOut_payload_0_346 : _zz_dataOut_payload_0_345);
  assign _zz_dataOut_payload_0_1038 = (_zz_dataOut_payload_0_1033 < _zz_dataOut_payload_0_1036);
  assign _zz_dataOut_payload_0_1039 = (_zz_dataOut_payload_0_1037 < _zz_dataOut_payload_0_1034);
  assign _zz_dataOut_payload_0_1044 = (_zz_dataOut_payload_0_348 < _zz_dataOut_payload_0_351);
  assign _zz_dataOut_payload_0_1045 = (_zz_dataOut_payload_0_1044 ? _zz_dataOut_payload_0_348 : _zz_dataOut_payload_0_351);
  assign _zz_dataOut_payload_0_1046 = (_zz_dataOut_payload_0_1044 ? _zz_dataOut_payload_0_351 : _zz_dataOut_payload_0_348);
  assign _zz_dataOut_payload_0_1047 = (_zz_dataOut_payload_0_349 < _zz_dataOut_payload_0_350);
  assign _zz_dataOut_payload_0_1048 = (_zz_dataOut_payload_0_1047 ? _zz_dataOut_payload_0_349 : _zz_dataOut_payload_0_350);
  assign _zz_dataOut_payload_0_1049 = (_zz_dataOut_payload_0_1047 ? _zz_dataOut_payload_0_350 : _zz_dataOut_payload_0_349);
  assign _zz_dataOut_payload_0_1050 = (_zz_dataOut_payload_0_1045 < _zz_dataOut_payload_0_1048);
  assign _zz_dataOut_payload_0_1051 = (_zz_dataOut_payload_0_1049 < _zz_dataOut_payload_0_1046);
  assign _zz_dataOut_payload_0_1056 = (_zz_dataOut_payload_0_352 < _zz_dataOut_payload_0_355);
  assign _zz_dataOut_payload_0_1057 = (_zz_dataOut_payload_0_1056 ? _zz_dataOut_payload_0_352 : _zz_dataOut_payload_0_355);
  assign _zz_dataOut_payload_0_1058 = (_zz_dataOut_payload_0_1056 ? _zz_dataOut_payload_0_355 : _zz_dataOut_payload_0_352);
  assign _zz_dataOut_payload_0_1059 = (_zz_dataOut_payload_0_353 < _zz_dataOut_payload_0_354);
  assign _zz_dataOut_payload_0_1060 = (_zz_dataOut_payload_0_1059 ? _zz_dataOut_payload_0_353 : _zz_dataOut_payload_0_354);
  assign _zz_dataOut_payload_0_1061 = (_zz_dataOut_payload_0_1059 ? _zz_dataOut_payload_0_354 : _zz_dataOut_payload_0_353);
  assign _zz_dataOut_payload_0_1062 = (_zz_dataOut_payload_0_1057 < _zz_dataOut_payload_0_1060);
  assign _zz_dataOut_payload_0_1063 = (_zz_dataOut_payload_0_1061 < _zz_dataOut_payload_0_1058);
  assign _zz_dataOut_payload_0_1068 = (_zz_dataOut_payload_0_356 < _zz_dataOut_payload_0_359);
  assign _zz_dataOut_payload_0_1069 = (_zz_dataOut_payload_0_1068 ? _zz_dataOut_payload_0_356 : _zz_dataOut_payload_0_359);
  assign _zz_dataOut_payload_0_1070 = (_zz_dataOut_payload_0_1068 ? _zz_dataOut_payload_0_359 : _zz_dataOut_payload_0_356);
  assign _zz_dataOut_payload_0_1071 = (_zz_dataOut_payload_0_357 < _zz_dataOut_payload_0_358);
  assign _zz_dataOut_payload_0_1072 = (_zz_dataOut_payload_0_1071 ? _zz_dataOut_payload_0_357 : _zz_dataOut_payload_0_358);
  assign _zz_dataOut_payload_0_1073 = (_zz_dataOut_payload_0_1071 ? _zz_dataOut_payload_0_358 : _zz_dataOut_payload_0_357);
  assign _zz_dataOut_payload_0_1074 = (_zz_dataOut_payload_0_1069 < _zz_dataOut_payload_0_1072);
  assign _zz_dataOut_payload_0_1075 = (_zz_dataOut_payload_0_1073 < _zz_dataOut_payload_0_1070);
  assign _zz_dataOut_payload_0_1080 = (_zz_dataOut_payload_0_360 < _zz_dataOut_payload_0_363);
  assign _zz_dataOut_payload_0_1081 = (_zz_dataOut_payload_0_1080 ? _zz_dataOut_payload_0_360 : _zz_dataOut_payload_0_363);
  assign _zz_dataOut_payload_0_1082 = (_zz_dataOut_payload_0_1080 ? _zz_dataOut_payload_0_363 : _zz_dataOut_payload_0_360);
  assign _zz_dataOut_payload_0_1083 = (_zz_dataOut_payload_0_361 < _zz_dataOut_payload_0_362);
  assign _zz_dataOut_payload_0_1084 = (_zz_dataOut_payload_0_1083 ? _zz_dataOut_payload_0_361 : _zz_dataOut_payload_0_362);
  assign _zz_dataOut_payload_0_1085 = (_zz_dataOut_payload_0_1083 ? _zz_dataOut_payload_0_362 : _zz_dataOut_payload_0_361);
  assign _zz_dataOut_payload_0_1086 = (_zz_dataOut_payload_0_1081 < _zz_dataOut_payload_0_1084);
  assign _zz_dataOut_payload_0_1087 = (_zz_dataOut_payload_0_1085 < _zz_dataOut_payload_0_1082);
  assign _zz_dataOut_payload_0_1092 = (_zz_dataOut_payload_0_364 < _zz_dataOut_payload_0_367);
  assign _zz_dataOut_payload_0_1093 = (_zz_dataOut_payload_0_1092 ? _zz_dataOut_payload_0_364 : _zz_dataOut_payload_0_367);
  assign _zz_dataOut_payload_0_1094 = (_zz_dataOut_payload_0_1092 ? _zz_dataOut_payload_0_367 : _zz_dataOut_payload_0_364);
  assign _zz_dataOut_payload_0_1095 = (_zz_dataOut_payload_0_365 < _zz_dataOut_payload_0_366);
  assign _zz_dataOut_payload_0_1096 = (_zz_dataOut_payload_0_1095 ? _zz_dataOut_payload_0_365 : _zz_dataOut_payload_0_366);
  assign _zz_dataOut_payload_0_1097 = (_zz_dataOut_payload_0_1095 ? _zz_dataOut_payload_0_366 : _zz_dataOut_payload_0_365);
  assign _zz_dataOut_payload_0_1098 = (_zz_dataOut_payload_0_1093 < _zz_dataOut_payload_0_1096);
  assign _zz_dataOut_payload_0_1099 = (_zz_dataOut_payload_0_1097 < _zz_dataOut_payload_0_1094);
  assign _zz_dataOut_payload_0_1104 = (_zz_dataOut_payload_0_368 < _zz_dataOut_payload_0_371);
  assign _zz_dataOut_payload_0_1105 = (_zz_dataOut_payload_0_1104 ? _zz_dataOut_payload_0_368 : _zz_dataOut_payload_0_371);
  assign _zz_dataOut_payload_0_1106 = (_zz_dataOut_payload_0_1104 ? _zz_dataOut_payload_0_371 : _zz_dataOut_payload_0_368);
  assign _zz_dataOut_payload_0_1107 = (_zz_dataOut_payload_0_369 < _zz_dataOut_payload_0_370);
  assign _zz_dataOut_payload_0_1108 = (_zz_dataOut_payload_0_1107 ? _zz_dataOut_payload_0_369 : _zz_dataOut_payload_0_370);
  assign _zz_dataOut_payload_0_1109 = (_zz_dataOut_payload_0_1107 ? _zz_dataOut_payload_0_370 : _zz_dataOut_payload_0_369);
  assign _zz_dataOut_payload_0_1110 = (_zz_dataOut_payload_0_1105 < _zz_dataOut_payload_0_1108);
  assign _zz_dataOut_payload_0_1111 = (_zz_dataOut_payload_0_1109 < _zz_dataOut_payload_0_1106);
  assign _zz_dataOut_payload_0_1116 = (_zz_dataOut_payload_0_372 < _zz_dataOut_payload_0_375);
  assign _zz_dataOut_payload_0_1117 = (_zz_dataOut_payload_0_1116 ? _zz_dataOut_payload_0_372 : _zz_dataOut_payload_0_375);
  assign _zz_dataOut_payload_0_1118 = (_zz_dataOut_payload_0_1116 ? _zz_dataOut_payload_0_375 : _zz_dataOut_payload_0_372);
  assign _zz_dataOut_payload_0_1119 = (_zz_dataOut_payload_0_373 < _zz_dataOut_payload_0_374);
  assign _zz_dataOut_payload_0_1120 = (_zz_dataOut_payload_0_1119 ? _zz_dataOut_payload_0_373 : _zz_dataOut_payload_0_374);
  assign _zz_dataOut_payload_0_1121 = (_zz_dataOut_payload_0_1119 ? _zz_dataOut_payload_0_374 : _zz_dataOut_payload_0_373);
  assign _zz_dataOut_payload_0_1122 = (_zz_dataOut_payload_0_1117 < _zz_dataOut_payload_0_1120);
  assign _zz_dataOut_payload_0_1123 = (_zz_dataOut_payload_0_1121 < _zz_dataOut_payload_0_1118);
  assign _zz_dataOut_payload_0_1128 = (_zz_dataOut_payload_0_376 < _zz_dataOut_payload_0_379);
  assign _zz_dataOut_payload_0_1129 = (_zz_dataOut_payload_0_1128 ? _zz_dataOut_payload_0_376 : _zz_dataOut_payload_0_379);
  assign _zz_dataOut_payload_0_1130 = (_zz_dataOut_payload_0_1128 ? _zz_dataOut_payload_0_379 : _zz_dataOut_payload_0_376);
  assign _zz_dataOut_payload_0_1131 = (_zz_dataOut_payload_0_377 < _zz_dataOut_payload_0_378);
  assign _zz_dataOut_payload_0_1132 = (_zz_dataOut_payload_0_1131 ? _zz_dataOut_payload_0_377 : _zz_dataOut_payload_0_378);
  assign _zz_dataOut_payload_0_1133 = (_zz_dataOut_payload_0_1131 ? _zz_dataOut_payload_0_378 : _zz_dataOut_payload_0_377);
  assign _zz_dataOut_payload_0_1134 = (_zz_dataOut_payload_0_1129 < _zz_dataOut_payload_0_1132);
  assign _zz_dataOut_payload_0_1135 = (_zz_dataOut_payload_0_1133 < _zz_dataOut_payload_0_1130);
  assign _zz_dataOut_payload_0_1140 = (_zz_dataOut_payload_0_380 < _zz_dataOut_payload_0_383);
  assign _zz_dataOut_payload_0_1141 = (_zz_dataOut_payload_0_1140 ? _zz_dataOut_payload_0_380 : _zz_dataOut_payload_0_383);
  assign _zz_dataOut_payload_0_1142 = (_zz_dataOut_payload_0_1140 ? _zz_dataOut_payload_0_383 : _zz_dataOut_payload_0_380);
  assign _zz_dataOut_payload_0_1143 = (_zz_dataOut_payload_0_381 < _zz_dataOut_payload_0_382);
  assign _zz_dataOut_payload_0_1144 = (_zz_dataOut_payload_0_1143 ? _zz_dataOut_payload_0_381 : _zz_dataOut_payload_0_382);
  assign _zz_dataOut_payload_0_1145 = (_zz_dataOut_payload_0_1143 ? _zz_dataOut_payload_0_382 : _zz_dataOut_payload_0_381);
  assign _zz_dataOut_payload_0_1146 = (_zz_dataOut_payload_0_1141 < _zz_dataOut_payload_0_1144);
  assign _zz_dataOut_payload_0_1147 = (_zz_dataOut_payload_0_1145 < _zz_dataOut_payload_0_1142);
  assign _zz_dataOut_payload_0_1408 = (_zz_dataOut_payload_0_1152 < _zz_dataOut_payload_0_1159);
  assign _zz_dataOut_payload_0_1409 = (_zz_dataOut_payload_0_1408 ? _zz_dataOut_payload_0_1152 : _zz_dataOut_payload_0_1159);
  assign _zz_dataOut_payload_0_1410 = (_zz_dataOut_payload_0_1408 ? _zz_dataOut_payload_0_1159 : _zz_dataOut_payload_0_1152);
  assign _zz_dataOut_payload_0_1411 = (_zz_dataOut_payload_0_1153 < _zz_dataOut_payload_0_1158);
  assign _zz_dataOut_payload_0_1412 = (_zz_dataOut_payload_0_1411 ? _zz_dataOut_payload_0_1153 : _zz_dataOut_payload_0_1158);
  assign _zz_dataOut_payload_0_1413 = (_zz_dataOut_payload_0_1411 ? _zz_dataOut_payload_0_1158 : _zz_dataOut_payload_0_1153);
  assign _zz_dataOut_payload_0_1414 = (_zz_dataOut_payload_0_1154 < _zz_dataOut_payload_0_1157);
  assign _zz_dataOut_payload_0_1415 = (_zz_dataOut_payload_0_1414 ? _zz_dataOut_payload_0_1154 : _zz_dataOut_payload_0_1157);
  assign _zz_dataOut_payload_0_1416 = (_zz_dataOut_payload_0_1414 ? _zz_dataOut_payload_0_1157 : _zz_dataOut_payload_0_1154);
  assign _zz_dataOut_payload_0_1417 = (_zz_dataOut_payload_0_1155 < _zz_dataOut_payload_0_1156);
  assign _zz_dataOut_payload_0_1418 = (_zz_dataOut_payload_0_1417 ? _zz_dataOut_payload_0_1155 : _zz_dataOut_payload_0_1156);
  assign _zz_dataOut_payload_0_1419 = (_zz_dataOut_payload_0_1417 ? _zz_dataOut_payload_0_1156 : _zz_dataOut_payload_0_1155);
  assign _zz_dataOut_payload_0_1420 = (_zz_dataOut_payload_0_1409 < _zz_dataOut_payload_0_1415);
  assign _zz_dataOut_payload_0_1421 = (_zz_dataOut_payload_0_1420 ? _zz_dataOut_payload_0_1409 : _zz_dataOut_payload_0_1415);
  assign _zz_dataOut_payload_0_1422 = (_zz_dataOut_payload_0_1420 ? _zz_dataOut_payload_0_1415 : _zz_dataOut_payload_0_1409);
  assign _zz_dataOut_payload_0_1423 = (_zz_dataOut_payload_0_1412 < _zz_dataOut_payload_0_1418);
  assign _zz_dataOut_payload_0_1424 = (_zz_dataOut_payload_0_1423 ? _zz_dataOut_payload_0_1412 : _zz_dataOut_payload_0_1418);
  assign _zz_dataOut_payload_0_1425 = (_zz_dataOut_payload_0_1423 ? _zz_dataOut_payload_0_1418 : _zz_dataOut_payload_0_1412);
  assign _zz_dataOut_payload_0_1426 = (_zz_dataOut_payload_0_1421 < _zz_dataOut_payload_0_1424);
  assign _zz_dataOut_payload_0_1427 = (_zz_dataOut_payload_0_1422 < _zz_dataOut_payload_0_1425);
  assign _zz_dataOut_payload_0_1432 = (_zz_dataOut_payload_0_1419 < _zz_dataOut_payload_0_1413);
  assign _zz_dataOut_payload_0_1433 = (_zz_dataOut_payload_0_1432 ? _zz_dataOut_payload_0_1419 : _zz_dataOut_payload_0_1413);
  assign _zz_dataOut_payload_0_1434 = (_zz_dataOut_payload_0_1432 ? _zz_dataOut_payload_0_1413 : _zz_dataOut_payload_0_1419);
  assign _zz_dataOut_payload_0_1435 = (_zz_dataOut_payload_0_1416 < _zz_dataOut_payload_0_1410);
  assign _zz_dataOut_payload_0_1436 = (_zz_dataOut_payload_0_1435 ? _zz_dataOut_payload_0_1416 : _zz_dataOut_payload_0_1410);
  assign _zz_dataOut_payload_0_1437 = (_zz_dataOut_payload_0_1435 ? _zz_dataOut_payload_0_1410 : _zz_dataOut_payload_0_1416);
  assign _zz_dataOut_payload_0_1438 = (_zz_dataOut_payload_0_1433 < _zz_dataOut_payload_0_1436);
  assign _zz_dataOut_payload_0_1439 = (_zz_dataOut_payload_0_1434 < _zz_dataOut_payload_0_1437);
  assign _zz_dataOut_payload_0_1452 = (_zz_dataOut_payload_0_1160 < _zz_dataOut_payload_0_1167);
  assign _zz_dataOut_payload_0_1453 = (_zz_dataOut_payload_0_1452 ? _zz_dataOut_payload_0_1160 : _zz_dataOut_payload_0_1167);
  assign _zz_dataOut_payload_0_1454 = (_zz_dataOut_payload_0_1452 ? _zz_dataOut_payload_0_1167 : _zz_dataOut_payload_0_1160);
  assign _zz_dataOut_payload_0_1455 = (_zz_dataOut_payload_0_1161 < _zz_dataOut_payload_0_1166);
  assign _zz_dataOut_payload_0_1456 = (_zz_dataOut_payload_0_1455 ? _zz_dataOut_payload_0_1161 : _zz_dataOut_payload_0_1166);
  assign _zz_dataOut_payload_0_1457 = (_zz_dataOut_payload_0_1455 ? _zz_dataOut_payload_0_1166 : _zz_dataOut_payload_0_1161);
  assign _zz_dataOut_payload_0_1458 = (_zz_dataOut_payload_0_1162 < _zz_dataOut_payload_0_1165);
  assign _zz_dataOut_payload_0_1459 = (_zz_dataOut_payload_0_1458 ? _zz_dataOut_payload_0_1162 : _zz_dataOut_payload_0_1165);
  assign _zz_dataOut_payload_0_1460 = (_zz_dataOut_payload_0_1458 ? _zz_dataOut_payload_0_1165 : _zz_dataOut_payload_0_1162);
  assign _zz_dataOut_payload_0_1461 = (_zz_dataOut_payload_0_1163 < _zz_dataOut_payload_0_1164);
  assign _zz_dataOut_payload_0_1462 = (_zz_dataOut_payload_0_1461 ? _zz_dataOut_payload_0_1163 : _zz_dataOut_payload_0_1164);
  assign _zz_dataOut_payload_0_1463 = (_zz_dataOut_payload_0_1461 ? _zz_dataOut_payload_0_1164 : _zz_dataOut_payload_0_1163);
  assign _zz_dataOut_payload_0_1464 = (_zz_dataOut_payload_0_1453 < _zz_dataOut_payload_0_1459);
  assign _zz_dataOut_payload_0_1465 = (_zz_dataOut_payload_0_1464 ? _zz_dataOut_payload_0_1453 : _zz_dataOut_payload_0_1459);
  assign _zz_dataOut_payload_0_1466 = (_zz_dataOut_payload_0_1464 ? _zz_dataOut_payload_0_1459 : _zz_dataOut_payload_0_1453);
  assign _zz_dataOut_payload_0_1467 = (_zz_dataOut_payload_0_1456 < _zz_dataOut_payload_0_1462);
  assign _zz_dataOut_payload_0_1468 = (_zz_dataOut_payload_0_1467 ? _zz_dataOut_payload_0_1456 : _zz_dataOut_payload_0_1462);
  assign _zz_dataOut_payload_0_1469 = (_zz_dataOut_payload_0_1467 ? _zz_dataOut_payload_0_1462 : _zz_dataOut_payload_0_1456);
  assign _zz_dataOut_payload_0_1470 = (_zz_dataOut_payload_0_1465 < _zz_dataOut_payload_0_1468);
  assign _zz_dataOut_payload_0_1471 = (_zz_dataOut_payload_0_1466 < _zz_dataOut_payload_0_1469);
  assign _zz_dataOut_payload_0_1476 = (_zz_dataOut_payload_0_1463 < _zz_dataOut_payload_0_1457);
  assign _zz_dataOut_payload_0_1477 = (_zz_dataOut_payload_0_1476 ? _zz_dataOut_payload_0_1463 : _zz_dataOut_payload_0_1457);
  assign _zz_dataOut_payload_0_1478 = (_zz_dataOut_payload_0_1476 ? _zz_dataOut_payload_0_1457 : _zz_dataOut_payload_0_1463);
  assign _zz_dataOut_payload_0_1479 = (_zz_dataOut_payload_0_1460 < _zz_dataOut_payload_0_1454);
  assign _zz_dataOut_payload_0_1480 = (_zz_dataOut_payload_0_1479 ? _zz_dataOut_payload_0_1460 : _zz_dataOut_payload_0_1454);
  assign _zz_dataOut_payload_0_1481 = (_zz_dataOut_payload_0_1479 ? _zz_dataOut_payload_0_1454 : _zz_dataOut_payload_0_1460);
  assign _zz_dataOut_payload_0_1482 = (_zz_dataOut_payload_0_1477 < _zz_dataOut_payload_0_1480);
  assign _zz_dataOut_payload_0_1483 = (_zz_dataOut_payload_0_1478 < _zz_dataOut_payload_0_1481);
  assign _zz_dataOut_payload_0_1496 = (_zz_dataOut_payload_0_1168 < _zz_dataOut_payload_0_1175);
  assign _zz_dataOut_payload_0_1497 = (_zz_dataOut_payload_0_1496 ? _zz_dataOut_payload_0_1168 : _zz_dataOut_payload_0_1175);
  assign _zz_dataOut_payload_0_1498 = (_zz_dataOut_payload_0_1496 ? _zz_dataOut_payload_0_1175 : _zz_dataOut_payload_0_1168);
  assign _zz_dataOut_payload_0_1499 = (_zz_dataOut_payload_0_1169 < _zz_dataOut_payload_0_1174);
  assign _zz_dataOut_payload_0_1500 = (_zz_dataOut_payload_0_1499 ? _zz_dataOut_payload_0_1169 : _zz_dataOut_payload_0_1174);
  assign _zz_dataOut_payload_0_1501 = (_zz_dataOut_payload_0_1499 ? _zz_dataOut_payload_0_1174 : _zz_dataOut_payload_0_1169);
  assign _zz_dataOut_payload_0_1502 = (_zz_dataOut_payload_0_1170 < _zz_dataOut_payload_0_1173);
  assign _zz_dataOut_payload_0_1503 = (_zz_dataOut_payload_0_1502 ? _zz_dataOut_payload_0_1170 : _zz_dataOut_payload_0_1173);
  assign _zz_dataOut_payload_0_1504 = (_zz_dataOut_payload_0_1502 ? _zz_dataOut_payload_0_1173 : _zz_dataOut_payload_0_1170);
  assign _zz_dataOut_payload_0_1505 = (_zz_dataOut_payload_0_1171 < _zz_dataOut_payload_0_1172);
  assign _zz_dataOut_payload_0_1506 = (_zz_dataOut_payload_0_1505 ? _zz_dataOut_payload_0_1171 : _zz_dataOut_payload_0_1172);
  assign _zz_dataOut_payload_0_1507 = (_zz_dataOut_payload_0_1505 ? _zz_dataOut_payload_0_1172 : _zz_dataOut_payload_0_1171);
  assign _zz_dataOut_payload_0_1508 = (_zz_dataOut_payload_0_1497 < _zz_dataOut_payload_0_1503);
  assign _zz_dataOut_payload_0_1509 = (_zz_dataOut_payload_0_1508 ? _zz_dataOut_payload_0_1497 : _zz_dataOut_payload_0_1503);
  assign _zz_dataOut_payload_0_1510 = (_zz_dataOut_payload_0_1508 ? _zz_dataOut_payload_0_1503 : _zz_dataOut_payload_0_1497);
  assign _zz_dataOut_payload_0_1511 = (_zz_dataOut_payload_0_1500 < _zz_dataOut_payload_0_1506);
  assign _zz_dataOut_payload_0_1512 = (_zz_dataOut_payload_0_1511 ? _zz_dataOut_payload_0_1500 : _zz_dataOut_payload_0_1506);
  assign _zz_dataOut_payload_0_1513 = (_zz_dataOut_payload_0_1511 ? _zz_dataOut_payload_0_1506 : _zz_dataOut_payload_0_1500);
  assign _zz_dataOut_payload_0_1514 = (_zz_dataOut_payload_0_1509 < _zz_dataOut_payload_0_1512);
  assign _zz_dataOut_payload_0_1515 = (_zz_dataOut_payload_0_1510 < _zz_dataOut_payload_0_1513);
  assign _zz_dataOut_payload_0_1520 = (_zz_dataOut_payload_0_1507 < _zz_dataOut_payload_0_1501);
  assign _zz_dataOut_payload_0_1521 = (_zz_dataOut_payload_0_1520 ? _zz_dataOut_payload_0_1507 : _zz_dataOut_payload_0_1501);
  assign _zz_dataOut_payload_0_1522 = (_zz_dataOut_payload_0_1520 ? _zz_dataOut_payload_0_1501 : _zz_dataOut_payload_0_1507);
  assign _zz_dataOut_payload_0_1523 = (_zz_dataOut_payload_0_1504 < _zz_dataOut_payload_0_1498);
  assign _zz_dataOut_payload_0_1524 = (_zz_dataOut_payload_0_1523 ? _zz_dataOut_payload_0_1504 : _zz_dataOut_payload_0_1498);
  assign _zz_dataOut_payload_0_1525 = (_zz_dataOut_payload_0_1523 ? _zz_dataOut_payload_0_1498 : _zz_dataOut_payload_0_1504);
  assign _zz_dataOut_payload_0_1526 = (_zz_dataOut_payload_0_1521 < _zz_dataOut_payload_0_1524);
  assign _zz_dataOut_payload_0_1527 = (_zz_dataOut_payload_0_1522 < _zz_dataOut_payload_0_1525);
  assign _zz_dataOut_payload_0_1540 = (_zz_dataOut_payload_0_1176 < _zz_dataOut_payload_0_1183);
  assign _zz_dataOut_payload_0_1541 = (_zz_dataOut_payload_0_1540 ? _zz_dataOut_payload_0_1176 : _zz_dataOut_payload_0_1183);
  assign _zz_dataOut_payload_0_1542 = (_zz_dataOut_payload_0_1540 ? _zz_dataOut_payload_0_1183 : _zz_dataOut_payload_0_1176);
  assign _zz_dataOut_payload_0_1543 = (_zz_dataOut_payload_0_1177 < _zz_dataOut_payload_0_1182);
  assign _zz_dataOut_payload_0_1544 = (_zz_dataOut_payload_0_1543 ? _zz_dataOut_payload_0_1177 : _zz_dataOut_payload_0_1182);
  assign _zz_dataOut_payload_0_1545 = (_zz_dataOut_payload_0_1543 ? _zz_dataOut_payload_0_1182 : _zz_dataOut_payload_0_1177);
  assign _zz_dataOut_payload_0_1546 = (_zz_dataOut_payload_0_1178 < _zz_dataOut_payload_0_1181);
  assign _zz_dataOut_payload_0_1547 = (_zz_dataOut_payload_0_1546 ? _zz_dataOut_payload_0_1178 : _zz_dataOut_payload_0_1181);
  assign _zz_dataOut_payload_0_1548 = (_zz_dataOut_payload_0_1546 ? _zz_dataOut_payload_0_1181 : _zz_dataOut_payload_0_1178);
  assign _zz_dataOut_payload_0_1549 = (_zz_dataOut_payload_0_1179 < _zz_dataOut_payload_0_1180);
  assign _zz_dataOut_payload_0_1550 = (_zz_dataOut_payload_0_1549 ? _zz_dataOut_payload_0_1179 : _zz_dataOut_payload_0_1180);
  assign _zz_dataOut_payload_0_1551 = (_zz_dataOut_payload_0_1549 ? _zz_dataOut_payload_0_1180 : _zz_dataOut_payload_0_1179);
  assign _zz_dataOut_payload_0_1552 = (_zz_dataOut_payload_0_1541 < _zz_dataOut_payload_0_1547);
  assign _zz_dataOut_payload_0_1553 = (_zz_dataOut_payload_0_1552 ? _zz_dataOut_payload_0_1541 : _zz_dataOut_payload_0_1547);
  assign _zz_dataOut_payload_0_1554 = (_zz_dataOut_payload_0_1552 ? _zz_dataOut_payload_0_1547 : _zz_dataOut_payload_0_1541);
  assign _zz_dataOut_payload_0_1555 = (_zz_dataOut_payload_0_1544 < _zz_dataOut_payload_0_1550);
  assign _zz_dataOut_payload_0_1556 = (_zz_dataOut_payload_0_1555 ? _zz_dataOut_payload_0_1544 : _zz_dataOut_payload_0_1550);
  assign _zz_dataOut_payload_0_1557 = (_zz_dataOut_payload_0_1555 ? _zz_dataOut_payload_0_1550 : _zz_dataOut_payload_0_1544);
  assign _zz_dataOut_payload_0_1558 = (_zz_dataOut_payload_0_1553 < _zz_dataOut_payload_0_1556);
  assign _zz_dataOut_payload_0_1559 = (_zz_dataOut_payload_0_1554 < _zz_dataOut_payload_0_1557);
  assign _zz_dataOut_payload_0_1564 = (_zz_dataOut_payload_0_1551 < _zz_dataOut_payload_0_1545);
  assign _zz_dataOut_payload_0_1565 = (_zz_dataOut_payload_0_1564 ? _zz_dataOut_payload_0_1551 : _zz_dataOut_payload_0_1545);
  assign _zz_dataOut_payload_0_1566 = (_zz_dataOut_payload_0_1564 ? _zz_dataOut_payload_0_1545 : _zz_dataOut_payload_0_1551);
  assign _zz_dataOut_payload_0_1567 = (_zz_dataOut_payload_0_1548 < _zz_dataOut_payload_0_1542);
  assign _zz_dataOut_payload_0_1568 = (_zz_dataOut_payload_0_1567 ? _zz_dataOut_payload_0_1548 : _zz_dataOut_payload_0_1542);
  assign _zz_dataOut_payload_0_1569 = (_zz_dataOut_payload_0_1567 ? _zz_dataOut_payload_0_1542 : _zz_dataOut_payload_0_1548);
  assign _zz_dataOut_payload_0_1570 = (_zz_dataOut_payload_0_1565 < _zz_dataOut_payload_0_1568);
  assign _zz_dataOut_payload_0_1571 = (_zz_dataOut_payload_0_1566 < _zz_dataOut_payload_0_1569);
  assign _zz_dataOut_payload_0_1584 = (_zz_dataOut_payload_0_1184 < _zz_dataOut_payload_0_1191);
  assign _zz_dataOut_payload_0_1585 = (_zz_dataOut_payload_0_1584 ? _zz_dataOut_payload_0_1184 : _zz_dataOut_payload_0_1191);
  assign _zz_dataOut_payload_0_1586 = (_zz_dataOut_payload_0_1584 ? _zz_dataOut_payload_0_1191 : _zz_dataOut_payload_0_1184);
  assign _zz_dataOut_payload_0_1587 = (_zz_dataOut_payload_0_1185 < _zz_dataOut_payload_0_1190);
  assign _zz_dataOut_payload_0_1588 = (_zz_dataOut_payload_0_1587 ? _zz_dataOut_payload_0_1185 : _zz_dataOut_payload_0_1190);
  assign _zz_dataOut_payload_0_1589 = (_zz_dataOut_payload_0_1587 ? _zz_dataOut_payload_0_1190 : _zz_dataOut_payload_0_1185);
  assign _zz_dataOut_payload_0_1590 = (_zz_dataOut_payload_0_1186 < _zz_dataOut_payload_0_1189);
  assign _zz_dataOut_payload_0_1591 = (_zz_dataOut_payload_0_1590 ? _zz_dataOut_payload_0_1186 : _zz_dataOut_payload_0_1189);
  assign _zz_dataOut_payload_0_1592 = (_zz_dataOut_payload_0_1590 ? _zz_dataOut_payload_0_1189 : _zz_dataOut_payload_0_1186);
  assign _zz_dataOut_payload_0_1593 = (_zz_dataOut_payload_0_1187 < _zz_dataOut_payload_0_1188);
  assign _zz_dataOut_payload_0_1594 = (_zz_dataOut_payload_0_1593 ? _zz_dataOut_payload_0_1187 : _zz_dataOut_payload_0_1188);
  assign _zz_dataOut_payload_0_1595 = (_zz_dataOut_payload_0_1593 ? _zz_dataOut_payload_0_1188 : _zz_dataOut_payload_0_1187);
  assign _zz_dataOut_payload_0_1596 = (_zz_dataOut_payload_0_1585 < _zz_dataOut_payload_0_1591);
  assign _zz_dataOut_payload_0_1597 = (_zz_dataOut_payload_0_1596 ? _zz_dataOut_payload_0_1585 : _zz_dataOut_payload_0_1591);
  assign _zz_dataOut_payload_0_1598 = (_zz_dataOut_payload_0_1596 ? _zz_dataOut_payload_0_1591 : _zz_dataOut_payload_0_1585);
  assign _zz_dataOut_payload_0_1599 = (_zz_dataOut_payload_0_1588 < _zz_dataOut_payload_0_1594);
  assign _zz_dataOut_payload_0_1600 = (_zz_dataOut_payload_0_1599 ? _zz_dataOut_payload_0_1588 : _zz_dataOut_payload_0_1594);
  assign _zz_dataOut_payload_0_1601 = (_zz_dataOut_payload_0_1599 ? _zz_dataOut_payload_0_1594 : _zz_dataOut_payload_0_1588);
  assign _zz_dataOut_payload_0_1602 = (_zz_dataOut_payload_0_1597 < _zz_dataOut_payload_0_1600);
  assign _zz_dataOut_payload_0_1603 = (_zz_dataOut_payload_0_1598 < _zz_dataOut_payload_0_1601);
  assign _zz_dataOut_payload_0_1608 = (_zz_dataOut_payload_0_1595 < _zz_dataOut_payload_0_1589);
  assign _zz_dataOut_payload_0_1609 = (_zz_dataOut_payload_0_1608 ? _zz_dataOut_payload_0_1595 : _zz_dataOut_payload_0_1589);
  assign _zz_dataOut_payload_0_1610 = (_zz_dataOut_payload_0_1608 ? _zz_dataOut_payload_0_1589 : _zz_dataOut_payload_0_1595);
  assign _zz_dataOut_payload_0_1611 = (_zz_dataOut_payload_0_1592 < _zz_dataOut_payload_0_1586);
  assign _zz_dataOut_payload_0_1612 = (_zz_dataOut_payload_0_1611 ? _zz_dataOut_payload_0_1592 : _zz_dataOut_payload_0_1586);
  assign _zz_dataOut_payload_0_1613 = (_zz_dataOut_payload_0_1611 ? _zz_dataOut_payload_0_1586 : _zz_dataOut_payload_0_1592);
  assign _zz_dataOut_payload_0_1614 = (_zz_dataOut_payload_0_1609 < _zz_dataOut_payload_0_1612);
  assign _zz_dataOut_payload_0_1615 = (_zz_dataOut_payload_0_1610 < _zz_dataOut_payload_0_1613);
  assign _zz_dataOut_payload_0_1628 = (_zz_dataOut_payload_0_1192 < _zz_dataOut_payload_0_1199);
  assign _zz_dataOut_payload_0_1629 = (_zz_dataOut_payload_0_1628 ? _zz_dataOut_payload_0_1192 : _zz_dataOut_payload_0_1199);
  assign _zz_dataOut_payload_0_1630 = (_zz_dataOut_payload_0_1628 ? _zz_dataOut_payload_0_1199 : _zz_dataOut_payload_0_1192);
  assign _zz_dataOut_payload_0_1631 = (_zz_dataOut_payload_0_1193 < _zz_dataOut_payload_0_1198);
  assign _zz_dataOut_payload_0_1632 = (_zz_dataOut_payload_0_1631 ? _zz_dataOut_payload_0_1193 : _zz_dataOut_payload_0_1198);
  assign _zz_dataOut_payload_0_1633 = (_zz_dataOut_payload_0_1631 ? _zz_dataOut_payload_0_1198 : _zz_dataOut_payload_0_1193);
  assign _zz_dataOut_payload_0_1634 = (_zz_dataOut_payload_0_1194 < _zz_dataOut_payload_0_1197);
  assign _zz_dataOut_payload_0_1635 = (_zz_dataOut_payload_0_1634 ? _zz_dataOut_payload_0_1194 : _zz_dataOut_payload_0_1197);
  assign _zz_dataOut_payload_0_1636 = (_zz_dataOut_payload_0_1634 ? _zz_dataOut_payload_0_1197 : _zz_dataOut_payload_0_1194);
  assign _zz_dataOut_payload_0_1637 = (_zz_dataOut_payload_0_1195 < _zz_dataOut_payload_0_1196);
  assign _zz_dataOut_payload_0_1638 = (_zz_dataOut_payload_0_1637 ? _zz_dataOut_payload_0_1195 : _zz_dataOut_payload_0_1196);
  assign _zz_dataOut_payload_0_1639 = (_zz_dataOut_payload_0_1637 ? _zz_dataOut_payload_0_1196 : _zz_dataOut_payload_0_1195);
  assign _zz_dataOut_payload_0_1640 = (_zz_dataOut_payload_0_1629 < _zz_dataOut_payload_0_1635);
  assign _zz_dataOut_payload_0_1641 = (_zz_dataOut_payload_0_1640 ? _zz_dataOut_payload_0_1629 : _zz_dataOut_payload_0_1635);
  assign _zz_dataOut_payload_0_1642 = (_zz_dataOut_payload_0_1640 ? _zz_dataOut_payload_0_1635 : _zz_dataOut_payload_0_1629);
  assign _zz_dataOut_payload_0_1643 = (_zz_dataOut_payload_0_1632 < _zz_dataOut_payload_0_1638);
  assign _zz_dataOut_payload_0_1644 = (_zz_dataOut_payload_0_1643 ? _zz_dataOut_payload_0_1632 : _zz_dataOut_payload_0_1638);
  assign _zz_dataOut_payload_0_1645 = (_zz_dataOut_payload_0_1643 ? _zz_dataOut_payload_0_1638 : _zz_dataOut_payload_0_1632);
  assign _zz_dataOut_payload_0_1646 = (_zz_dataOut_payload_0_1641 < _zz_dataOut_payload_0_1644);
  assign _zz_dataOut_payload_0_1647 = (_zz_dataOut_payload_0_1642 < _zz_dataOut_payload_0_1645);
  assign _zz_dataOut_payload_0_1652 = (_zz_dataOut_payload_0_1639 < _zz_dataOut_payload_0_1633);
  assign _zz_dataOut_payload_0_1653 = (_zz_dataOut_payload_0_1652 ? _zz_dataOut_payload_0_1639 : _zz_dataOut_payload_0_1633);
  assign _zz_dataOut_payload_0_1654 = (_zz_dataOut_payload_0_1652 ? _zz_dataOut_payload_0_1633 : _zz_dataOut_payload_0_1639);
  assign _zz_dataOut_payload_0_1655 = (_zz_dataOut_payload_0_1636 < _zz_dataOut_payload_0_1630);
  assign _zz_dataOut_payload_0_1656 = (_zz_dataOut_payload_0_1655 ? _zz_dataOut_payload_0_1636 : _zz_dataOut_payload_0_1630);
  assign _zz_dataOut_payload_0_1657 = (_zz_dataOut_payload_0_1655 ? _zz_dataOut_payload_0_1630 : _zz_dataOut_payload_0_1636);
  assign _zz_dataOut_payload_0_1658 = (_zz_dataOut_payload_0_1653 < _zz_dataOut_payload_0_1656);
  assign _zz_dataOut_payload_0_1659 = (_zz_dataOut_payload_0_1654 < _zz_dataOut_payload_0_1657);
  assign _zz_dataOut_payload_0_1672 = (_zz_dataOut_payload_0_1200 < _zz_dataOut_payload_0_1207);
  assign _zz_dataOut_payload_0_1673 = (_zz_dataOut_payload_0_1672 ? _zz_dataOut_payload_0_1200 : _zz_dataOut_payload_0_1207);
  assign _zz_dataOut_payload_0_1674 = (_zz_dataOut_payload_0_1672 ? _zz_dataOut_payload_0_1207 : _zz_dataOut_payload_0_1200);
  assign _zz_dataOut_payload_0_1675 = (_zz_dataOut_payload_0_1201 < _zz_dataOut_payload_0_1206);
  assign _zz_dataOut_payload_0_1676 = (_zz_dataOut_payload_0_1675 ? _zz_dataOut_payload_0_1201 : _zz_dataOut_payload_0_1206);
  assign _zz_dataOut_payload_0_1677 = (_zz_dataOut_payload_0_1675 ? _zz_dataOut_payload_0_1206 : _zz_dataOut_payload_0_1201);
  assign _zz_dataOut_payload_0_1678 = (_zz_dataOut_payload_0_1202 < _zz_dataOut_payload_0_1205);
  assign _zz_dataOut_payload_0_1679 = (_zz_dataOut_payload_0_1678 ? _zz_dataOut_payload_0_1202 : _zz_dataOut_payload_0_1205);
  assign _zz_dataOut_payload_0_1680 = (_zz_dataOut_payload_0_1678 ? _zz_dataOut_payload_0_1205 : _zz_dataOut_payload_0_1202);
  assign _zz_dataOut_payload_0_1681 = (_zz_dataOut_payload_0_1203 < _zz_dataOut_payload_0_1204);
  assign _zz_dataOut_payload_0_1682 = (_zz_dataOut_payload_0_1681 ? _zz_dataOut_payload_0_1203 : _zz_dataOut_payload_0_1204);
  assign _zz_dataOut_payload_0_1683 = (_zz_dataOut_payload_0_1681 ? _zz_dataOut_payload_0_1204 : _zz_dataOut_payload_0_1203);
  assign _zz_dataOut_payload_0_1684 = (_zz_dataOut_payload_0_1673 < _zz_dataOut_payload_0_1679);
  assign _zz_dataOut_payload_0_1685 = (_zz_dataOut_payload_0_1684 ? _zz_dataOut_payload_0_1673 : _zz_dataOut_payload_0_1679);
  assign _zz_dataOut_payload_0_1686 = (_zz_dataOut_payload_0_1684 ? _zz_dataOut_payload_0_1679 : _zz_dataOut_payload_0_1673);
  assign _zz_dataOut_payload_0_1687 = (_zz_dataOut_payload_0_1676 < _zz_dataOut_payload_0_1682);
  assign _zz_dataOut_payload_0_1688 = (_zz_dataOut_payload_0_1687 ? _zz_dataOut_payload_0_1676 : _zz_dataOut_payload_0_1682);
  assign _zz_dataOut_payload_0_1689 = (_zz_dataOut_payload_0_1687 ? _zz_dataOut_payload_0_1682 : _zz_dataOut_payload_0_1676);
  assign _zz_dataOut_payload_0_1690 = (_zz_dataOut_payload_0_1685 < _zz_dataOut_payload_0_1688);
  assign _zz_dataOut_payload_0_1691 = (_zz_dataOut_payload_0_1686 < _zz_dataOut_payload_0_1689);
  assign _zz_dataOut_payload_0_1696 = (_zz_dataOut_payload_0_1683 < _zz_dataOut_payload_0_1677);
  assign _zz_dataOut_payload_0_1697 = (_zz_dataOut_payload_0_1696 ? _zz_dataOut_payload_0_1683 : _zz_dataOut_payload_0_1677);
  assign _zz_dataOut_payload_0_1698 = (_zz_dataOut_payload_0_1696 ? _zz_dataOut_payload_0_1677 : _zz_dataOut_payload_0_1683);
  assign _zz_dataOut_payload_0_1699 = (_zz_dataOut_payload_0_1680 < _zz_dataOut_payload_0_1674);
  assign _zz_dataOut_payload_0_1700 = (_zz_dataOut_payload_0_1699 ? _zz_dataOut_payload_0_1680 : _zz_dataOut_payload_0_1674);
  assign _zz_dataOut_payload_0_1701 = (_zz_dataOut_payload_0_1699 ? _zz_dataOut_payload_0_1674 : _zz_dataOut_payload_0_1680);
  assign _zz_dataOut_payload_0_1702 = (_zz_dataOut_payload_0_1697 < _zz_dataOut_payload_0_1700);
  assign _zz_dataOut_payload_0_1703 = (_zz_dataOut_payload_0_1698 < _zz_dataOut_payload_0_1701);
  assign _zz_dataOut_payload_0_1716 = (_zz_dataOut_payload_0_1208 < _zz_dataOut_payload_0_1215);
  assign _zz_dataOut_payload_0_1717 = (_zz_dataOut_payload_0_1716 ? _zz_dataOut_payload_0_1208 : _zz_dataOut_payload_0_1215);
  assign _zz_dataOut_payload_0_1718 = (_zz_dataOut_payload_0_1716 ? _zz_dataOut_payload_0_1215 : _zz_dataOut_payload_0_1208);
  assign _zz_dataOut_payload_0_1719 = (_zz_dataOut_payload_0_1209 < _zz_dataOut_payload_0_1214);
  assign _zz_dataOut_payload_0_1720 = (_zz_dataOut_payload_0_1719 ? _zz_dataOut_payload_0_1209 : _zz_dataOut_payload_0_1214);
  assign _zz_dataOut_payload_0_1721 = (_zz_dataOut_payload_0_1719 ? _zz_dataOut_payload_0_1214 : _zz_dataOut_payload_0_1209);
  assign _zz_dataOut_payload_0_1722 = (_zz_dataOut_payload_0_1210 < _zz_dataOut_payload_0_1213);
  assign _zz_dataOut_payload_0_1723 = (_zz_dataOut_payload_0_1722 ? _zz_dataOut_payload_0_1210 : _zz_dataOut_payload_0_1213);
  assign _zz_dataOut_payload_0_1724 = (_zz_dataOut_payload_0_1722 ? _zz_dataOut_payload_0_1213 : _zz_dataOut_payload_0_1210);
  assign _zz_dataOut_payload_0_1725 = (_zz_dataOut_payload_0_1211 < _zz_dataOut_payload_0_1212);
  assign _zz_dataOut_payload_0_1726 = (_zz_dataOut_payload_0_1725 ? _zz_dataOut_payload_0_1211 : _zz_dataOut_payload_0_1212);
  assign _zz_dataOut_payload_0_1727 = (_zz_dataOut_payload_0_1725 ? _zz_dataOut_payload_0_1212 : _zz_dataOut_payload_0_1211);
  assign _zz_dataOut_payload_0_1728 = (_zz_dataOut_payload_0_1717 < _zz_dataOut_payload_0_1723);
  assign _zz_dataOut_payload_0_1729 = (_zz_dataOut_payload_0_1728 ? _zz_dataOut_payload_0_1717 : _zz_dataOut_payload_0_1723);
  assign _zz_dataOut_payload_0_1730 = (_zz_dataOut_payload_0_1728 ? _zz_dataOut_payload_0_1723 : _zz_dataOut_payload_0_1717);
  assign _zz_dataOut_payload_0_1731 = (_zz_dataOut_payload_0_1720 < _zz_dataOut_payload_0_1726);
  assign _zz_dataOut_payload_0_1732 = (_zz_dataOut_payload_0_1731 ? _zz_dataOut_payload_0_1720 : _zz_dataOut_payload_0_1726);
  assign _zz_dataOut_payload_0_1733 = (_zz_dataOut_payload_0_1731 ? _zz_dataOut_payload_0_1726 : _zz_dataOut_payload_0_1720);
  assign _zz_dataOut_payload_0_1734 = (_zz_dataOut_payload_0_1729 < _zz_dataOut_payload_0_1732);
  assign _zz_dataOut_payload_0_1735 = (_zz_dataOut_payload_0_1730 < _zz_dataOut_payload_0_1733);
  assign _zz_dataOut_payload_0_1740 = (_zz_dataOut_payload_0_1727 < _zz_dataOut_payload_0_1721);
  assign _zz_dataOut_payload_0_1741 = (_zz_dataOut_payload_0_1740 ? _zz_dataOut_payload_0_1727 : _zz_dataOut_payload_0_1721);
  assign _zz_dataOut_payload_0_1742 = (_zz_dataOut_payload_0_1740 ? _zz_dataOut_payload_0_1721 : _zz_dataOut_payload_0_1727);
  assign _zz_dataOut_payload_0_1743 = (_zz_dataOut_payload_0_1724 < _zz_dataOut_payload_0_1718);
  assign _zz_dataOut_payload_0_1744 = (_zz_dataOut_payload_0_1743 ? _zz_dataOut_payload_0_1724 : _zz_dataOut_payload_0_1718);
  assign _zz_dataOut_payload_0_1745 = (_zz_dataOut_payload_0_1743 ? _zz_dataOut_payload_0_1718 : _zz_dataOut_payload_0_1724);
  assign _zz_dataOut_payload_0_1746 = (_zz_dataOut_payload_0_1741 < _zz_dataOut_payload_0_1744);
  assign _zz_dataOut_payload_0_1747 = (_zz_dataOut_payload_0_1742 < _zz_dataOut_payload_0_1745);
  assign _zz_dataOut_payload_0_1760 = (_zz_dataOut_payload_0_1216 < _zz_dataOut_payload_0_1223);
  assign _zz_dataOut_payload_0_1761 = (_zz_dataOut_payload_0_1760 ? _zz_dataOut_payload_0_1216 : _zz_dataOut_payload_0_1223);
  assign _zz_dataOut_payload_0_1762 = (_zz_dataOut_payload_0_1760 ? _zz_dataOut_payload_0_1223 : _zz_dataOut_payload_0_1216);
  assign _zz_dataOut_payload_0_1763 = (_zz_dataOut_payload_0_1217 < _zz_dataOut_payload_0_1222);
  assign _zz_dataOut_payload_0_1764 = (_zz_dataOut_payload_0_1763 ? _zz_dataOut_payload_0_1217 : _zz_dataOut_payload_0_1222);
  assign _zz_dataOut_payload_0_1765 = (_zz_dataOut_payload_0_1763 ? _zz_dataOut_payload_0_1222 : _zz_dataOut_payload_0_1217);
  assign _zz_dataOut_payload_0_1766 = (_zz_dataOut_payload_0_1218 < _zz_dataOut_payload_0_1221);
  assign _zz_dataOut_payload_0_1767 = (_zz_dataOut_payload_0_1766 ? _zz_dataOut_payload_0_1218 : _zz_dataOut_payload_0_1221);
  assign _zz_dataOut_payload_0_1768 = (_zz_dataOut_payload_0_1766 ? _zz_dataOut_payload_0_1221 : _zz_dataOut_payload_0_1218);
  assign _zz_dataOut_payload_0_1769 = (_zz_dataOut_payload_0_1219 < _zz_dataOut_payload_0_1220);
  assign _zz_dataOut_payload_0_1770 = (_zz_dataOut_payload_0_1769 ? _zz_dataOut_payload_0_1219 : _zz_dataOut_payload_0_1220);
  assign _zz_dataOut_payload_0_1771 = (_zz_dataOut_payload_0_1769 ? _zz_dataOut_payload_0_1220 : _zz_dataOut_payload_0_1219);
  assign _zz_dataOut_payload_0_1772 = (_zz_dataOut_payload_0_1761 < _zz_dataOut_payload_0_1767);
  assign _zz_dataOut_payload_0_1773 = (_zz_dataOut_payload_0_1772 ? _zz_dataOut_payload_0_1761 : _zz_dataOut_payload_0_1767);
  assign _zz_dataOut_payload_0_1774 = (_zz_dataOut_payload_0_1772 ? _zz_dataOut_payload_0_1767 : _zz_dataOut_payload_0_1761);
  assign _zz_dataOut_payload_0_1775 = (_zz_dataOut_payload_0_1764 < _zz_dataOut_payload_0_1770);
  assign _zz_dataOut_payload_0_1776 = (_zz_dataOut_payload_0_1775 ? _zz_dataOut_payload_0_1764 : _zz_dataOut_payload_0_1770);
  assign _zz_dataOut_payload_0_1777 = (_zz_dataOut_payload_0_1775 ? _zz_dataOut_payload_0_1770 : _zz_dataOut_payload_0_1764);
  assign _zz_dataOut_payload_0_1778 = (_zz_dataOut_payload_0_1773 < _zz_dataOut_payload_0_1776);
  assign _zz_dataOut_payload_0_1779 = (_zz_dataOut_payload_0_1774 < _zz_dataOut_payload_0_1777);
  assign _zz_dataOut_payload_0_1784 = (_zz_dataOut_payload_0_1771 < _zz_dataOut_payload_0_1765);
  assign _zz_dataOut_payload_0_1785 = (_zz_dataOut_payload_0_1784 ? _zz_dataOut_payload_0_1771 : _zz_dataOut_payload_0_1765);
  assign _zz_dataOut_payload_0_1786 = (_zz_dataOut_payload_0_1784 ? _zz_dataOut_payload_0_1765 : _zz_dataOut_payload_0_1771);
  assign _zz_dataOut_payload_0_1787 = (_zz_dataOut_payload_0_1768 < _zz_dataOut_payload_0_1762);
  assign _zz_dataOut_payload_0_1788 = (_zz_dataOut_payload_0_1787 ? _zz_dataOut_payload_0_1768 : _zz_dataOut_payload_0_1762);
  assign _zz_dataOut_payload_0_1789 = (_zz_dataOut_payload_0_1787 ? _zz_dataOut_payload_0_1762 : _zz_dataOut_payload_0_1768);
  assign _zz_dataOut_payload_0_1790 = (_zz_dataOut_payload_0_1785 < _zz_dataOut_payload_0_1788);
  assign _zz_dataOut_payload_0_1791 = (_zz_dataOut_payload_0_1786 < _zz_dataOut_payload_0_1789);
  assign _zz_dataOut_payload_0_1804 = (_zz_dataOut_payload_0_1224 < _zz_dataOut_payload_0_1231);
  assign _zz_dataOut_payload_0_1805 = (_zz_dataOut_payload_0_1804 ? _zz_dataOut_payload_0_1224 : _zz_dataOut_payload_0_1231);
  assign _zz_dataOut_payload_0_1806 = (_zz_dataOut_payload_0_1804 ? _zz_dataOut_payload_0_1231 : _zz_dataOut_payload_0_1224);
  assign _zz_dataOut_payload_0_1807 = (_zz_dataOut_payload_0_1225 < _zz_dataOut_payload_0_1230);
  assign _zz_dataOut_payload_0_1808 = (_zz_dataOut_payload_0_1807 ? _zz_dataOut_payload_0_1225 : _zz_dataOut_payload_0_1230);
  assign _zz_dataOut_payload_0_1809 = (_zz_dataOut_payload_0_1807 ? _zz_dataOut_payload_0_1230 : _zz_dataOut_payload_0_1225);
  assign _zz_dataOut_payload_0_1810 = (_zz_dataOut_payload_0_1226 < _zz_dataOut_payload_0_1229);
  assign _zz_dataOut_payload_0_1811 = (_zz_dataOut_payload_0_1810 ? _zz_dataOut_payload_0_1226 : _zz_dataOut_payload_0_1229);
  assign _zz_dataOut_payload_0_1812 = (_zz_dataOut_payload_0_1810 ? _zz_dataOut_payload_0_1229 : _zz_dataOut_payload_0_1226);
  assign _zz_dataOut_payload_0_1813 = (_zz_dataOut_payload_0_1227 < _zz_dataOut_payload_0_1228);
  assign _zz_dataOut_payload_0_1814 = (_zz_dataOut_payload_0_1813 ? _zz_dataOut_payload_0_1227 : _zz_dataOut_payload_0_1228);
  assign _zz_dataOut_payload_0_1815 = (_zz_dataOut_payload_0_1813 ? _zz_dataOut_payload_0_1228 : _zz_dataOut_payload_0_1227);
  assign _zz_dataOut_payload_0_1816 = (_zz_dataOut_payload_0_1805 < _zz_dataOut_payload_0_1811);
  assign _zz_dataOut_payload_0_1817 = (_zz_dataOut_payload_0_1816 ? _zz_dataOut_payload_0_1805 : _zz_dataOut_payload_0_1811);
  assign _zz_dataOut_payload_0_1818 = (_zz_dataOut_payload_0_1816 ? _zz_dataOut_payload_0_1811 : _zz_dataOut_payload_0_1805);
  assign _zz_dataOut_payload_0_1819 = (_zz_dataOut_payload_0_1808 < _zz_dataOut_payload_0_1814);
  assign _zz_dataOut_payload_0_1820 = (_zz_dataOut_payload_0_1819 ? _zz_dataOut_payload_0_1808 : _zz_dataOut_payload_0_1814);
  assign _zz_dataOut_payload_0_1821 = (_zz_dataOut_payload_0_1819 ? _zz_dataOut_payload_0_1814 : _zz_dataOut_payload_0_1808);
  assign _zz_dataOut_payload_0_1822 = (_zz_dataOut_payload_0_1817 < _zz_dataOut_payload_0_1820);
  assign _zz_dataOut_payload_0_1823 = (_zz_dataOut_payload_0_1818 < _zz_dataOut_payload_0_1821);
  assign _zz_dataOut_payload_0_1828 = (_zz_dataOut_payload_0_1815 < _zz_dataOut_payload_0_1809);
  assign _zz_dataOut_payload_0_1829 = (_zz_dataOut_payload_0_1828 ? _zz_dataOut_payload_0_1815 : _zz_dataOut_payload_0_1809);
  assign _zz_dataOut_payload_0_1830 = (_zz_dataOut_payload_0_1828 ? _zz_dataOut_payload_0_1809 : _zz_dataOut_payload_0_1815);
  assign _zz_dataOut_payload_0_1831 = (_zz_dataOut_payload_0_1812 < _zz_dataOut_payload_0_1806);
  assign _zz_dataOut_payload_0_1832 = (_zz_dataOut_payload_0_1831 ? _zz_dataOut_payload_0_1812 : _zz_dataOut_payload_0_1806);
  assign _zz_dataOut_payload_0_1833 = (_zz_dataOut_payload_0_1831 ? _zz_dataOut_payload_0_1806 : _zz_dataOut_payload_0_1812);
  assign _zz_dataOut_payload_0_1834 = (_zz_dataOut_payload_0_1829 < _zz_dataOut_payload_0_1832);
  assign _zz_dataOut_payload_0_1835 = (_zz_dataOut_payload_0_1830 < _zz_dataOut_payload_0_1833);
  assign _zz_dataOut_payload_0_1848 = (_zz_dataOut_payload_0_1232 < _zz_dataOut_payload_0_1239);
  assign _zz_dataOut_payload_0_1849 = (_zz_dataOut_payload_0_1848 ? _zz_dataOut_payload_0_1232 : _zz_dataOut_payload_0_1239);
  assign _zz_dataOut_payload_0_1850 = (_zz_dataOut_payload_0_1848 ? _zz_dataOut_payload_0_1239 : _zz_dataOut_payload_0_1232);
  assign _zz_dataOut_payload_0_1851 = (_zz_dataOut_payload_0_1233 < _zz_dataOut_payload_0_1238);
  assign _zz_dataOut_payload_0_1852 = (_zz_dataOut_payload_0_1851 ? _zz_dataOut_payload_0_1233 : _zz_dataOut_payload_0_1238);
  assign _zz_dataOut_payload_0_1853 = (_zz_dataOut_payload_0_1851 ? _zz_dataOut_payload_0_1238 : _zz_dataOut_payload_0_1233);
  assign _zz_dataOut_payload_0_1854 = (_zz_dataOut_payload_0_1234 < _zz_dataOut_payload_0_1237);
  assign _zz_dataOut_payload_0_1855 = (_zz_dataOut_payload_0_1854 ? _zz_dataOut_payload_0_1234 : _zz_dataOut_payload_0_1237);
  assign _zz_dataOut_payload_0_1856 = (_zz_dataOut_payload_0_1854 ? _zz_dataOut_payload_0_1237 : _zz_dataOut_payload_0_1234);
  assign _zz_dataOut_payload_0_1857 = (_zz_dataOut_payload_0_1235 < _zz_dataOut_payload_0_1236);
  assign _zz_dataOut_payload_0_1858 = (_zz_dataOut_payload_0_1857 ? _zz_dataOut_payload_0_1235 : _zz_dataOut_payload_0_1236);
  assign _zz_dataOut_payload_0_1859 = (_zz_dataOut_payload_0_1857 ? _zz_dataOut_payload_0_1236 : _zz_dataOut_payload_0_1235);
  assign _zz_dataOut_payload_0_1860 = (_zz_dataOut_payload_0_1849 < _zz_dataOut_payload_0_1855);
  assign _zz_dataOut_payload_0_1861 = (_zz_dataOut_payload_0_1860 ? _zz_dataOut_payload_0_1849 : _zz_dataOut_payload_0_1855);
  assign _zz_dataOut_payload_0_1862 = (_zz_dataOut_payload_0_1860 ? _zz_dataOut_payload_0_1855 : _zz_dataOut_payload_0_1849);
  assign _zz_dataOut_payload_0_1863 = (_zz_dataOut_payload_0_1852 < _zz_dataOut_payload_0_1858);
  assign _zz_dataOut_payload_0_1864 = (_zz_dataOut_payload_0_1863 ? _zz_dataOut_payload_0_1852 : _zz_dataOut_payload_0_1858);
  assign _zz_dataOut_payload_0_1865 = (_zz_dataOut_payload_0_1863 ? _zz_dataOut_payload_0_1858 : _zz_dataOut_payload_0_1852);
  assign _zz_dataOut_payload_0_1866 = (_zz_dataOut_payload_0_1861 < _zz_dataOut_payload_0_1864);
  assign _zz_dataOut_payload_0_1867 = (_zz_dataOut_payload_0_1862 < _zz_dataOut_payload_0_1865);
  assign _zz_dataOut_payload_0_1872 = (_zz_dataOut_payload_0_1859 < _zz_dataOut_payload_0_1853);
  assign _zz_dataOut_payload_0_1873 = (_zz_dataOut_payload_0_1872 ? _zz_dataOut_payload_0_1859 : _zz_dataOut_payload_0_1853);
  assign _zz_dataOut_payload_0_1874 = (_zz_dataOut_payload_0_1872 ? _zz_dataOut_payload_0_1853 : _zz_dataOut_payload_0_1859);
  assign _zz_dataOut_payload_0_1875 = (_zz_dataOut_payload_0_1856 < _zz_dataOut_payload_0_1850);
  assign _zz_dataOut_payload_0_1876 = (_zz_dataOut_payload_0_1875 ? _zz_dataOut_payload_0_1856 : _zz_dataOut_payload_0_1850);
  assign _zz_dataOut_payload_0_1877 = (_zz_dataOut_payload_0_1875 ? _zz_dataOut_payload_0_1850 : _zz_dataOut_payload_0_1856);
  assign _zz_dataOut_payload_0_1878 = (_zz_dataOut_payload_0_1873 < _zz_dataOut_payload_0_1876);
  assign _zz_dataOut_payload_0_1879 = (_zz_dataOut_payload_0_1874 < _zz_dataOut_payload_0_1877);
  assign _zz_dataOut_payload_0_1892 = (_zz_dataOut_payload_0_1240 < _zz_dataOut_payload_0_1247);
  assign _zz_dataOut_payload_0_1893 = (_zz_dataOut_payload_0_1892 ? _zz_dataOut_payload_0_1240 : _zz_dataOut_payload_0_1247);
  assign _zz_dataOut_payload_0_1894 = (_zz_dataOut_payload_0_1892 ? _zz_dataOut_payload_0_1247 : _zz_dataOut_payload_0_1240);
  assign _zz_dataOut_payload_0_1895 = (_zz_dataOut_payload_0_1241 < _zz_dataOut_payload_0_1246);
  assign _zz_dataOut_payload_0_1896 = (_zz_dataOut_payload_0_1895 ? _zz_dataOut_payload_0_1241 : _zz_dataOut_payload_0_1246);
  assign _zz_dataOut_payload_0_1897 = (_zz_dataOut_payload_0_1895 ? _zz_dataOut_payload_0_1246 : _zz_dataOut_payload_0_1241);
  assign _zz_dataOut_payload_0_1898 = (_zz_dataOut_payload_0_1242 < _zz_dataOut_payload_0_1245);
  assign _zz_dataOut_payload_0_1899 = (_zz_dataOut_payload_0_1898 ? _zz_dataOut_payload_0_1242 : _zz_dataOut_payload_0_1245);
  assign _zz_dataOut_payload_0_1900 = (_zz_dataOut_payload_0_1898 ? _zz_dataOut_payload_0_1245 : _zz_dataOut_payload_0_1242);
  assign _zz_dataOut_payload_0_1901 = (_zz_dataOut_payload_0_1243 < _zz_dataOut_payload_0_1244);
  assign _zz_dataOut_payload_0_1902 = (_zz_dataOut_payload_0_1901 ? _zz_dataOut_payload_0_1243 : _zz_dataOut_payload_0_1244);
  assign _zz_dataOut_payload_0_1903 = (_zz_dataOut_payload_0_1901 ? _zz_dataOut_payload_0_1244 : _zz_dataOut_payload_0_1243);
  assign _zz_dataOut_payload_0_1904 = (_zz_dataOut_payload_0_1893 < _zz_dataOut_payload_0_1899);
  assign _zz_dataOut_payload_0_1905 = (_zz_dataOut_payload_0_1904 ? _zz_dataOut_payload_0_1893 : _zz_dataOut_payload_0_1899);
  assign _zz_dataOut_payload_0_1906 = (_zz_dataOut_payload_0_1904 ? _zz_dataOut_payload_0_1899 : _zz_dataOut_payload_0_1893);
  assign _zz_dataOut_payload_0_1907 = (_zz_dataOut_payload_0_1896 < _zz_dataOut_payload_0_1902);
  assign _zz_dataOut_payload_0_1908 = (_zz_dataOut_payload_0_1907 ? _zz_dataOut_payload_0_1896 : _zz_dataOut_payload_0_1902);
  assign _zz_dataOut_payload_0_1909 = (_zz_dataOut_payload_0_1907 ? _zz_dataOut_payload_0_1902 : _zz_dataOut_payload_0_1896);
  assign _zz_dataOut_payload_0_1910 = (_zz_dataOut_payload_0_1905 < _zz_dataOut_payload_0_1908);
  assign _zz_dataOut_payload_0_1911 = (_zz_dataOut_payload_0_1906 < _zz_dataOut_payload_0_1909);
  assign _zz_dataOut_payload_0_1916 = (_zz_dataOut_payload_0_1903 < _zz_dataOut_payload_0_1897);
  assign _zz_dataOut_payload_0_1917 = (_zz_dataOut_payload_0_1916 ? _zz_dataOut_payload_0_1903 : _zz_dataOut_payload_0_1897);
  assign _zz_dataOut_payload_0_1918 = (_zz_dataOut_payload_0_1916 ? _zz_dataOut_payload_0_1897 : _zz_dataOut_payload_0_1903);
  assign _zz_dataOut_payload_0_1919 = (_zz_dataOut_payload_0_1900 < _zz_dataOut_payload_0_1894);
  assign _zz_dataOut_payload_0_1920 = (_zz_dataOut_payload_0_1919 ? _zz_dataOut_payload_0_1900 : _zz_dataOut_payload_0_1894);
  assign _zz_dataOut_payload_0_1921 = (_zz_dataOut_payload_0_1919 ? _zz_dataOut_payload_0_1894 : _zz_dataOut_payload_0_1900);
  assign _zz_dataOut_payload_0_1922 = (_zz_dataOut_payload_0_1917 < _zz_dataOut_payload_0_1920);
  assign _zz_dataOut_payload_0_1923 = (_zz_dataOut_payload_0_1918 < _zz_dataOut_payload_0_1921);
  assign _zz_dataOut_payload_0_1936 = (_zz_dataOut_payload_0_1248 < _zz_dataOut_payload_0_1255);
  assign _zz_dataOut_payload_0_1937 = (_zz_dataOut_payload_0_1936 ? _zz_dataOut_payload_0_1248 : _zz_dataOut_payload_0_1255);
  assign _zz_dataOut_payload_0_1938 = (_zz_dataOut_payload_0_1936 ? _zz_dataOut_payload_0_1255 : _zz_dataOut_payload_0_1248);
  assign _zz_dataOut_payload_0_1939 = (_zz_dataOut_payload_0_1249 < _zz_dataOut_payload_0_1254);
  assign _zz_dataOut_payload_0_1940 = (_zz_dataOut_payload_0_1939 ? _zz_dataOut_payload_0_1249 : _zz_dataOut_payload_0_1254);
  assign _zz_dataOut_payload_0_1941 = (_zz_dataOut_payload_0_1939 ? _zz_dataOut_payload_0_1254 : _zz_dataOut_payload_0_1249);
  assign _zz_dataOut_payload_0_1942 = (_zz_dataOut_payload_0_1250 < _zz_dataOut_payload_0_1253);
  assign _zz_dataOut_payload_0_1943 = (_zz_dataOut_payload_0_1942 ? _zz_dataOut_payload_0_1250 : _zz_dataOut_payload_0_1253);
  assign _zz_dataOut_payload_0_1944 = (_zz_dataOut_payload_0_1942 ? _zz_dataOut_payload_0_1253 : _zz_dataOut_payload_0_1250);
  assign _zz_dataOut_payload_0_1945 = (_zz_dataOut_payload_0_1251 < _zz_dataOut_payload_0_1252);
  assign _zz_dataOut_payload_0_1946 = (_zz_dataOut_payload_0_1945 ? _zz_dataOut_payload_0_1251 : _zz_dataOut_payload_0_1252);
  assign _zz_dataOut_payload_0_1947 = (_zz_dataOut_payload_0_1945 ? _zz_dataOut_payload_0_1252 : _zz_dataOut_payload_0_1251);
  assign _zz_dataOut_payload_0_1948 = (_zz_dataOut_payload_0_1937 < _zz_dataOut_payload_0_1943);
  assign _zz_dataOut_payload_0_1949 = (_zz_dataOut_payload_0_1948 ? _zz_dataOut_payload_0_1937 : _zz_dataOut_payload_0_1943);
  assign _zz_dataOut_payload_0_1950 = (_zz_dataOut_payload_0_1948 ? _zz_dataOut_payload_0_1943 : _zz_dataOut_payload_0_1937);
  assign _zz_dataOut_payload_0_1951 = (_zz_dataOut_payload_0_1940 < _zz_dataOut_payload_0_1946);
  assign _zz_dataOut_payload_0_1952 = (_zz_dataOut_payload_0_1951 ? _zz_dataOut_payload_0_1940 : _zz_dataOut_payload_0_1946);
  assign _zz_dataOut_payload_0_1953 = (_zz_dataOut_payload_0_1951 ? _zz_dataOut_payload_0_1946 : _zz_dataOut_payload_0_1940);
  assign _zz_dataOut_payload_0_1954 = (_zz_dataOut_payload_0_1949 < _zz_dataOut_payload_0_1952);
  assign _zz_dataOut_payload_0_1955 = (_zz_dataOut_payload_0_1950 < _zz_dataOut_payload_0_1953);
  assign _zz_dataOut_payload_0_1960 = (_zz_dataOut_payload_0_1947 < _zz_dataOut_payload_0_1941);
  assign _zz_dataOut_payload_0_1961 = (_zz_dataOut_payload_0_1960 ? _zz_dataOut_payload_0_1947 : _zz_dataOut_payload_0_1941);
  assign _zz_dataOut_payload_0_1962 = (_zz_dataOut_payload_0_1960 ? _zz_dataOut_payload_0_1941 : _zz_dataOut_payload_0_1947);
  assign _zz_dataOut_payload_0_1963 = (_zz_dataOut_payload_0_1944 < _zz_dataOut_payload_0_1938);
  assign _zz_dataOut_payload_0_1964 = (_zz_dataOut_payload_0_1963 ? _zz_dataOut_payload_0_1944 : _zz_dataOut_payload_0_1938);
  assign _zz_dataOut_payload_0_1965 = (_zz_dataOut_payload_0_1963 ? _zz_dataOut_payload_0_1938 : _zz_dataOut_payload_0_1944);
  assign _zz_dataOut_payload_0_1966 = (_zz_dataOut_payload_0_1961 < _zz_dataOut_payload_0_1964);
  assign _zz_dataOut_payload_0_1967 = (_zz_dataOut_payload_0_1962 < _zz_dataOut_payload_0_1965);
  assign _zz_dataOut_payload_0_1980 = (_zz_dataOut_payload_0_1256 < _zz_dataOut_payload_0_1263);
  assign _zz_dataOut_payload_0_1981 = (_zz_dataOut_payload_0_1980 ? _zz_dataOut_payload_0_1256 : _zz_dataOut_payload_0_1263);
  assign _zz_dataOut_payload_0_1982 = (_zz_dataOut_payload_0_1980 ? _zz_dataOut_payload_0_1263 : _zz_dataOut_payload_0_1256);
  assign _zz_dataOut_payload_0_1983 = (_zz_dataOut_payload_0_1257 < _zz_dataOut_payload_0_1262);
  assign _zz_dataOut_payload_0_1984 = (_zz_dataOut_payload_0_1983 ? _zz_dataOut_payload_0_1257 : _zz_dataOut_payload_0_1262);
  assign _zz_dataOut_payload_0_1985 = (_zz_dataOut_payload_0_1983 ? _zz_dataOut_payload_0_1262 : _zz_dataOut_payload_0_1257);
  assign _zz_dataOut_payload_0_1986 = (_zz_dataOut_payload_0_1258 < _zz_dataOut_payload_0_1261);
  assign _zz_dataOut_payload_0_1987 = (_zz_dataOut_payload_0_1986 ? _zz_dataOut_payload_0_1258 : _zz_dataOut_payload_0_1261);
  assign _zz_dataOut_payload_0_1988 = (_zz_dataOut_payload_0_1986 ? _zz_dataOut_payload_0_1261 : _zz_dataOut_payload_0_1258);
  assign _zz_dataOut_payload_0_1989 = (_zz_dataOut_payload_0_1259 < _zz_dataOut_payload_0_1260);
  assign _zz_dataOut_payload_0_1990 = (_zz_dataOut_payload_0_1989 ? _zz_dataOut_payload_0_1259 : _zz_dataOut_payload_0_1260);
  assign _zz_dataOut_payload_0_1991 = (_zz_dataOut_payload_0_1989 ? _zz_dataOut_payload_0_1260 : _zz_dataOut_payload_0_1259);
  assign _zz_dataOut_payload_0_1992 = (_zz_dataOut_payload_0_1981 < _zz_dataOut_payload_0_1987);
  assign _zz_dataOut_payload_0_1993 = (_zz_dataOut_payload_0_1992 ? _zz_dataOut_payload_0_1981 : _zz_dataOut_payload_0_1987);
  assign _zz_dataOut_payload_0_1994 = (_zz_dataOut_payload_0_1992 ? _zz_dataOut_payload_0_1987 : _zz_dataOut_payload_0_1981);
  assign _zz_dataOut_payload_0_1995 = (_zz_dataOut_payload_0_1984 < _zz_dataOut_payload_0_1990);
  assign _zz_dataOut_payload_0_1996 = (_zz_dataOut_payload_0_1995 ? _zz_dataOut_payload_0_1984 : _zz_dataOut_payload_0_1990);
  assign _zz_dataOut_payload_0_1997 = (_zz_dataOut_payload_0_1995 ? _zz_dataOut_payload_0_1990 : _zz_dataOut_payload_0_1984);
  assign _zz_dataOut_payload_0_1998 = (_zz_dataOut_payload_0_1993 < _zz_dataOut_payload_0_1996);
  assign _zz_dataOut_payload_0_1999 = (_zz_dataOut_payload_0_1994 < _zz_dataOut_payload_0_1997);
  assign _zz_dataOut_payload_0_2004 = (_zz_dataOut_payload_0_1991 < _zz_dataOut_payload_0_1985);
  assign _zz_dataOut_payload_0_2005 = (_zz_dataOut_payload_0_2004 ? _zz_dataOut_payload_0_1991 : _zz_dataOut_payload_0_1985);
  assign _zz_dataOut_payload_0_2006 = (_zz_dataOut_payload_0_2004 ? _zz_dataOut_payload_0_1985 : _zz_dataOut_payload_0_1991);
  assign _zz_dataOut_payload_0_2007 = (_zz_dataOut_payload_0_1988 < _zz_dataOut_payload_0_1982);
  assign _zz_dataOut_payload_0_2008 = (_zz_dataOut_payload_0_2007 ? _zz_dataOut_payload_0_1988 : _zz_dataOut_payload_0_1982);
  assign _zz_dataOut_payload_0_2009 = (_zz_dataOut_payload_0_2007 ? _zz_dataOut_payload_0_1982 : _zz_dataOut_payload_0_1988);
  assign _zz_dataOut_payload_0_2010 = (_zz_dataOut_payload_0_2005 < _zz_dataOut_payload_0_2008);
  assign _zz_dataOut_payload_0_2011 = (_zz_dataOut_payload_0_2006 < _zz_dataOut_payload_0_2009);
  assign _zz_dataOut_payload_0_2024 = (_zz_dataOut_payload_0_1264 < _zz_dataOut_payload_0_1271);
  assign _zz_dataOut_payload_0_2025 = (_zz_dataOut_payload_0_2024 ? _zz_dataOut_payload_0_1264 : _zz_dataOut_payload_0_1271);
  assign _zz_dataOut_payload_0_2026 = (_zz_dataOut_payload_0_2024 ? _zz_dataOut_payload_0_1271 : _zz_dataOut_payload_0_1264);
  assign _zz_dataOut_payload_0_2027 = (_zz_dataOut_payload_0_1265 < _zz_dataOut_payload_0_1270);
  assign _zz_dataOut_payload_0_2028 = (_zz_dataOut_payload_0_2027 ? _zz_dataOut_payload_0_1265 : _zz_dataOut_payload_0_1270);
  assign _zz_dataOut_payload_0_2029 = (_zz_dataOut_payload_0_2027 ? _zz_dataOut_payload_0_1270 : _zz_dataOut_payload_0_1265);
  assign _zz_dataOut_payload_0_2030 = (_zz_dataOut_payload_0_1266 < _zz_dataOut_payload_0_1269);
  assign _zz_dataOut_payload_0_2031 = (_zz_dataOut_payload_0_2030 ? _zz_dataOut_payload_0_1266 : _zz_dataOut_payload_0_1269);
  assign _zz_dataOut_payload_0_2032 = (_zz_dataOut_payload_0_2030 ? _zz_dataOut_payload_0_1269 : _zz_dataOut_payload_0_1266);
  assign _zz_dataOut_payload_0_2033 = (_zz_dataOut_payload_0_1267 < _zz_dataOut_payload_0_1268);
  assign _zz_dataOut_payload_0_2034 = (_zz_dataOut_payload_0_2033 ? _zz_dataOut_payload_0_1267 : _zz_dataOut_payload_0_1268);
  assign _zz_dataOut_payload_0_2035 = (_zz_dataOut_payload_0_2033 ? _zz_dataOut_payload_0_1268 : _zz_dataOut_payload_0_1267);
  assign _zz_dataOut_payload_0_2036 = (_zz_dataOut_payload_0_2025 < _zz_dataOut_payload_0_2031);
  assign _zz_dataOut_payload_0_2037 = (_zz_dataOut_payload_0_2036 ? _zz_dataOut_payload_0_2025 : _zz_dataOut_payload_0_2031);
  assign _zz_dataOut_payload_0_2038 = (_zz_dataOut_payload_0_2036 ? _zz_dataOut_payload_0_2031 : _zz_dataOut_payload_0_2025);
  assign _zz_dataOut_payload_0_2039 = (_zz_dataOut_payload_0_2028 < _zz_dataOut_payload_0_2034);
  assign _zz_dataOut_payload_0_2040 = (_zz_dataOut_payload_0_2039 ? _zz_dataOut_payload_0_2028 : _zz_dataOut_payload_0_2034);
  assign _zz_dataOut_payload_0_2041 = (_zz_dataOut_payload_0_2039 ? _zz_dataOut_payload_0_2034 : _zz_dataOut_payload_0_2028);
  assign _zz_dataOut_payload_0_2042 = (_zz_dataOut_payload_0_2037 < _zz_dataOut_payload_0_2040);
  assign _zz_dataOut_payload_0_2043 = (_zz_dataOut_payload_0_2038 < _zz_dataOut_payload_0_2041);
  assign _zz_dataOut_payload_0_2048 = (_zz_dataOut_payload_0_2035 < _zz_dataOut_payload_0_2029);
  assign _zz_dataOut_payload_0_2049 = (_zz_dataOut_payload_0_2048 ? _zz_dataOut_payload_0_2035 : _zz_dataOut_payload_0_2029);
  assign _zz_dataOut_payload_0_2050 = (_zz_dataOut_payload_0_2048 ? _zz_dataOut_payload_0_2029 : _zz_dataOut_payload_0_2035);
  assign _zz_dataOut_payload_0_2051 = (_zz_dataOut_payload_0_2032 < _zz_dataOut_payload_0_2026);
  assign _zz_dataOut_payload_0_2052 = (_zz_dataOut_payload_0_2051 ? _zz_dataOut_payload_0_2032 : _zz_dataOut_payload_0_2026);
  assign _zz_dataOut_payload_0_2053 = (_zz_dataOut_payload_0_2051 ? _zz_dataOut_payload_0_2026 : _zz_dataOut_payload_0_2032);
  assign _zz_dataOut_payload_0_2054 = (_zz_dataOut_payload_0_2049 < _zz_dataOut_payload_0_2052);
  assign _zz_dataOut_payload_0_2055 = (_zz_dataOut_payload_0_2050 < _zz_dataOut_payload_0_2053);
  assign _zz_dataOut_payload_0_2068 = (_zz_dataOut_payload_0_1272 < _zz_dataOut_payload_0_1279);
  assign _zz_dataOut_payload_0_2069 = (_zz_dataOut_payload_0_2068 ? _zz_dataOut_payload_0_1272 : _zz_dataOut_payload_0_1279);
  assign _zz_dataOut_payload_0_2070 = (_zz_dataOut_payload_0_2068 ? _zz_dataOut_payload_0_1279 : _zz_dataOut_payload_0_1272);
  assign _zz_dataOut_payload_0_2071 = (_zz_dataOut_payload_0_1273 < _zz_dataOut_payload_0_1278);
  assign _zz_dataOut_payload_0_2072 = (_zz_dataOut_payload_0_2071 ? _zz_dataOut_payload_0_1273 : _zz_dataOut_payload_0_1278);
  assign _zz_dataOut_payload_0_2073 = (_zz_dataOut_payload_0_2071 ? _zz_dataOut_payload_0_1278 : _zz_dataOut_payload_0_1273);
  assign _zz_dataOut_payload_0_2074 = (_zz_dataOut_payload_0_1274 < _zz_dataOut_payload_0_1277);
  assign _zz_dataOut_payload_0_2075 = (_zz_dataOut_payload_0_2074 ? _zz_dataOut_payload_0_1274 : _zz_dataOut_payload_0_1277);
  assign _zz_dataOut_payload_0_2076 = (_zz_dataOut_payload_0_2074 ? _zz_dataOut_payload_0_1277 : _zz_dataOut_payload_0_1274);
  assign _zz_dataOut_payload_0_2077 = (_zz_dataOut_payload_0_1275 < _zz_dataOut_payload_0_1276);
  assign _zz_dataOut_payload_0_2078 = (_zz_dataOut_payload_0_2077 ? _zz_dataOut_payload_0_1275 : _zz_dataOut_payload_0_1276);
  assign _zz_dataOut_payload_0_2079 = (_zz_dataOut_payload_0_2077 ? _zz_dataOut_payload_0_1276 : _zz_dataOut_payload_0_1275);
  assign _zz_dataOut_payload_0_2080 = (_zz_dataOut_payload_0_2069 < _zz_dataOut_payload_0_2075);
  assign _zz_dataOut_payload_0_2081 = (_zz_dataOut_payload_0_2080 ? _zz_dataOut_payload_0_2069 : _zz_dataOut_payload_0_2075);
  assign _zz_dataOut_payload_0_2082 = (_zz_dataOut_payload_0_2080 ? _zz_dataOut_payload_0_2075 : _zz_dataOut_payload_0_2069);
  assign _zz_dataOut_payload_0_2083 = (_zz_dataOut_payload_0_2072 < _zz_dataOut_payload_0_2078);
  assign _zz_dataOut_payload_0_2084 = (_zz_dataOut_payload_0_2083 ? _zz_dataOut_payload_0_2072 : _zz_dataOut_payload_0_2078);
  assign _zz_dataOut_payload_0_2085 = (_zz_dataOut_payload_0_2083 ? _zz_dataOut_payload_0_2078 : _zz_dataOut_payload_0_2072);
  assign _zz_dataOut_payload_0_2086 = (_zz_dataOut_payload_0_2081 < _zz_dataOut_payload_0_2084);
  assign _zz_dataOut_payload_0_2087 = (_zz_dataOut_payload_0_2082 < _zz_dataOut_payload_0_2085);
  assign _zz_dataOut_payload_0_2092 = (_zz_dataOut_payload_0_2079 < _zz_dataOut_payload_0_2073);
  assign _zz_dataOut_payload_0_2093 = (_zz_dataOut_payload_0_2092 ? _zz_dataOut_payload_0_2079 : _zz_dataOut_payload_0_2073);
  assign _zz_dataOut_payload_0_2094 = (_zz_dataOut_payload_0_2092 ? _zz_dataOut_payload_0_2073 : _zz_dataOut_payload_0_2079);
  assign _zz_dataOut_payload_0_2095 = (_zz_dataOut_payload_0_2076 < _zz_dataOut_payload_0_2070);
  assign _zz_dataOut_payload_0_2096 = (_zz_dataOut_payload_0_2095 ? _zz_dataOut_payload_0_2076 : _zz_dataOut_payload_0_2070);
  assign _zz_dataOut_payload_0_2097 = (_zz_dataOut_payload_0_2095 ? _zz_dataOut_payload_0_2070 : _zz_dataOut_payload_0_2076);
  assign _zz_dataOut_payload_0_2098 = (_zz_dataOut_payload_0_2093 < _zz_dataOut_payload_0_2096);
  assign _zz_dataOut_payload_0_2099 = (_zz_dataOut_payload_0_2094 < _zz_dataOut_payload_0_2097);
  assign _zz_dataOut_payload_0_2112 = (_zz_dataOut_payload_0_1280 < _zz_dataOut_payload_0_1287);
  assign _zz_dataOut_payload_0_2113 = (_zz_dataOut_payload_0_2112 ? _zz_dataOut_payload_0_1280 : _zz_dataOut_payload_0_1287);
  assign _zz_dataOut_payload_0_2114 = (_zz_dataOut_payload_0_2112 ? _zz_dataOut_payload_0_1287 : _zz_dataOut_payload_0_1280);
  assign _zz_dataOut_payload_0_2115 = (_zz_dataOut_payload_0_1281 < _zz_dataOut_payload_0_1286);
  assign _zz_dataOut_payload_0_2116 = (_zz_dataOut_payload_0_2115 ? _zz_dataOut_payload_0_1281 : _zz_dataOut_payload_0_1286);
  assign _zz_dataOut_payload_0_2117 = (_zz_dataOut_payload_0_2115 ? _zz_dataOut_payload_0_1286 : _zz_dataOut_payload_0_1281);
  assign _zz_dataOut_payload_0_2118 = (_zz_dataOut_payload_0_1282 < _zz_dataOut_payload_0_1285);
  assign _zz_dataOut_payload_0_2119 = (_zz_dataOut_payload_0_2118 ? _zz_dataOut_payload_0_1282 : _zz_dataOut_payload_0_1285);
  assign _zz_dataOut_payload_0_2120 = (_zz_dataOut_payload_0_2118 ? _zz_dataOut_payload_0_1285 : _zz_dataOut_payload_0_1282);
  assign _zz_dataOut_payload_0_2121 = (_zz_dataOut_payload_0_1283 < _zz_dataOut_payload_0_1284);
  assign _zz_dataOut_payload_0_2122 = (_zz_dataOut_payload_0_2121 ? _zz_dataOut_payload_0_1283 : _zz_dataOut_payload_0_1284);
  assign _zz_dataOut_payload_0_2123 = (_zz_dataOut_payload_0_2121 ? _zz_dataOut_payload_0_1284 : _zz_dataOut_payload_0_1283);
  assign _zz_dataOut_payload_0_2124 = (_zz_dataOut_payload_0_2113 < _zz_dataOut_payload_0_2119);
  assign _zz_dataOut_payload_0_2125 = (_zz_dataOut_payload_0_2124 ? _zz_dataOut_payload_0_2113 : _zz_dataOut_payload_0_2119);
  assign _zz_dataOut_payload_0_2126 = (_zz_dataOut_payload_0_2124 ? _zz_dataOut_payload_0_2119 : _zz_dataOut_payload_0_2113);
  assign _zz_dataOut_payload_0_2127 = (_zz_dataOut_payload_0_2116 < _zz_dataOut_payload_0_2122);
  assign _zz_dataOut_payload_0_2128 = (_zz_dataOut_payload_0_2127 ? _zz_dataOut_payload_0_2116 : _zz_dataOut_payload_0_2122);
  assign _zz_dataOut_payload_0_2129 = (_zz_dataOut_payload_0_2127 ? _zz_dataOut_payload_0_2122 : _zz_dataOut_payload_0_2116);
  assign _zz_dataOut_payload_0_2130 = (_zz_dataOut_payload_0_2125 < _zz_dataOut_payload_0_2128);
  assign _zz_dataOut_payload_0_2131 = (_zz_dataOut_payload_0_2126 < _zz_dataOut_payload_0_2129);
  assign _zz_dataOut_payload_0_2136 = (_zz_dataOut_payload_0_2123 < _zz_dataOut_payload_0_2117);
  assign _zz_dataOut_payload_0_2137 = (_zz_dataOut_payload_0_2136 ? _zz_dataOut_payload_0_2123 : _zz_dataOut_payload_0_2117);
  assign _zz_dataOut_payload_0_2138 = (_zz_dataOut_payload_0_2136 ? _zz_dataOut_payload_0_2117 : _zz_dataOut_payload_0_2123);
  assign _zz_dataOut_payload_0_2139 = (_zz_dataOut_payload_0_2120 < _zz_dataOut_payload_0_2114);
  assign _zz_dataOut_payload_0_2140 = (_zz_dataOut_payload_0_2139 ? _zz_dataOut_payload_0_2120 : _zz_dataOut_payload_0_2114);
  assign _zz_dataOut_payload_0_2141 = (_zz_dataOut_payload_0_2139 ? _zz_dataOut_payload_0_2114 : _zz_dataOut_payload_0_2120);
  assign _zz_dataOut_payload_0_2142 = (_zz_dataOut_payload_0_2137 < _zz_dataOut_payload_0_2140);
  assign _zz_dataOut_payload_0_2143 = (_zz_dataOut_payload_0_2138 < _zz_dataOut_payload_0_2141);
  assign _zz_dataOut_payload_0_2156 = (_zz_dataOut_payload_0_1288 < _zz_dataOut_payload_0_1295);
  assign _zz_dataOut_payload_0_2157 = (_zz_dataOut_payload_0_2156 ? _zz_dataOut_payload_0_1288 : _zz_dataOut_payload_0_1295);
  assign _zz_dataOut_payload_0_2158 = (_zz_dataOut_payload_0_2156 ? _zz_dataOut_payload_0_1295 : _zz_dataOut_payload_0_1288);
  assign _zz_dataOut_payload_0_2159 = (_zz_dataOut_payload_0_1289 < _zz_dataOut_payload_0_1294);
  assign _zz_dataOut_payload_0_2160 = (_zz_dataOut_payload_0_2159 ? _zz_dataOut_payload_0_1289 : _zz_dataOut_payload_0_1294);
  assign _zz_dataOut_payload_0_2161 = (_zz_dataOut_payload_0_2159 ? _zz_dataOut_payload_0_1294 : _zz_dataOut_payload_0_1289);
  assign _zz_dataOut_payload_0_2162 = (_zz_dataOut_payload_0_1290 < _zz_dataOut_payload_0_1293);
  assign _zz_dataOut_payload_0_2163 = (_zz_dataOut_payload_0_2162 ? _zz_dataOut_payload_0_1290 : _zz_dataOut_payload_0_1293);
  assign _zz_dataOut_payload_0_2164 = (_zz_dataOut_payload_0_2162 ? _zz_dataOut_payload_0_1293 : _zz_dataOut_payload_0_1290);
  assign _zz_dataOut_payload_0_2165 = (_zz_dataOut_payload_0_1291 < _zz_dataOut_payload_0_1292);
  assign _zz_dataOut_payload_0_2166 = (_zz_dataOut_payload_0_2165 ? _zz_dataOut_payload_0_1291 : _zz_dataOut_payload_0_1292);
  assign _zz_dataOut_payload_0_2167 = (_zz_dataOut_payload_0_2165 ? _zz_dataOut_payload_0_1292 : _zz_dataOut_payload_0_1291);
  assign _zz_dataOut_payload_0_2168 = (_zz_dataOut_payload_0_2157 < _zz_dataOut_payload_0_2163);
  assign _zz_dataOut_payload_0_2169 = (_zz_dataOut_payload_0_2168 ? _zz_dataOut_payload_0_2157 : _zz_dataOut_payload_0_2163);
  assign _zz_dataOut_payload_0_2170 = (_zz_dataOut_payload_0_2168 ? _zz_dataOut_payload_0_2163 : _zz_dataOut_payload_0_2157);
  assign _zz_dataOut_payload_0_2171 = (_zz_dataOut_payload_0_2160 < _zz_dataOut_payload_0_2166);
  assign _zz_dataOut_payload_0_2172 = (_zz_dataOut_payload_0_2171 ? _zz_dataOut_payload_0_2160 : _zz_dataOut_payload_0_2166);
  assign _zz_dataOut_payload_0_2173 = (_zz_dataOut_payload_0_2171 ? _zz_dataOut_payload_0_2166 : _zz_dataOut_payload_0_2160);
  assign _zz_dataOut_payload_0_2174 = (_zz_dataOut_payload_0_2169 < _zz_dataOut_payload_0_2172);
  assign _zz_dataOut_payload_0_2175 = (_zz_dataOut_payload_0_2170 < _zz_dataOut_payload_0_2173);
  assign _zz_dataOut_payload_0_2180 = (_zz_dataOut_payload_0_2167 < _zz_dataOut_payload_0_2161);
  assign _zz_dataOut_payload_0_2181 = (_zz_dataOut_payload_0_2180 ? _zz_dataOut_payload_0_2167 : _zz_dataOut_payload_0_2161);
  assign _zz_dataOut_payload_0_2182 = (_zz_dataOut_payload_0_2180 ? _zz_dataOut_payload_0_2161 : _zz_dataOut_payload_0_2167);
  assign _zz_dataOut_payload_0_2183 = (_zz_dataOut_payload_0_2164 < _zz_dataOut_payload_0_2158);
  assign _zz_dataOut_payload_0_2184 = (_zz_dataOut_payload_0_2183 ? _zz_dataOut_payload_0_2164 : _zz_dataOut_payload_0_2158);
  assign _zz_dataOut_payload_0_2185 = (_zz_dataOut_payload_0_2183 ? _zz_dataOut_payload_0_2158 : _zz_dataOut_payload_0_2164);
  assign _zz_dataOut_payload_0_2186 = (_zz_dataOut_payload_0_2181 < _zz_dataOut_payload_0_2184);
  assign _zz_dataOut_payload_0_2187 = (_zz_dataOut_payload_0_2182 < _zz_dataOut_payload_0_2185);
  assign _zz_dataOut_payload_0_2200 = (_zz_dataOut_payload_0_1296 < _zz_dataOut_payload_0_1303);
  assign _zz_dataOut_payload_0_2201 = (_zz_dataOut_payload_0_2200 ? _zz_dataOut_payload_0_1296 : _zz_dataOut_payload_0_1303);
  assign _zz_dataOut_payload_0_2202 = (_zz_dataOut_payload_0_2200 ? _zz_dataOut_payload_0_1303 : _zz_dataOut_payload_0_1296);
  assign _zz_dataOut_payload_0_2203 = (_zz_dataOut_payload_0_1297 < _zz_dataOut_payload_0_1302);
  assign _zz_dataOut_payload_0_2204 = (_zz_dataOut_payload_0_2203 ? _zz_dataOut_payload_0_1297 : _zz_dataOut_payload_0_1302);
  assign _zz_dataOut_payload_0_2205 = (_zz_dataOut_payload_0_2203 ? _zz_dataOut_payload_0_1302 : _zz_dataOut_payload_0_1297);
  assign _zz_dataOut_payload_0_2206 = (_zz_dataOut_payload_0_1298 < _zz_dataOut_payload_0_1301);
  assign _zz_dataOut_payload_0_2207 = (_zz_dataOut_payload_0_2206 ? _zz_dataOut_payload_0_1298 : _zz_dataOut_payload_0_1301);
  assign _zz_dataOut_payload_0_2208 = (_zz_dataOut_payload_0_2206 ? _zz_dataOut_payload_0_1301 : _zz_dataOut_payload_0_1298);
  assign _zz_dataOut_payload_0_2209 = (_zz_dataOut_payload_0_1299 < _zz_dataOut_payload_0_1300);
  assign _zz_dataOut_payload_0_2210 = (_zz_dataOut_payload_0_2209 ? _zz_dataOut_payload_0_1299 : _zz_dataOut_payload_0_1300);
  assign _zz_dataOut_payload_0_2211 = (_zz_dataOut_payload_0_2209 ? _zz_dataOut_payload_0_1300 : _zz_dataOut_payload_0_1299);
  assign _zz_dataOut_payload_0_2212 = (_zz_dataOut_payload_0_2201 < _zz_dataOut_payload_0_2207);
  assign _zz_dataOut_payload_0_2213 = (_zz_dataOut_payload_0_2212 ? _zz_dataOut_payload_0_2201 : _zz_dataOut_payload_0_2207);
  assign _zz_dataOut_payload_0_2214 = (_zz_dataOut_payload_0_2212 ? _zz_dataOut_payload_0_2207 : _zz_dataOut_payload_0_2201);
  assign _zz_dataOut_payload_0_2215 = (_zz_dataOut_payload_0_2204 < _zz_dataOut_payload_0_2210);
  assign _zz_dataOut_payload_0_2216 = (_zz_dataOut_payload_0_2215 ? _zz_dataOut_payload_0_2204 : _zz_dataOut_payload_0_2210);
  assign _zz_dataOut_payload_0_2217 = (_zz_dataOut_payload_0_2215 ? _zz_dataOut_payload_0_2210 : _zz_dataOut_payload_0_2204);
  assign _zz_dataOut_payload_0_2218 = (_zz_dataOut_payload_0_2213 < _zz_dataOut_payload_0_2216);
  assign _zz_dataOut_payload_0_2219 = (_zz_dataOut_payload_0_2214 < _zz_dataOut_payload_0_2217);
  assign _zz_dataOut_payload_0_2224 = (_zz_dataOut_payload_0_2211 < _zz_dataOut_payload_0_2205);
  assign _zz_dataOut_payload_0_2225 = (_zz_dataOut_payload_0_2224 ? _zz_dataOut_payload_0_2211 : _zz_dataOut_payload_0_2205);
  assign _zz_dataOut_payload_0_2226 = (_zz_dataOut_payload_0_2224 ? _zz_dataOut_payload_0_2205 : _zz_dataOut_payload_0_2211);
  assign _zz_dataOut_payload_0_2227 = (_zz_dataOut_payload_0_2208 < _zz_dataOut_payload_0_2202);
  assign _zz_dataOut_payload_0_2228 = (_zz_dataOut_payload_0_2227 ? _zz_dataOut_payload_0_2208 : _zz_dataOut_payload_0_2202);
  assign _zz_dataOut_payload_0_2229 = (_zz_dataOut_payload_0_2227 ? _zz_dataOut_payload_0_2202 : _zz_dataOut_payload_0_2208);
  assign _zz_dataOut_payload_0_2230 = (_zz_dataOut_payload_0_2225 < _zz_dataOut_payload_0_2228);
  assign _zz_dataOut_payload_0_2231 = (_zz_dataOut_payload_0_2226 < _zz_dataOut_payload_0_2229);
  assign _zz_dataOut_payload_0_2244 = (_zz_dataOut_payload_0_1304 < _zz_dataOut_payload_0_1311);
  assign _zz_dataOut_payload_0_2245 = (_zz_dataOut_payload_0_2244 ? _zz_dataOut_payload_0_1304 : _zz_dataOut_payload_0_1311);
  assign _zz_dataOut_payload_0_2246 = (_zz_dataOut_payload_0_2244 ? _zz_dataOut_payload_0_1311 : _zz_dataOut_payload_0_1304);
  assign _zz_dataOut_payload_0_2247 = (_zz_dataOut_payload_0_1305 < _zz_dataOut_payload_0_1310);
  assign _zz_dataOut_payload_0_2248 = (_zz_dataOut_payload_0_2247 ? _zz_dataOut_payload_0_1305 : _zz_dataOut_payload_0_1310);
  assign _zz_dataOut_payload_0_2249 = (_zz_dataOut_payload_0_2247 ? _zz_dataOut_payload_0_1310 : _zz_dataOut_payload_0_1305);
  assign _zz_dataOut_payload_0_2250 = (_zz_dataOut_payload_0_1306 < _zz_dataOut_payload_0_1309);
  assign _zz_dataOut_payload_0_2251 = (_zz_dataOut_payload_0_2250 ? _zz_dataOut_payload_0_1306 : _zz_dataOut_payload_0_1309);
  assign _zz_dataOut_payload_0_2252 = (_zz_dataOut_payload_0_2250 ? _zz_dataOut_payload_0_1309 : _zz_dataOut_payload_0_1306);
  assign _zz_dataOut_payload_0_2253 = (_zz_dataOut_payload_0_1307 < _zz_dataOut_payload_0_1308);
  assign _zz_dataOut_payload_0_2254 = (_zz_dataOut_payload_0_2253 ? _zz_dataOut_payload_0_1307 : _zz_dataOut_payload_0_1308);
  assign _zz_dataOut_payload_0_2255 = (_zz_dataOut_payload_0_2253 ? _zz_dataOut_payload_0_1308 : _zz_dataOut_payload_0_1307);
  assign _zz_dataOut_payload_0_2256 = (_zz_dataOut_payload_0_2245 < _zz_dataOut_payload_0_2251);
  assign _zz_dataOut_payload_0_2257 = (_zz_dataOut_payload_0_2256 ? _zz_dataOut_payload_0_2245 : _zz_dataOut_payload_0_2251);
  assign _zz_dataOut_payload_0_2258 = (_zz_dataOut_payload_0_2256 ? _zz_dataOut_payload_0_2251 : _zz_dataOut_payload_0_2245);
  assign _zz_dataOut_payload_0_2259 = (_zz_dataOut_payload_0_2248 < _zz_dataOut_payload_0_2254);
  assign _zz_dataOut_payload_0_2260 = (_zz_dataOut_payload_0_2259 ? _zz_dataOut_payload_0_2248 : _zz_dataOut_payload_0_2254);
  assign _zz_dataOut_payload_0_2261 = (_zz_dataOut_payload_0_2259 ? _zz_dataOut_payload_0_2254 : _zz_dataOut_payload_0_2248);
  assign _zz_dataOut_payload_0_2262 = (_zz_dataOut_payload_0_2257 < _zz_dataOut_payload_0_2260);
  assign _zz_dataOut_payload_0_2263 = (_zz_dataOut_payload_0_2258 < _zz_dataOut_payload_0_2261);
  assign _zz_dataOut_payload_0_2268 = (_zz_dataOut_payload_0_2255 < _zz_dataOut_payload_0_2249);
  assign _zz_dataOut_payload_0_2269 = (_zz_dataOut_payload_0_2268 ? _zz_dataOut_payload_0_2255 : _zz_dataOut_payload_0_2249);
  assign _zz_dataOut_payload_0_2270 = (_zz_dataOut_payload_0_2268 ? _zz_dataOut_payload_0_2249 : _zz_dataOut_payload_0_2255);
  assign _zz_dataOut_payload_0_2271 = (_zz_dataOut_payload_0_2252 < _zz_dataOut_payload_0_2246);
  assign _zz_dataOut_payload_0_2272 = (_zz_dataOut_payload_0_2271 ? _zz_dataOut_payload_0_2252 : _zz_dataOut_payload_0_2246);
  assign _zz_dataOut_payload_0_2273 = (_zz_dataOut_payload_0_2271 ? _zz_dataOut_payload_0_2246 : _zz_dataOut_payload_0_2252);
  assign _zz_dataOut_payload_0_2274 = (_zz_dataOut_payload_0_2269 < _zz_dataOut_payload_0_2272);
  assign _zz_dataOut_payload_0_2275 = (_zz_dataOut_payload_0_2270 < _zz_dataOut_payload_0_2273);
  assign _zz_dataOut_payload_0_2288 = (_zz_dataOut_payload_0_1312 < _zz_dataOut_payload_0_1319);
  assign _zz_dataOut_payload_0_2289 = (_zz_dataOut_payload_0_2288 ? _zz_dataOut_payload_0_1312 : _zz_dataOut_payload_0_1319);
  assign _zz_dataOut_payload_0_2290 = (_zz_dataOut_payload_0_2288 ? _zz_dataOut_payload_0_1319 : _zz_dataOut_payload_0_1312);
  assign _zz_dataOut_payload_0_2291 = (_zz_dataOut_payload_0_1313 < _zz_dataOut_payload_0_1318);
  assign _zz_dataOut_payload_0_2292 = (_zz_dataOut_payload_0_2291 ? _zz_dataOut_payload_0_1313 : _zz_dataOut_payload_0_1318);
  assign _zz_dataOut_payload_0_2293 = (_zz_dataOut_payload_0_2291 ? _zz_dataOut_payload_0_1318 : _zz_dataOut_payload_0_1313);
  assign _zz_dataOut_payload_0_2294 = (_zz_dataOut_payload_0_1314 < _zz_dataOut_payload_0_1317);
  assign _zz_dataOut_payload_0_2295 = (_zz_dataOut_payload_0_2294 ? _zz_dataOut_payload_0_1314 : _zz_dataOut_payload_0_1317);
  assign _zz_dataOut_payload_0_2296 = (_zz_dataOut_payload_0_2294 ? _zz_dataOut_payload_0_1317 : _zz_dataOut_payload_0_1314);
  assign _zz_dataOut_payload_0_2297 = (_zz_dataOut_payload_0_1315 < _zz_dataOut_payload_0_1316);
  assign _zz_dataOut_payload_0_2298 = (_zz_dataOut_payload_0_2297 ? _zz_dataOut_payload_0_1315 : _zz_dataOut_payload_0_1316);
  assign _zz_dataOut_payload_0_2299 = (_zz_dataOut_payload_0_2297 ? _zz_dataOut_payload_0_1316 : _zz_dataOut_payload_0_1315);
  assign _zz_dataOut_payload_0_2300 = (_zz_dataOut_payload_0_2289 < _zz_dataOut_payload_0_2295);
  assign _zz_dataOut_payload_0_2301 = (_zz_dataOut_payload_0_2300 ? _zz_dataOut_payload_0_2289 : _zz_dataOut_payload_0_2295);
  assign _zz_dataOut_payload_0_2302 = (_zz_dataOut_payload_0_2300 ? _zz_dataOut_payload_0_2295 : _zz_dataOut_payload_0_2289);
  assign _zz_dataOut_payload_0_2303 = (_zz_dataOut_payload_0_2292 < _zz_dataOut_payload_0_2298);
  assign _zz_dataOut_payload_0_2304 = (_zz_dataOut_payload_0_2303 ? _zz_dataOut_payload_0_2292 : _zz_dataOut_payload_0_2298);
  assign _zz_dataOut_payload_0_2305 = (_zz_dataOut_payload_0_2303 ? _zz_dataOut_payload_0_2298 : _zz_dataOut_payload_0_2292);
  assign _zz_dataOut_payload_0_2306 = (_zz_dataOut_payload_0_2301 < _zz_dataOut_payload_0_2304);
  assign _zz_dataOut_payload_0_2307 = (_zz_dataOut_payload_0_2302 < _zz_dataOut_payload_0_2305);
  assign _zz_dataOut_payload_0_2312 = (_zz_dataOut_payload_0_2299 < _zz_dataOut_payload_0_2293);
  assign _zz_dataOut_payload_0_2313 = (_zz_dataOut_payload_0_2312 ? _zz_dataOut_payload_0_2299 : _zz_dataOut_payload_0_2293);
  assign _zz_dataOut_payload_0_2314 = (_zz_dataOut_payload_0_2312 ? _zz_dataOut_payload_0_2293 : _zz_dataOut_payload_0_2299);
  assign _zz_dataOut_payload_0_2315 = (_zz_dataOut_payload_0_2296 < _zz_dataOut_payload_0_2290);
  assign _zz_dataOut_payload_0_2316 = (_zz_dataOut_payload_0_2315 ? _zz_dataOut_payload_0_2296 : _zz_dataOut_payload_0_2290);
  assign _zz_dataOut_payload_0_2317 = (_zz_dataOut_payload_0_2315 ? _zz_dataOut_payload_0_2290 : _zz_dataOut_payload_0_2296);
  assign _zz_dataOut_payload_0_2318 = (_zz_dataOut_payload_0_2313 < _zz_dataOut_payload_0_2316);
  assign _zz_dataOut_payload_0_2319 = (_zz_dataOut_payload_0_2314 < _zz_dataOut_payload_0_2317);
  assign _zz_dataOut_payload_0_2332 = (_zz_dataOut_payload_0_1320 < _zz_dataOut_payload_0_1327);
  assign _zz_dataOut_payload_0_2333 = (_zz_dataOut_payload_0_2332 ? _zz_dataOut_payload_0_1320 : _zz_dataOut_payload_0_1327);
  assign _zz_dataOut_payload_0_2334 = (_zz_dataOut_payload_0_2332 ? _zz_dataOut_payload_0_1327 : _zz_dataOut_payload_0_1320);
  assign _zz_dataOut_payload_0_2335 = (_zz_dataOut_payload_0_1321 < _zz_dataOut_payload_0_1326);
  assign _zz_dataOut_payload_0_2336 = (_zz_dataOut_payload_0_2335 ? _zz_dataOut_payload_0_1321 : _zz_dataOut_payload_0_1326);
  assign _zz_dataOut_payload_0_2337 = (_zz_dataOut_payload_0_2335 ? _zz_dataOut_payload_0_1326 : _zz_dataOut_payload_0_1321);
  assign _zz_dataOut_payload_0_2338 = (_zz_dataOut_payload_0_1322 < _zz_dataOut_payload_0_1325);
  assign _zz_dataOut_payload_0_2339 = (_zz_dataOut_payload_0_2338 ? _zz_dataOut_payload_0_1322 : _zz_dataOut_payload_0_1325);
  assign _zz_dataOut_payload_0_2340 = (_zz_dataOut_payload_0_2338 ? _zz_dataOut_payload_0_1325 : _zz_dataOut_payload_0_1322);
  assign _zz_dataOut_payload_0_2341 = (_zz_dataOut_payload_0_1323 < _zz_dataOut_payload_0_1324);
  assign _zz_dataOut_payload_0_2342 = (_zz_dataOut_payload_0_2341 ? _zz_dataOut_payload_0_1323 : _zz_dataOut_payload_0_1324);
  assign _zz_dataOut_payload_0_2343 = (_zz_dataOut_payload_0_2341 ? _zz_dataOut_payload_0_1324 : _zz_dataOut_payload_0_1323);
  assign _zz_dataOut_payload_0_2344 = (_zz_dataOut_payload_0_2333 < _zz_dataOut_payload_0_2339);
  assign _zz_dataOut_payload_0_2345 = (_zz_dataOut_payload_0_2344 ? _zz_dataOut_payload_0_2333 : _zz_dataOut_payload_0_2339);
  assign _zz_dataOut_payload_0_2346 = (_zz_dataOut_payload_0_2344 ? _zz_dataOut_payload_0_2339 : _zz_dataOut_payload_0_2333);
  assign _zz_dataOut_payload_0_2347 = (_zz_dataOut_payload_0_2336 < _zz_dataOut_payload_0_2342);
  assign _zz_dataOut_payload_0_2348 = (_zz_dataOut_payload_0_2347 ? _zz_dataOut_payload_0_2336 : _zz_dataOut_payload_0_2342);
  assign _zz_dataOut_payload_0_2349 = (_zz_dataOut_payload_0_2347 ? _zz_dataOut_payload_0_2342 : _zz_dataOut_payload_0_2336);
  assign _zz_dataOut_payload_0_2350 = (_zz_dataOut_payload_0_2345 < _zz_dataOut_payload_0_2348);
  assign _zz_dataOut_payload_0_2351 = (_zz_dataOut_payload_0_2346 < _zz_dataOut_payload_0_2349);
  assign _zz_dataOut_payload_0_2356 = (_zz_dataOut_payload_0_2343 < _zz_dataOut_payload_0_2337);
  assign _zz_dataOut_payload_0_2357 = (_zz_dataOut_payload_0_2356 ? _zz_dataOut_payload_0_2343 : _zz_dataOut_payload_0_2337);
  assign _zz_dataOut_payload_0_2358 = (_zz_dataOut_payload_0_2356 ? _zz_dataOut_payload_0_2337 : _zz_dataOut_payload_0_2343);
  assign _zz_dataOut_payload_0_2359 = (_zz_dataOut_payload_0_2340 < _zz_dataOut_payload_0_2334);
  assign _zz_dataOut_payload_0_2360 = (_zz_dataOut_payload_0_2359 ? _zz_dataOut_payload_0_2340 : _zz_dataOut_payload_0_2334);
  assign _zz_dataOut_payload_0_2361 = (_zz_dataOut_payload_0_2359 ? _zz_dataOut_payload_0_2334 : _zz_dataOut_payload_0_2340);
  assign _zz_dataOut_payload_0_2362 = (_zz_dataOut_payload_0_2357 < _zz_dataOut_payload_0_2360);
  assign _zz_dataOut_payload_0_2363 = (_zz_dataOut_payload_0_2358 < _zz_dataOut_payload_0_2361);
  assign _zz_dataOut_payload_0_2376 = (_zz_dataOut_payload_0_1328 < _zz_dataOut_payload_0_1335);
  assign _zz_dataOut_payload_0_2377 = (_zz_dataOut_payload_0_2376 ? _zz_dataOut_payload_0_1328 : _zz_dataOut_payload_0_1335);
  assign _zz_dataOut_payload_0_2378 = (_zz_dataOut_payload_0_2376 ? _zz_dataOut_payload_0_1335 : _zz_dataOut_payload_0_1328);
  assign _zz_dataOut_payload_0_2379 = (_zz_dataOut_payload_0_1329 < _zz_dataOut_payload_0_1334);
  assign _zz_dataOut_payload_0_2380 = (_zz_dataOut_payload_0_2379 ? _zz_dataOut_payload_0_1329 : _zz_dataOut_payload_0_1334);
  assign _zz_dataOut_payload_0_2381 = (_zz_dataOut_payload_0_2379 ? _zz_dataOut_payload_0_1334 : _zz_dataOut_payload_0_1329);
  assign _zz_dataOut_payload_0_2382 = (_zz_dataOut_payload_0_1330 < _zz_dataOut_payload_0_1333);
  assign _zz_dataOut_payload_0_2383 = (_zz_dataOut_payload_0_2382 ? _zz_dataOut_payload_0_1330 : _zz_dataOut_payload_0_1333);
  assign _zz_dataOut_payload_0_2384 = (_zz_dataOut_payload_0_2382 ? _zz_dataOut_payload_0_1333 : _zz_dataOut_payload_0_1330);
  assign _zz_dataOut_payload_0_2385 = (_zz_dataOut_payload_0_1331 < _zz_dataOut_payload_0_1332);
  assign _zz_dataOut_payload_0_2386 = (_zz_dataOut_payload_0_2385 ? _zz_dataOut_payload_0_1331 : _zz_dataOut_payload_0_1332);
  assign _zz_dataOut_payload_0_2387 = (_zz_dataOut_payload_0_2385 ? _zz_dataOut_payload_0_1332 : _zz_dataOut_payload_0_1331);
  assign _zz_dataOut_payload_0_2388 = (_zz_dataOut_payload_0_2377 < _zz_dataOut_payload_0_2383);
  assign _zz_dataOut_payload_0_2389 = (_zz_dataOut_payload_0_2388 ? _zz_dataOut_payload_0_2377 : _zz_dataOut_payload_0_2383);
  assign _zz_dataOut_payload_0_2390 = (_zz_dataOut_payload_0_2388 ? _zz_dataOut_payload_0_2383 : _zz_dataOut_payload_0_2377);
  assign _zz_dataOut_payload_0_2391 = (_zz_dataOut_payload_0_2380 < _zz_dataOut_payload_0_2386);
  assign _zz_dataOut_payload_0_2392 = (_zz_dataOut_payload_0_2391 ? _zz_dataOut_payload_0_2380 : _zz_dataOut_payload_0_2386);
  assign _zz_dataOut_payload_0_2393 = (_zz_dataOut_payload_0_2391 ? _zz_dataOut_payload_0_2386 : _zz_dataOut_payload_0_2380);
  assign _zz_dataOut_payload_0_2394 = (_zz_dataOut_payload_0_2389 < _zz_dataOut_payload_0_2392);
  assign _zz_dataOut_payload_0_2395 = (_zz_dataOut_payload_0_2390 < _zz_dataOut_payload_0_2393);
  assign _zz_dataOut_payload_0_2400 = (_zz_dataOut_payload_0_2387 < _zz_dataOut_payload_0_2381);
  assign _zz_dataOut_payload_0_2401 = (_zz_dataOut_payload_0_2400 ? _zz_dataOut_payload_0_2387 : _zz_dataOut_payload_0_2381);
  assign _zz_dataOut_payload_0_2402 = (_zz_dataOut_payload_0_2400 ? _zz_dataOut_payload_0_2381 : _zz_dataOut_payload_0_2387);
  assign _zz_dataOut_payload_0_2403 = (_zz_dataOut_payload_0_2384 < _zz_dataOut_payload_0_2378);
  assign _zz_dataOut_payload_0_2404 = (_zz_dataOut_payload_0_2403 ? _zz_dataOut_payload_0_2384 : _zz_dataOut_payload_0_2378);
  assign _zz_dataOut_payload_0_2405 = (_zz_dataOut_payload_0_2403 ? _zz_dataOut_payload_0_2378 : _zz_dataOut_payload_0_2384);
  assign _zz_dataOut_payload_0_2406 = (_zz_dataOut_payload_0_2401 < _zz_dataOut_payload_0_2404);
  assign _zz_dataOut_payload_0_2407 = (_zz_dataOut_payload_0_2402 < _zz_dataOut_payload_0_2405);
  assign _zz_dataOut_payload_0_2420 = (_zz_dataOut_payload_0_1336 < _zz_dataOut_payload_0_1343);
  assign _zz_dataOut_payload_0_2421 = (_zz_dataOut_payload_0_2420 ? _zz_dataOut_payload_0_1336 : _zz_dataOut_payload_0_1343);
  assign _zz_dataOut_payload_0_2422 = (_zz_dataOut_payload_0_2420 ? _zz_dataOut_payload_0_1343 : _zz_dataOut_payload_0_1336);
  assign _zz_dataOut_payload_0_2423 = (_zz_dataOut_payload_0_1337 < _zz_dataOut_payload_0_1342);
  assign _zz_dataOut_payload_0_2424 = (_zz_dataOut_payload_0_2423 ? _zz_dataOut_payload_0_1337 : _zz_dataOut_payload_0_1342);
  assign _zz_dataOut_payload_0_2425 = (_zz_dataOut_payload_0_2423 ? _zz_dataOut_payload_0_1342 : _zz_dataOut_payload_0_1337);
  assign _zz_dataOut_payload_0_2426 = (_zz_dataOut_payload_0_1338 < _zz_dataOut_payload_0_1341);
  assign _zz_dataOut_payload_0_2427 = (_zz_dataOut_payload_0_2426 ? _zz_dataOut_payload_0_1338 : _zz_dataOut_payload_0_1341);
  assign _zz_dataOut_payload_0_2428 = (_zz_dataOut_payload_0_2426 ? _zz_dataOut_payload_0_1341 : _zz_dataOut_payload_0_1338);
  assign _zz_dataOut_payload_0_2429 = (_zz_dataOut_payload_0_1339 < _zz_dataOut_payload_0_1340);
  assign _zz_dataOut_payload_0_2430 = (_zz_dataOut_payload_0_2429 ? _zz_dataOut_payload_0_1339 : _zz_dataOut_payload_0_1340);
  assign _zz_dataOut_payload_0_2431 = (_zz_dataOut_payload_0_2429 ? _zz_dataOut_payload_0_1340 : _zz_dataOut_payload_0_1339);
  assign _zz_dataOut_payload_0_2432 = (_zz_dataOut_payload_0_2421 < _zz_dataOut_payload_0_2427);
  assign _zz_dataOut_payload_0_2433 = (_zz_dataOut_payload_0_2432 ? _zz_dataOut_payload_0_2421 : _zz_dataOut_payload_0_2427);
  assign _zz_dataOut_payload_0_2434 = (_zz_dataOut_payload_0_2432 ? _zz_dataOut_payload_0_2427 : _zz_dataOut_payload_0_2421);
  assign _zz_dataOut_payload_0_2435 = (_zz_dataOut_payload_0_2424 < _zz_dataOut_payload_0_2430);
  assign _zz_dataOut_payload_0_2436 = (_zz_dataOut_payload_0_2435 ? _zz_dataOut_payload_0_2424 : _zz_dataOut_payload_0_2430);
  assign _zz_dataOut_payload_0_2437 = (_zz_dataOut_payload_0_2435 ? _zz_dataOut_payload_0_2430 : _zz_dataOut_payload_0_2424);
  assign _zz_dataOut_payload_0_2438 = (_zz_dataOut_payload_0_2433 < _zz_dataOut_payload_0_2436);
  assign _zz_dataOut_payload_0_2439 = (_zz_dataOut_payload_0_2434 < _zz_dataOut_payload_0_2437);
  assign _zz_dataOut_payload_0_2444 = (_zz_dataOut_payload_0_2431 < _zz_dataOut_payload_0_2425);
  assign _zz_dataOut_payload_0_2445 = (_zz_dataOut_payload_0_2444 ? _zz_dataOut_payload_0_2431 : _zz_dataOut_payload_0_2425);
  assign _zz_dataOut_payload_0_2446 = (_zz_dataOut_payload_0_2444 ? _zz_dataOut_payload_0_2425 : _zz_dataOut_payload_0_2431);
  assign _zz_dataOut_payload_0_2447 = (_zz_dataOut_payload_0_2428 < _zz_dataOut_payload_0_2422);
  assign _zz_dataOut_payload_0_2448 = (_zz_dataOut_payload_0_2447 ? _zz_dataOut_payload_0_2428 : _zz_dataOut_payload_0_2422);
  assign _zz_dataOut_payload_0_2449 = (_zz_dataOut_payload_0_2447 ? _zz_dataOut_payload_0_2422 : _zz_dataOut_payload_0_2428);
  assign _zz_dataOut_payload_0_2450 = (_zz_dataOut_payload_0_2445 < _zz_dataOut_payload_0_2448);
  assign _zz_dataOut_payload_0_2451 = (_zz_dataOut_payload_0_2446 < _zz_dataOut_payload_0_2449);
  assign _zz_dataOut_payload_0_2464 = (_zz_dataOut_payload_0_1344 < _zz_dataOut_payload_0_1351);
  assign _zz_dataOut_payload_0_2465 = (_zz_dataOut_payload_0_2464 ? _zz_dataOut_payload_0_1344 : _zz_dataOut_payload_0_1351);
  assign _zz_dataOut_payload_0_2466 = (_zz_dataOut_payload_0_2464 ? _zz_dataOut_payload_0_1351 : _zz_dataOut_payload_0_1344);
  assign _zz_dataOut_payload_0_2467 = (_zz_dataOut_payload_0_1345 < _zz_dataOut_payload_0_1350);
  assign _zz_dataOut_payload_0_2468 = (_zz_dataOut_payload_0_2467 ? _zz_dataOut_payload_0_1345 : _zz_dataOut_payload_0_1350);
  assign _zz_dataOut_payload_0_2469 = (_zz_dataOut_payload_0_2467 ? _zz_dataOut_payload_0_1350 : _zz_dataOut_payload_0_1345);
  assign _zz_dataOut_payload_0_2470 = (_zz_dataOut_payload_0_1346 < _zz_dataOut_payload_0_1349);
  assign _zz_dataOut_payload_0_2471 = (_zz_dataOut_payload_0_2470 ? _zz_dataOut_payload_0_1346 : _zz_dataOut_payload_0_1349);
  assign _zz_dataOut_payload_0_2472 = (_zz_dataOut_payload_0_2470 ? _zz_dataOut_payload_0_1349 : _zz_dataOut_payload_0_1346);
  assign _zz_dataOut_payload_0_2473 = (_zz_dataOut_payload_0_1347 < _zz_dataOut_payload_0_1348);
  assign _zz_dataOut_payload_0_2474 = (_zz_dataOut_payload_0_2473 ? _zz_dataOut_payload_0_1347 : _zz_dataOut_payload_0_1348);
  assign _zz_dataOut_payload_0_2475 = (_zz_dataOut_payload_0_2473 ? _zz_dataOut_payload_0_1348 : _zz_dataOut_payload_0_1347);
  assign _zz_dataOut_payload_0_2476 = (_zz_dataOut_payload_0_2465 < _zz_dataOut_payload_0_2471);
  assign _zz_dataOut_payload_0_2477 = (_zz_dataOut_payload_0_2476 ? _zz_dataOut_payload_0_2465 : _zz_dataOut_payload_0_2471);
  assign _zz_dataOut_payload_0_2478 = (_zz_dataOut_payload_0_2476 ? _zz_dataOut_payload_0_2471 : _zz_dataOut_payload_0_2465);
  assign _zz_dataOut_payload_0_2479 = (_zz_dataOut_payload_0_2468 < _zz_dataOut_payload_0_2474);
  assign _zz_dataOut_payload_0_2480 = (_zz_dataOut_payload_0_2479 ? _zz_dataOut_payload_0_2468 : _zz_dataOut_payload_0_2474);
  assign _zz_dataOut_payload_0_2481 = (_zz_dataOut_payload_0_2479 ? _zz_dataOut_payload_0_2474 : _zz_dataOut_payload_0_2468);
  assign _zz_dataOut_payload_0_2482 = (_zz_dataOut_payload_0_2477 < _zz_dataOut_payload_0_2480);
  assign _zz_dataOut_payload_0_2483 = (_zz_dataOut_payload_0_2478 < _zz_dataOut_payload_0_2481);
  assign _zz_dataOut_payload_0_2488 = (_zz_dataOut_payload_0_2475 < _zz_dataOut_payload_0_2469);
  assign _zz_dataOut_payload_0_2489 = (_zz_dataOut_payload_0_2488 ? _zz_dataOut_payload_0_2475 : _zz_dataOut_payload_0_2469);
  assign _zz_dataOut_payload_0_2490 = (_zz_dataOut_payload_0_2488 ? _zz_dataOut_payload_0_2469 : _zz_dataOut_payload_0_2475);
  assign _zz_dataOut_payload_0_2491 = (_zz_dataOut_payload_0_2472 < _zz_dataOut_payload_0_2466);
  assign _zz_dataOut_payload_0_2492 = (_zz_dataOut_payload_0_2491 ? _zz_dataOut_payload_0_2472 : _zz_dataOut_payload_0_2466);
  assign _zz_dataOut_payload_0_2493 = (_zz_dataOut_payload_0_2491 ? _zz_dataOut_payload_0_2466 : _zz_dataOut_payload_0_2472);
  assign _zz_dataOut_payload_0_2494 = (_zz_dataOut_payload_0_2489 < _zz_dataOut_payload_0_2492);
  assign _zz_dataOut_payload_0_2495 = (_zz_dataOut_payload_0_2490 < _zz_dataOut_payload_0_2493);
  assign _zz_dataOut_payload_0_2508 = (_zz_dataOut_payload_0_1352 < _zz_dataOut_payload_0_1359);
  assign _zz_dataOut_payload_0_2509 = (_zz_dataOut_payload_0_2508 ? _zz_dataOut_payload_0_1352 : _zz_dataOut_payload_0_1359);
  assign _zz_dataOut_payload_0_2510 = (_zz_dataOut_payload_0_2508 ? _zz_dataOut_payload_0_1359 : _zz_dataOut_payload_0_1352);
  assign _zz_dataOut_payload_0_2511 = (_zz_dataOut_payload_0_1353 < _zz_dataOut_payload_0_1358);
  assign _zz_dataOut_payload_0_2512 = (_zz_dataOut_payload_0_2511 ? _zz_dataOut_payload_0_1353 : _zz_dataOut_payload_0_1358);
  assign _zz_dataOut_payload_0_2513 = (_zz_dataOut_payload_0_2511 ? _zz_dataOut_payload_0_1358 : _zz_dataOut_payload_0_1353);
  assign _zz_dataOut_payload_0_2514 = (_zz_dataOut_payload_0_1354 < _zz_dataOut_payload_0_1357);
  assign _zz_dataOut_payload_0_2515 = (_zz_dataOut_payload_0_2514 ? _zz_dataOut_payload_0_1354 : _zz_dataOut_payload_0_1357);
  assign _zz_dataOut_payload_0_2516 = (_zz_dataOut_payload_0_2514 ? _zz_dataOut_payload_0_1357 : _zz_dataOut_payload_0_1354);
  assign _zz_dataOut_payload_0_2517 = (_zz_dataOut_payload_0_1355 < _zz_dataOut_payload_0_1356);
  assign _zz_dataOut_payload_0_2518 = (_zz_dataOut_payload_0_2517 ? _zz_dataOut_payload_0_1355 : _zz_dataOut_payload_0_1356);
  assign _zz_dataOut_payload_0_2519 = (_zz_dataOut_payload_0_2517 ? _zz_dataOut_payload_0_1356 : _zz_dataOut_payload_0_1355);
  assign _zz_dataOut_payload_0_2520 = (_zz_dataOut_payload_0_2509 < _zz_dataOut_payload_0_2515);
  assign _zz_dataOut_payload_0_2521 = (_zz_dataOut_payload_0_2520 ? _zz_dataOut_payload_0_2509 : _zz_dataOut_payload_0_2515);
  assign _zz_dataOut_payload_0_2522 = (_zz_dataOut_payload_0_2520 ? _zz_dataOut_payload_0_2515 : _zz_dataOut_payload_0_2509);
  assign _zz_dataOut_payload_0_2523 = (_zz_dataOut_payload_0_2512 < _zz_dataOut_payload_0_2518);
  assign _zz_dataOut_payload_0_2524 = (_zz_dataOut_payload_0_2523 ? _zz_dataOut_payload_0_2512 : _zz_dataOut_payload_0_2518);
  assign _zz_dataOut_payload_0_2525 = (_zz_dataOut_payload_0_2523 ? _zz_dataOut_payload_0_2518 : _zz_dataOut_payload_0_2512);
  assign _zz_dataOut_payload_0_2526 = (_zz_dataOut_payload_0_2521 < _zz_dataOut_payload_0_2524);
  assign _zz_dataOut_payload_0_2527 = (_zz_dataOut_payload_0_2522 < _zz_dataOut_payload_0_2525);
  assign _zz_dataOut_payload_0_2532 = (_zz_dataOut_payload_0_2519 < _zz_dataOut_payload_0_2513);
  assign _zz_dataOut_payload_0_2533 = (_zz_dataOut_payload_0_2532 ? _zz_dataOut_payload_0_2519 : _zz_dataOut_payload_0_2513);
  assign _zz_dataOut_payload_0_2534 = (_zz_dataOut_payload_0_2532 ? _zz_dataOut_payload_0_2513 : _zz_dataOut_payload_0_2519);
  assign _zz_dataOut_payload_0_2535 = (_zz_dataOut_payload_0_2516 < _zz_dataOut_payload_0_2510);
  assign _zz_dataOut_payload_0_2536 = (_zz_dataOut_payload_0_2535 ? _zz_dataOut_payload_0_2516 : _zz_dataOut_payload_0_2510);
  assign _zz_dataOut_payload_0_2537 = (_zz_dataOut_payload_0_2535 ? _zz_dataOut_payload_0_2510 : _zz_dataOut_payload_0_2516);
  assign _zz_dataOut_payload_0_2538 = (_zz_dataOut_payload_0_2533 < _zz_dataOut_payload_0_2536);
  assign _zz_dataOut_payload_0_2539 = (_zz_dataOut_payload_0_2534 < _zz_dataOut_payload_0_2537);
  assign _zz_dataOut_payload_0_2552 = (_zz_dataOut_payload_0_1360 < _zz_dataOut_payload_0_1367);
  assign _zz_dataOut_payload_0_2553 = (_zz_dataOut_payload_0_2552 ? _zz_dataOut_payload_0_1360 : _zz_dataOut_payload_0_1367);
  assign _zz_dataOut_payload_0_2554 = (_zz_dataOut_payload_0_2552 ? _zz_dataOut_payload_0_1367 : _zz_dataOut_payload_0_1360);
  assign _zz_dataOut_payload_0_2555 = (_zz_dataOut_payload_0_1361 < _zz_dataOut_payload_0_1366);
  assign _zz_dataOut_payload_0_2556 = (_zz_dataOut_payload_0_2555 ? _zz_dataOut_payload_0_1361 : _zz_dataOut_payload_0_1366);
  assign _zz_dataOut_payload_0_2557 = (_zz_dataOut_payload_0_2555 ? _zz_dataOut_payload_0_1366 : _zz_dataOut_payload_0_1361);
  assign _zz_dataOut_payload_0_2558 = (_zz_dataOut_payload_0_1362 < _zz_dataOut_payload_0_1365);
  assign _zz_dataOut_payload_0_2559 = (_zz_dataOut_payload_0_2558 ? _zz_dataOut_payload_0_1362 : _zz_dataOut_payload_0_1365);
  assign _zz_dataOut_payload_0_2560 = (_zz_dataOut_payload_0_2558 ? _zz_dataOut_payload_0_1365 : _zz_dataOut_payload_0_1362);
  assign _zz_dataOut_payload_0_2561 = (_zz_dataOut_payload_0_1363 < _zz_dataOut_payload_0_1364);
  assign _zz_dataOut_payload_0_2562 = (_zz_dataOut_payload_0_2561 ? _zz_dataOut_payload_0_1363 : _zz_dataOut_payload_0_1364);
  assign _zz_dataOut_payload_0_2563 = (_zz_dataOut_payload_0_2561 ? _zz_dataOut_payload_0_1364 : _zz_dataOut_payload_0_1363);
  assign _zz_dataOut_payload_0_2564 = (_zz_dataOut_payload_0_2553 < _zz_dataOut_payload_0_2559);
  assign _zz_dataOut_payload_0_2565 = (_zz_dataOut_payload_0_2564 ? _zz_dataOut_payload_0_2553 : _zz_dataOut_payload_0_2559);
  assign _zz_dataOut_payload_0_2566 = (_zz_dataOut_payload_0_2564 ? _zz_dataOut_payload_0_2559 : _zz_dataOut_payload_0_2553);
  assign _zz_dataOut_payload_0_2567 = (_zz_dataOut_payload_0_2556 < _zz_dataOut_payload_0_2562);
  assign _zz_dataOut_payload_0_2568 = (_zz_dataOut_payload_0_2567 ? _zz_dataOut_payload_0_2556 : _zz_dataOut_payload_0_2562);
  assign _zz_dataOut_payload_0_2569 = (_zz_dataOut_payload_0_2567 ? _zz_dataOut_payload_0_2562 : _zz_dataOut_payload_0_2556);
  assign _zz_dataOut_payload_0_2570 = (_zz_dataOut_payload_0_2565 < _zz_dataOut_payload_0_2568);
  assign _zz_dataOut_payload_0_2571 = (_zz_dataOut_payload_0_2566 < _zz_dataOut_payload_0_2569);
  assign _zz_dataOut_payload_0_2576 = (_zz_dataOut_payload_0_2563 < _zz_dataOut_payload_0_2557);
  assign _zz_dataOut_payload_0_2577 = (_zz_dataOut_payload_0_2576 ? _zz_dataOut_payload_0_2563 : _zz_dataOut_payload_0_2557);
  assign _zz_dataOut_payload_0_2578 = (_zz_dataOut_payload_0_2576 ? _zz_dataOut_payload_0_2557 : _zz_dataOut_payload_0_2563);
  assign _zz_dataOut_payload_0_2579 = (_zz_dataOut_payload_0_2560 < _zz_dataOut_payload_0_2554);
  assign _zz_dataOut_payload_0_2580 = (_zz_dataOut_payload_0_2579 ? _zz_dataOut_payload_0_2560 : _zz_dataOut_payload_0_2554);
  assign _zz_dataOut_payload_0_2581 = (_zz_dataOut_payload_0_2579 ? _zz_dataOut_payload_0_2554 : _zz_dataOut_payload_0_2560);
  assign _zz_dataOut_payload_0_2582 = (_zz_dataOut_payload_0_2577 < _zz_dataOut_payload_0_2580);
  assign _zz_dataOut_payload_0_2583 = (_zz_dataOut_payload_0_2578 < _zz_dataOut_payload_0_2581);
  assign _zz_dataOut_payload_0_2596 = (_zz_dataOut_payload_0_1368 < _zz_dataOut_payload_0_1375);
  assign _zz_dataOut_payload_0_2597 = (_zz_dataOut_payload_0_2596 ? _zz_dataOut_payload_0_1368 : _zz_dataOut_payload_0_1375);
  assign _zz_dataOut_payload_0_2598 = (_zz_dataOut_payload_0_2596 ? _zz_dataOut_payload_0_1375 : _zz_dataOut_payload_0_1368);
  assign _zz_dataOut_payload_0_2599 = (_zz_dataOut_payload_0_1369 < _zz_dataOut_payload_0_1374);
  assign _zz_dataOut_payload_0_2600 = (_zz_dataOut_payload_0_2599 ? _zz_dataOut_payload_0_1369 : _zz_dataOut_payload_0_1374);
  assign _zz_dataOut_payload_0_2601 = (_zz_dataOut_payload_0_2599 ? _zz_dataOut_payload_0_1374 : _zz_dataOut_payload_0_1369);
  assign _zz_dataOut_payload_0_2602 = (_zz_dataOut_payload_0_1370 < _zz_dataOut_payload_0_1373);
  assign _zz_dataOut_payload_0_2603 = (_zz_dataOut_payload_0_2602 ? _zz_dataOut_payload_0_1370 : _zz_dataOut_payload_0_1373);
  assign _zz_dataOut_payload_0_2604 = (_zz_dataOut_payload_0_2602 ? _zz_dataOut_payload_0_1373 : _zz_dataOut_payload_0_1370);
  assign _zz_dataOut_payload_0_2605 = (_zz_dataOut_payload_0_1371 < _zz_dataOut_payload_0_1372);
  assign _zz_dataOut_payload_0_2606 = (_zz_dataOut_payload_0_2605 ? _zz_dataOut_payload_0_1371 : _zz_dataOut_payload_0_1372);
  assign _zz_dataOut_payload_0_2607 = (_zz_dataOut_payload_0_2605 ? _zz_dataOut_payload_0_1372 : _zz_dataOut_payload_0_1371);
  assign _zz_dataOut_payload_0_2608 = (_zz_dataOut_payload_0_2597 < _zz_dataOut_payload_0_2603);
  assign _zz_dataOut_payload_0_2609 = (_zz_dataOut_payload_0_2608 ? _zz_dataOut_payload_0_2597 : _zz_dataOut_payload_0_2603);
  assign _zz_dataOut_payload_0_2610 = (_zz_dataOut_payload_0_2608 ? _zz_dataOut_payload_0_2603 : _zz_dataOut_payload_0_2597);
  assign _zz_dataOut_payload_0_2611 = (_zz_dataOut_payload_0_2600 < _zz_dataOut_payload_0_2606);
  assign _zz_dataOut_payload_0_2612 = (_zz_dataOut_payload_0_2611 ? _zz_dataOut_payload_0_2600 : _zz_dataOut_payload_0_2606);
  assign _zz_dataOut_payload_0_2613 = (_zz_dataOut_payload_0_2611 ? _zz_dataOut_payload_0_2606 : _zz_dataOut_payload_0_2600);
  assign _zz_dataOut_payload_0_2614 = (_zz_dataOut_payload_0_2609 < _zz_dataOut_payload_0_2612);
  assign _zz_dataOut_payload_0_2615 = (_zz_dataOut_payload_0_2610 < _zz_dataOut_payload_0_2613);
  assign _zz_dataOut_payload_0_2620 = (_zz_dataOut_payload_0_2607 < _zz_dataOut_payload_0_2601);
  assign _zz_dataOut_payload_0_2621 = (_zz_dataOut_payload_0_2620 ? _zz_dataOut_payload_0_2607 : _zz_dataOut_payload_0_2601);
  assign _zz_dataOut_payload_0_2622 = (_zz_dataOut_payload_0_2620 ? _zz_dataOut_payload_0_2601 : _zz_dataOut_payload_0_2607);
  assign _zz_dataOut_payload_0_2623 = (_zz_dataOut_payload_0_2604 < _zz_dataOut_payload_0_2598);
  assign _zz_dataOut_payload_0_2624 = (_zz_dataOut_payload_0_2623 ? _zz_dataOut_payload_0_2604 : _zz_dataOut_payload_0_2598);
  assign _zz_dataOut_payload_0_2625 = (_zz_dataOut_payload_0_2623 ? _zz_dataOut_payload_0_2598 : _zz_dataOut_payload_0_2604);
  assign _zz_dataOut_payload_0_2626 = (_zz_dataOut_payload_0_2621 < _zz_dataOut_payload_0_2624);
  assign _zz_dataOut_payload_0_2627 = (_zz_dataOut_payload_0_2622 < _zz_dataOut_payload_0_2625);
  assign _zz_dataOut_payload_0_2640 = (_zz_dataOut_payload_0_1376 < _zz_dataOut_payload_0_1383);
  assign _zz_dataOut_payload_0_2641 = (_zz_dataOut_payload_0_2640 ? _zz_dataOut_payload_0_1376 : _zz_dataOut_payload_0_1383);
  assign _zz_dataOut_payload_0_2642 = (_zz_dataOut_payload_0_2640 ? _zz_dataOut_payload_0_1383 : _zz_dataOut_payload_0_1376);
  assign _zz_dataOut_payload_0_2643 = (_zz_dataOut_payload_0_1377 < _zz_dataOut_payload_0_1382);
  assign _zz_dataOut_payload_0_2644 = (_zz_dataOut_payload_0_2643 ? _zz_dataOut_payload_0_1377 : _zz_dataOut_payload_0_1382);
  assign _zz_dataOut_payload_0_2645 = (_zz_dataOut_payload_0_2643 ? _zz_dataOut_payload_0_1382 : _zz_dataOut_payload_0_1377);
  assign _zz_dataOut_payload_0_2646 = (_zz_dataOut_payload_0_1378 < _zz_dataOut_payload_0_1381);
  assign _zz_dataOut_payload_0_2647 = (_zz_dataOut_payload_0_2646 ? _zz_dataOut_payload_0_1378 : _zz_dataOut_payload_0_1381);
  assign _zz_dataOut_payload_0_2648 = (_zz_dataOut_payload_0_2646 ? _zz_dataOut_payload_0_1381 : _zz_dataOut_payload_0_1378);
  assign _zz_dataOut_payload_0_2649 = (_zz_dataOut_payload_0_1379 < _zz_dataOut_payload_0_1380);
  assign _zz_dataOut_payload_0_2650 = (_zz_dataOut_payload_0_2649 ? _zz_dataOut_payload_0_1379 : _zz_dataOut_payload_0_1380);
  assign _zz_dataOut_payload_0_2651 = (_zz_dataOut_payload_0_2649 ? _zz_dataOut_payload_0_1380 : _zz_dataOut_payload_0_1379);
  assign _zz_dataOut_payload_0_2652 = (_zz_dataOut_payload_0_2641 < _zz_dataOut_payload_0_2647);
  assign _zz_dataOut_payload_0_2653 = (_zz_dataOut_payload_0_2652 ? _zz_dataOut_payload_0_2641 : _zz_dataOut_payload_0_2647);
  assign _zz_dataOut_payload_0_2654 = (_zz_dataOut_payload_0_2652 ? _zz_dataOut_payload_0_2647 : _zz_dataOut_payload_0_2641);
  assign _zz_dataOut_payload_0_2655 = (_zz_dataOut_payload_0_2644 < _zz_dataOut_payload_0_2650);
  assign _zz_dataOut_payload_0_2656 = (_zz_dataOut_payload_0_2655 ? _zz_dataOut_payload_0_2644 : _zz_dataOut_payload_0_2650);
  assign _zz_dataOut_payload_0_2657 = (_zz_dataOut_payload_0_2655 ? _zz_dataOut_payload_0_2650 : _zz_dataOut_payload_0_2644);
  assign _zz_dataOut_payload_0_2658 = (_zz_dataOut_payload_0_2653 < _zz_dataOut_payload_0_2656);
  assign _zz_dataOut_payload_0_2659 = (_zz_dataOut_payload_0_2654 < _zz_dataOut_payload_0_2657);
  assign _zz_dataOut_payload_0_2664 = (_zz_dataOut_payload_0_2651 < _zz_dataOut_payload_0_2645);
  assign _zz_dataOut_payload_0_2665 = (_zz_dataOut_payload_0_2664 ? _zz_dataOut_payload_0_2651 : _zz_dataOut_payload_0_2645);
  assign _zz_dataOut_payload_0_2666 = (_zz_dataOut_payload_0_2664 ? _zz_dataOut_payload_0_2645 : _zz_dataOut_payload_0_2651);
  assign _zz_dataOut_payload_0_2667 = (_zz_dataOut_payload_0_2648 < _zz_dataOut_payload_0_2642);
  assign _zz_dataOut_payload_0_2668 = (_zz_dataOut_payload_0_2667 ? _zz_dataOut_payload_0_2648 : _zz_dataOut_payload_0_2642);
  assign _zz_dataOut_payload_0_2669 = (_zz_dataOut_payload_0_2667 ? _zz_dataOut_payload_0_2642 : _zz_dataOut_payload_0_2648);
  assign _zz_dataOut_payload_0_2670 = (_zz_dataOut_payload_0_2665 < _zz_dataOut_payload_0_2668);
  assign _zz_dataOut_payload_0_2671 = (_zz_dataOut_payload_0_2666 < _zz_dataOut_payload_0_2669);
  assign _zz_dataOut_payload_0_2684 = (_zz_dataOut_payload_0_1384 < _zz_dataOut_payload_0_1391);
  assign _zz_dataOut_payload_0_2685 = (_zz_dataOut_payload_0_2684 ? _zz_dataOut_payload_0_1384 : _zz_dataOut_payload_0_1391);
  assign _zz_dataOut_payload_0_2686 = (_zz_dataOut_payload_0_2684 ? _zz_dataOut_payload_0_1391 : _zz_dataOut_payload_0_1384);
  assign _zz_dataOut_payload_0_2687 = (_zz_dataOut_payload_0_1385 < _zz_dataOut_payload_0_1390);
  assign _zz_dataOut_payload_0_2688 = (_zz_dataOut_payload_0_2687 ? _zz_dataOut_payload_0_1385 : _zz_dataOut_payload_0_1390);
  assign _zz_dataOut_payload_0_2689 = (_zz_dataOut_payload_0_2687 ? _zz_dataOut_payload_0_1390 : _zz_dataOut_payload_0_1385);
  assign _zz_dataOut_payload_0_2690 = (_zz_dataOut_payload_0_1386 < _zz_dataOut_payload_0_1389);
  assign _zz_dataOut_payload_0_2691 = (_zz_dataOut_payload_0_2690 ? _zz_dataOut_payload_0_1386 : _zz_dataOut_payload_0_1389);
  assign _zz_dataOut_payload_0_2692 = (_zz_dataOut_payload_0_2690 ? _zz_dataOut_payload_0_1389 : _zz_dataOut_payload_0_1386);
  assign _zz_dataOut_payload_0_2693 = (_zz_dataOut_payload_0_1387 < _zz_dataOut_payload_0_1388);
  assign _zz_dataOut_payload_0_2694 = (_zz_dataOut_payload_0_2693 ? _zz_dataOut_payload_0_1387 : _zz_dataOut_payload_0_1388);
  assign _zz_dataOut_payload_0_2695 = (_zz_dataOut_payload_0_2693 ? _zz_dataOut_payload_0_1388 : _zz_dataOut_payload_0_1387);
  assign _zz_dataOut_payload_0_2696 = (_zz_dataOut_payload_0_2685 < _zz_dataOut_payload_0_2691);
  assign _zz_dataOut_payload_0_2697 = (_zz_dataOut_payload_0_2696 ? _zz_dataOut_payload_0_2685 : _zz_dataOut_payload_0_2691);
  assign _zz_dataOut_payload_0_2698 = (_zz_dataOut_payload_0_2696 ? _zz_dataOut_payload_0_2691 : _zz_dataOut_payload_0_2685);
  assign _zz_dataOut_payload_0_2699 = (_zz_dataOut_payload_0_2688 < _zz_dataOut_payload_0_2694);
  assign _zz_dataOut_payload_0_2700 = (_zz_dataOut_payload_0_2699 ? _zz_dataOut_payload_0_2688 : _zz_dataOut_payload_0_2694);
  assign _zz_dataOut_payload_0_2701 = (_zz_dataOut_payload_0_2699 ? _zz_dataOut_payload_0_2694 : _zz_dataOut_payload_0_2688);
  assign _zz_dataOut_payload_0_2702 = (_zz_dataOut_payload_0_2697 < _zz_dataOut_payload_0_2700);
  assign _zz_dataOut_payload_0_2703 = (_zz_dataOut_payload_0_2698 < _zz_dataOut_payload_0_2701);
  assign _zz_dataOut_payload_0_2708 = (_zz_dataOut_payload_0_2695 < _zz_dataOut_payload_0_2689);
  assign _zz_dataOut_payload_0_2709 = (_zz_dataOut_payload_0_2708 ? _zz_dataOut_payload_0_2695 : _zz_dataOut_payload_0_2689);
  assign _zz_dataOut_payload_0_2710 = (_zz_dataOut_payload_0_2708 ? _zz_dataOut_payload_0_2689 : _zz_dataOut_payload_0_2695);
  assign _zz_dataOut_payload_0_2711 = (_zz_dataOut_payload_0_2692 < _zz_dataOut_payload_0_2686);
  assign _zz_dataOut_payload_0_2712 = (_zz_dataOut_payload_0_2711 ? _zz_dataOut_payload_0_2692 : _zz_dataOut_payload_0_2686);
  assign _zz_dataOut_payload_0_2713 = (_zz_dataOut_payload_0_2711 ? _zz_dataOut_payload_0_2686 : _zz_dataOut_payload_0_2692);
  assign _zz_dataOut_payload_0_2714 = (_zz_dataOut_payload_0_2709 < _zz_dataOut_payload_0_2712);
  assign _zz_dataOut_payload_0_2715 = (_zz_dataOut_payload_0_2710 < _zz_dataOut_payload_0_2713);
  assign _zz_dataOut_payload_0_2728 = (_zz_dataOut_payload_0_1392 < _zz_dataOut_payload_0_1399);
  assign _zz_dataOut_payload_0_2729 = (_zz_dataOut_payload_0_2728 ? _zz_dataOut_payload_0_1392 : _zz_dataOut_payload_0_1399);
  assign _zz_dataOut_payload_0_2730 = (_zz_dataOut_payload_0_2728 ? _zz_dataOut_payload_0_1399 : _zz_dataOut_payload_0_1392);
  assign _zz_dataOut_payload_0_2731 = (_zz_dataOut_payload_0_1393 < _zz_dataOut_payload_0_1398);
  assign _zz_dataOut_payload_0_2732 = (_zz_dataOut_payload_0_2731 ? _zz_dataOut_payload_0_1393 : _zz_dataOut_payload_0_1398);
  assign _zz_dataOut_payload_0_2733 = (_zz_dataOut_payload_0_2731 ? _zz_dataOut_payload_0_1398 : _zz_dataOut_payload_0_1393);
  assign _zz_dataOut_payload_0_2734 = (_zz_dataOut_payload_0_1394 < _zz_dataOut_payload_0_1397);
  assign _zz_dataOut_payload_0_2735 = (_zz_dataOut_payload_0_2734 ? _zz_dataOut_payload_0_1394 : _zz_dataOut_payload_0_1397);
  assign _zz_dataOut_payload_0_2736 = (_zz_dataOut_payload_0_2734 ? _zz_dataOut_payload_0_1397 : _zz_dataOut_payload_0_1394);
  assign _zz_dataOut_payload_0_2737 = (_zz_dataOut_payload_0_1395 < _zz_dataOut_payload_0_1396);
  assign _zz_dataOut_payload_0_2738 = (_zz_dataOut_payload_0_2737 ? _zz_dataOut_payload_0_1395 : _zz_dataOut_payload_0_1396);
  assign _zz_dataOut_payload_0_2739 = (_zz_dataOut_payload_0_2737 ? _zz_dataOut_payload_0_1396 : _zz_dataOut_payload_0_1395);
  assign _zz_dataOut_payload_0_2740 = (_zz_dataOut_payload_0_2729 < _zz_dataOut_payload_0_2735);
  assign _zz_dataOut_payload_0_2741 = (_zz_dataOut_payload_0_2740 ? _zz_dataOut_payload_0_2729 : _zz_dataOut_payload_0_2735);
  assign _zz_dataOut_payload_0_2742 = (_zz_dataOut_payload_0_2740 ? _zz_dataOut_payload_0_2735 : _zz_dataOut_payload_0_2729);
  assign _zz_dataOut_payload_0_2743 = (_zz_dataOut_payload_0_2732 < _zz_dataOut_payload_0_2738);
  assign _zz_dataOut_payload_0_2744 = (_zz_dataOut_payload_0_2743 ? _zz_dataOut_payload_0_2732 : _zz_dataOut_payload_0_2738);
  assign _zz_dataOut_payload_0_2745 = (_zz_dataOut_payload_0_2743 ? _zz_dataOut_payload_0_2738 : _zz_dataOut_payload_0_2732);
  assign _zz_dataOut_payload_0_2746 = (_zz_dataOut_payload_0_2741 < _zz_dataOut_payload_0_2744);
  assign _zz_dataOut_payload_0_2747 = (_zz_dataOut_payload_0_2742 < _zz_dataOut_payload_0_2745);
  assign _zz_dataOut_payload_0_2752 = (_zz_dataOut_payload_0_2739 < _zz_dataOut_payload_0_2733);
  assign _zz_dataOut_payload_0_2753 = (_zz_dataOut_payload_0_2752 ? _zz_dataOut_payload_0_2739 : _zz_dataOut_payload_0_2733);
  assign _zz_dataOut_payload_0_2754 = (_zz_dataOut_payload_0_2752 ? _zz_dataOut_payload_0_2733 : _zz_dataOut_payload_0_2739);
  assign _zz_dataOut_payload_0_2755 = (_zz_dataOut_payload_0_2736 < _zz_dataOut_payload_0_2730);
  assign _zz_dataOut_payload_0_2756 = (_zz_dataOut_payload_0_2755 ? _zz_dataOut_payload_0_2736 : _zz_dataOut_payload_0_2730);
  assign _zz_dataOut_payload_0_2757 = (_zz_dataOut_payload_0_2755 ? _zz_dataOut_payload_0_2730 : _zz_dataOut_payload_0_2736);
  assign _zz_dataOut_payload_0_2758 = (_zz_dataOut_payload_0_2753 < _zz_dataOut_payload_0_2756);
  assign _zz_dataOut_payload_0_2759 = (_zz_dataOut_payload_0_2754 < _zz_dataOut_payload_0_2757);
  assign _zz_dataOut_payload_0_2772 = (_zz_dataOut_payload_0_1400 < _zz_dataOut_payload_0_1407);
  assign _zz_dataOut_payload_0_2773 = (_zz_dataOut_payload_0_2772 ? _zz_dataOut_payload_0_1400 : _zz_dataOut_payload_0_1407);
  assign _zz_dataOut_payload_0_2774 = (_zz_dataOut_payload_0_2772 ? _zz_dataOut_payload_0_1407 : _zz_dataOut_payload_0_1400);
  assign _zz_dataOut_payload_0_2775 = (_zz_dataOut_payload_0_1401 < _zz_dataOut_payload_0_1406);
  assign _zz_dataOut_payload_0_2776 = (_zz_dataOut_payload_0_2775 ? _zz_dataOut_payload_0_1401 : _zz_dataOut_payload_0_1406);
  assign _zz_dataOut_payload_0_2777 = (_zz_dataOut_payload_0_2775 ? _zz_dataOut_payload_0_1406 : _zz_dataOut_payload_0_1401);
  assign _zz_dataOut_payload_0_2778 = (_zz_dataOut_payload_0_1402 < _zz_dataOut_payload_0_1405);
  assign _zz_dataOut_payload_0_2779 = (_zz_dataOut_payload_0_2778 ? _zz_dataOut_payload_0_1402 : _zz_dataOut_payload_0_1405);
  assign _zz_dataOut_payload_0_2780 = (_zz_dataOut_payload_0_2778 ? _zz_dataOut_payload_0_1405 : _zz_dataOut_payload_0_1402);
  assign _zz_dataOut_payload_0_2781 = (_zz_dataOut_payload_0_1403 < _zz_dataOut_payload_0_1404);
  assign _zz_dataOut_payload_0_2782 = (_zz_dataOut_payload_0_2781 ? _zz_dataOut_payload_0_1403 : _zz_dataOut_payload_0_1404);
  assign _zz_dataOut_payload_0_2783 = (_zz_dataOut_payload_0_2781 ? _zz_dataOut_payload_0_1404 : _zz_dataOut_payload_0_1403);
  assign _zz_dataOut_payload_0_2784 = (_zz_dataOut_payload_0_2773 < _zz_dataOut_payload_0_2779);
  assign _zz_dataOut_payload_0_2785 = (_zz_dataOut_payload_0_2784 ? _zz_dataOut_payload_0_2773 : _zz_dataOut_payload_0_2779);
  assign _zz_dataOut_payload_0_2786 = (_zz_dataOut_payload_0_2784 ? _zz_dataOut_payload_0_2779 : _zz_dataOut_payload_0_2773);
  assign _zz_dataOut_payload_0_2787 = (_zz_dataOut_payload_0_2776 < _zz_dataOut_payload_0_2782);
  assign _zz_dataOut_payload_0_2788 = (_zz_dataOut_payload_0_2787 ? _zz_dataOut_payload_0_2776 : _zz_dataOut_payload_0_2782);
  assign _zz_dataOut_payload_0_2789 = (_zz_dataOut_payload_0_2787 ? _zz_dataOut_payload_0_2782 : _zz_dataOut_payload_0_2776);
  assign _zz_dataOut_payload_0_2790 = (_zz_dataOut_payload_0_2785 < _zz_dataOut_payload_0_2788);
  assign _zz_dataOut_payload_0_2791 = (_zz_dataOut_payload_0_2786 < _zz_dataOut_payload_0_2789);
  assign _zz_dataOut_payload_0_2796 = (_zz_dataOut_payload_0_2783 < _zz_dataOut_payload_0_2777);
  assign _zz_dataOut_payload_0_2797 = (_zz_dataOut_payload_0_2796 ? _zz_dataOut_payload_0_2783 : _zz_dataOut_payload_0_2777);
  assign _zz_dataOut_payload_0_2798 = (_zz_dataOut_payload_0_2796 ? _zz_dataOut_payload_0_2777 : _zz_dataOut_payload_0_2783);
  assign _zz_dataOut_payload_0_2799 = (_zz_dataOut_payload_0_2780 < _zz_dataOut_payload_0_2774);
  assign _zz_dataOut_payload_0_2800 = (_zz_dataOut_payload_0_2799 ? _zz_dataOut_payload_0_2780 : _zz_dataOut_payload_0_2774);
  assign _zz_dataOut_payload_0_2801 = (_zz_dataOut_payload_0_2799 ? _zz_dataOut_payload_0_2774 : _zz_dataOut_payload_0_2780);
  assign _zz_dataOut_payload_0_2802 = (_zz_dataOut_payload_0_2797 < _zz_dataOut_payload_0_2800);
  assign _zz_dataOut_payload_0_2803 = (_zz_dataOut_payload_0_2798 < _zz_dataOut_payload_0_2801);
  assign _zz_dataOut_payload_0_3072 = (_zz_dataOut_payload_0_2816 < _zz_dataOut_payload_0_2831);
  assign _zz_dataOut_payload_0_3073 = (_zz_dataOut_payload_0_3072 ? _zz_dataOut_payload_0_2816 : _zz_dataOut_payload_0_2831);
  assign _zz_dataOut_payload_0_3074 = (_zz_dataOut_payload_0_3072 ? _zz_dataOut_payload_0_2831 : _zz_dataOut_payload_0_2816);
  assign _zz_dataOut_payload_0_3075 = (_zz_dataOut_payload_0_2817 < _zz_dataOut_payload_0_2830);
  assign _zz_dataOut_payload_0_3076 = (_zz_dataOut_payload_0_3075 ? _zz_dataOut_payload_0_2817 : _zz_dataOut_payload_0_2830);
  assign _zz_dataOut_payload_0_3077 = (_zz_dataOut_payload_0_3075 ? _zz_dataOut_payload_0_2830 : _zz_dataOut_payload_0_2817);
  assign _zz_dataOut_payload_0_3078 = (_zz_dataOut_payload_0_2818 < _zz_dataOut_payload_0_2829);
  assign _zz_dataOut_payload_0_3079 = (_zz_dataOut_payload_0_3078 ? _zz_dataOut_payload_0_2818 : _zz_dataOut_payload_0_2829);
  assign _zz_dataOut_payload_0_3080 = (_zz_dataOut_payload_0_3078 ? _zz_dataOut_payload_0_2829 : _zz_dataOut_payload_0_2818);
  assign _zz_dataOut_payload_0_3081 = (_zz_dataOut_payload_0_2819 < _zz_dataOut_payload_0_2828);
  assign _zz_dataOut_payload_0_3082 = (_zz_dataOut_payload_0_3081 ? _zz_dataOut_payload_0_2819 : _zz_dataOut_payload_0_2828);
  assign _zz_dataOut_payload_0_3083 = (_zz_dataOut_payload_0_3081 ? _zz_dataOut_payload_0_2828 : _zz_dataOut_payload_0_2819);
  assign _zz_dataOut_payload_0_3084 = (_zz_dataOut_payload_0_2820 < _zz_dataOut_payload_0_2827);
  assign _zz_dataOut_payload_0_3085 = (_zz_dataOut_payload_0_3084 ? _zz_dataOut_payload_0_2820 : _zz_dataOut_payload_0_2827);
  assign _zz_dataOut_payload_0_3086 = (_zz_dataOut_payload_0_3084 ? _zz_dataOut_payload_0_2827 : _zz_dataOut_payload_0_2820);
  assign _zz_dataOut_payload_0_3087 = (_zz_dataOut_payload_0_2821 < _zz_dataOut_payload_0_2826);
  assign _zz_dataOut_payload_0_3088 = (_zz_dataOut_payload_0_3087 ? _zz_dataOut_payload_0_2821 : _zz_dataOut_payload_0_2826);
  assign _zz_dataOut_payload_0_3089 = (_zz_dataOut_payload_0_3087 ? _zz_dataOut_payload_0_2826 : _zz_dataOut_payload_0_2821);
  assign _zz_dataOut_payload_0_3090 = (_zz_dataOut_payload_0_2822 < _zz_dataOut_payload_0_2825);
  assign _zz_dataOut_payload_0_3091 = (_zz_dataOut_payload_0_3090 ? _zz_dataOut_payload_0_2822 : _zz_dataOut_payload_0_2825);
  assign _zz_dataOut_payload_0_3092 = (_zz_dataOut_payload_0_3090 ? _zz_dataOut_payload_0_2825 : _zz_dataOut_payload_0_2822);
  assign _zz_dataOut_payload_0_3093 = (_zz_dataOut_payload_0_2823 < _zz_dataOut_payload_0_2824);
  assign _zz_dataOut_payload_0_3094 = (_zz_dataOut_payload_0_3093 ? _zz_dataOut_payload_0_2823 : _zz_dataOut_payload_0_2824);
  assign _zz_dataOut_payload_0_3095 = (_zz_dataOut_payload_0_3093 ? _zz_dataOut_payload_0_2824 : _zz_dataOut_payload_0_2823);
  assign _zz_dataOut_payload_0_3096 = (_zz_dataOut_payload_0_3073 < _zz_dataOut_payload_0_3085);
  assign _zz_dataOut_payload_0_3097 = (_zz_dataOut_payload_0_3096 ? _zz_dataOut_payload_0_3073 : _zz_dataOut_payload_0_3085);
  assign _zz_dataOut_payload_0_3098 = (_zz_dataOut_payload_0_3096 ? _zz_dataOut_payload_0_3085 : _zz_dataOut_payload_0_3073);
  assign _zz_dataOut_payload_0_3099 = (_zz_dataOut_payload_0_3076 < _zz_dataOut_payload_0_3088);
  assign _zz_dataOut_payload_0_3100 = (_zz_dataOut_payload_0_3099 ? _zz_dataOut_payload_0_3076 : _zz_dataOut_payload_0_3088);
  assign _zz_dataOut_payload_0_3101 = (_zz_dataOut_payload_0_3099 ? _zz_dataOut_payload_0_3088 : _zz_dataOut_payload_0_3076);
  assign _zz_dataOut_payload_0_3102 = (_zz_dataOut_payload_0_3079 < _zz_dataOut_payload_0_3091);
  assign _zz_dataOut_payload_0_3103 = (_zz_dataOut_payload_0_3102 ? _zz_dataOut_payload_0_3079 : _zz_dataOut_payload_0_3091);
  assign _zz_dataOut_payload_0_3104 = (_zz_dataOut_payload_0_3102 ? _zz_dataOut_payload_0_3091 : _zz_dataOut_payload_0_3079);
  assign _zz_dataOut_payload_0_3105 = (_zz_dataOut_payload_0_3082 < _zz_dataOut_payload_0_3094);
  assign _zz_dataOut_payload_0_3106 = (_zz_dataOut_payload_0_3105 ? _zz_dataOut_payload_0_3082 : _zz_dataOut_payload_0_3094);
  assign _zz_dataOut_payload_0_3107 = (_zz_dataOut_payload_0_3105 ? _zz_dataOut_payload_0_3094 : _zz_dataOut_payload_0_3082);
  assign _zz_dataOut_payload_0_3108 = (_zz_dataOut_payload_0_3097 < _zz_dataOut_payload_0_3103);
  assign _zz_dataOut_payload_0_3109 = (_zz_dataOut_payload_0_3108 ? _zz_dataOut_payload_0_3097 : _zz_dataOut_payload_0_3103);
  assign _zz_dataOut_payload_0_3110 = (_zz_dataOut_payload_0_3108 ? _zz_dataOut_payload_0_3103 : _zz_dataOut_payload_0_3097);
  assign _zz_dataOut_payload_0_3111 = (_zz_dataOut_payload_0_3100 < _zz_dataOut_payload_0_3106);
  assign _zz_dataOut_payload_0_3112 = (_zz_dataOut_payload_0_3111 ? _zz_dataOut_payload_0_3100 : _zz_dataOut_payload_0_3106);
  assign _zz_dataOut_payload_0_3113 = (_zz_dataOut_payload_0_3111 ? _zz_dataOut_payload_0_3106 : _zz_dataOut_payload_0_3100);
  assign _zz_dataOut_payload_0_3114 = (_zz_dataOut_payload_0_3109 < _zz_dataOut_payload_0_3112);
  assign _zz_dataOut_payload_0_3115 = (_zz_dataOut_payload_0_3110 < _zz_dataOut_payload_0_3113);
  assign _zz_dataOut_payload_0_3120 = (_zz_dataOut_payload_0_3098 < _zz_dataOut_payload_0_3104);
  assign _zz_dataOut_payload_0_3121 = (_zz_dataOut_payload_0_3120 ? _zz_dataOut_payload_0_3098 : _zz_dataOut_payload_0_3104);
  assign _zz_dataOut_payload_0_3122 = (_zz_dataOut_payload_0_3120 ? _zz_dataOut_payload_0_3104 : _zz_dataOut_payload_0_3098);
  assign _zz_dataOut_payload_0_3123 = (_zz_dataOut_payload_0_3101 < _zz_dataOut_payload_0_3107);
  assign _zz_dataOut_payload_0_3124 = (_zz_dataOut_payload_0_3123 ? _zz_dataOut_payload_0_3101 : _zz_dataOut_payload_0_3107);
  assign _zz_dataOut_payload_0_3125 = (_zz_dataOut_payload_0_3123 ? _zz_dataOut_payload_0_3107 : _zz_dataOut_payload_0_3101);
  assign _zz_dataOut_payload_0_3126 = (_zz_dataOut_payload_0_3121 < _zz_dataOut_payload_0_3124);
  assign _zz_dataOut_payload_0_3127 = (_zz_dataOut_payload_0_3122 < _zz_dataOut_payload_0_3125);
  assign _zz_dataOut_payload_0_3140 = (_zz_dataOut_payload_0_3095 < _zz_dataOut_payload_0_3083);
  assign _zz_dataOut_payload_0_3141 = (_zz_dataOut_payload_0_3140 ? _zz_dataOut_payload_0_3095 : _zz_dataOut_payload_0_3083);
  assign _zz_dataOut_payload_0_3142 = (_zz_dataOut_payload_0_3140 ? _zz_dataOut_payload_0_3083 : _zz_dataOut_payload_0_3095);
  assign _zz_dataOut_payload_0_3143 = (_zz_dataOut_payload_0_3092 < _zz_dataOut_payload_0_3080);
  assign _zz_dataOut_payload_0_3144 = (_zz_dataOut_payload_0_3143 ? _zz_dataOut_payload_0_3092 : _zz_dataOut_payload_0_3080);
  assign _zz_dataOut_payload_0_3145 = (_zz_dataOut_payload_0_3143 ? _zz_dataOut_payload_0_3080 : _zz_dataOut_payload_0_3092);
  assign _zz_dataOut_payload_0_3146 = (_zz_dataOut_payload_0_3089 < _zz_dataOut_payload_0_3077);
  assign _zz_dataOut_payload_0_3147 = (_zz_dataOut_payload_0_3146 ? _zz_dataOut_payload_0_3089 : _zz_dataOut_payload_0_3077);
  assign _zz_dataOut_payload_0_3148 = (_zz_dataOut_payload_0_3146 ? _zz_dataOut_payload_0_3077 : _zz_dataOut_payload_0_3089);
  assign _zz_dataOut_payload_0_3149 = (_zz_dataOut_payload_0_3086 < _zz_dataOut_payload_0_3074);
  assign _zz_dataOut_payload_0_3150 = (_zz_dataOut_payload_0_3149 ? _zz_dataOut_payload_0_3086 : _zz_dataOut_payload_0_3074);
  assign _zz_dataOut_payload_0_3151 = (_zz_dataOut_payload_0_3149 ? _zz_dataOut_payload_0_3074 : _zz_dataOut_payload_0_3086);
  assign _zz_dataOut_payload_0_3152 = (_zz_dataOut_payload_0_3141 < _zz_dataOut_payload_0_3147);
  assign _zz_dataOut_payload_0_3153 = (_zz_dataOut_payload_0_3152 ? _zz_dataOut_payload_0_3141 : _zz_dataOut_payload_0_3147);
  assign _zz_dataOut_payload_0_3154 = (_zz_dataOut_payload_0_3152 ? _zz_dataOut_payload_0_3147 : _zz_dataOut_payload_0_3141);
  assign _zz_dataOut_payload_0_3155 = (_zz_dataOut_payload_0_3144 < _zz_dataOut_payload_0_3150);
  assign _zz_dataOut_payload_0_3156 = (_zz_dataOut_payload_0_3155 ? _zz_dataOut_payload_0_3144 : _zz_dataOut_payload_0_3150);
  assign _zz_dataOut_payload_0_3157 = (_zz_dataOut_payload_0_3155 ? _zz_dataOut_payload_0_3150 : _zz_dataOut_payload_0_3144);
  assign _zz_dataOut_payload_0_3158 = (_zz_dataOut_payload_0_3153 < _zz_dataOut_payload_0_3156);
  assign _zz_dataOut_payload_0_3159 = (_zz_dataOut_payload_0_3154 < _zz_dataOut_payload_0_3157);
  assign _zz_dataOut_payload_0_3164 = (_zz_dataOut_payload_0_3142 < _zz_dataOut_payload_0_3148);
  assign _zz_dataOut_payload_0_3165 = (_zz_dataOut_payload_0_3164 ? _zz_dataOut_payload_0_3142 : _zz_dataOut_payload_0_3148);
  assign _zz_dataOut_payload_0_3166 = (_zz_dataOut_payload_0_3164 ? _zz_dataOut_payload_0_3148 : _zz_dataOut_payload_0_3142);
  assign _zz_dataOut_payload_0_3167 = (_zz_dataOut_payload_0_3145 < _zz_dataOut_payload_0_3151);
  assign _zz_dataOut_payload_0_3168 = (_zz_dataOut_payload_0_3167 ? _zz_dataOut_payload_0_3145 : _zz_dataOut_payload_0_3151);
  assign _zz_dataOut_payload_0_3169 = (_zz_dataOut_payload_0_3167 ? _zz_dataOut_payload_0_3151 : _zz_dataOut_payload_0_3145);
  assign _zz_dataOut_payload_0_3170 = (_zz_dataOut_payload_0_3165 < _zz_dataOut_payload_0_3168);
  assign _zz_dataOut_payload_0_3171 = (_zz_dataOut_payload_0_3166 < _zz_dataOut_payload_0_3169);
  assign _zz_dataOut_payload_0_3200 = (_zz_dataOut_payload_0_2832 < _zz_dataOut_payload_0_2847);
  assign _zz_dataOut_payload_0_3201 = (_zz_dataOut_payload_0_3200 ? _zz_dataOut_payload_0_2832 : _zz_dataOut_payload_0_2847);
  assign _zz_dataOut_payload_0_3202 = (_zz_dataOut_payload_0_3200 ? _zz_dataOut_payload_0_2847 : _zz_dataOut_payload_0_2832);
  assign _zz_dataOut_payload_0_3203 = (_zz_dataOut_payload_0_2833 < _zz_dataOut_payload_0_2846);
  assign _zz_dataOut_payload_0_3204 = (_zz_dataOut_payload_0_3203 ? _zz_dataOut_payload_0_2833 : _zz_dataOut_payload_0_2846);
  assign _zz_dataOut_payload_0_3205 = (_zz_dataOut_payload_0_3203 ? _zz_dataOut_payload_0_2846 : _zz_dataOut_payload_0_2833);
  assign _zz_dataOut_payload_0_3206 = (_zz_dataOut_payload_0_2834 < _zz_dataOut_payload_0_2845);
  assign _zz_dataOut_payload_0_3207 = (_zz_dataOut_payload_0_3206 ? _zz_dataOut_payload_0_2834 : _zz_dataOut_payload_0_2845);
  assign _zz_dataOut_payload_0_3208 = (_zz_dataOut_payload_0_3206 ? _zz_dataOut_payload_0_2845 : _zz_dataOut_payload_0_2834);
  assign _zz_dataOut_payload_0_3209 = (_zz_dataOut_payload_0_2835 < _zz_dataOut_payload_0_2844);
  assign _zz_dataOut_payload_0_3210 = (_zz_dataOut_payload_0_3209 ? _zz_dataOut_payload_0_2835 : _zz_dataOut_payload_0_2844);
  assign _zz_dataOut_payload_0_3211 = (_zz_dataOut_payload_0_3209 ? _zz_dataOut_payload_0_2844 : _zz_dataOut_payload_0_2835);
  assign _zz_dataOut_payload_0_3212 = (_zz_dataOut_payload_0_2836 < _zz_dataOut_payload_0_2843);
  assign _zz_dataOut_payload_0_3213 = (_zz_dataOut_payload_0_3212 ? _zz_dataOut_payload_0_2836 : _zz_dataOut_payload_0_2843);
  assign _zz_dataOut_payload_0_3214 = (_zz_dataOut_payload_0_3212 ? _zz_dataOut_payload_0_2843 : _zz_dataOut_payload_0_2836);
  assign _zz_dataOut_payload_0_3215 = (_zz_dataOut_payload_0_2837 < _zz_dataOut_payload_0_2842);
  assign _zz_dataOut_payload_0_3216 = (_zz_dataOut_payload_0_3215 ? _zz_dataOut_payload_0_2837 : _zz_dataOut_payload_0_2842);
  assign _zz_dataOut_payload_0_3217 = (_zz_dataOut_payload_0_3215 ? _zz_dataOut_payload_0_2842 : _zz_dataOut_payload_0_2837);
  assign _zz_dataOut_payload_0_3218 = (_zz_dataOut_payload_0_2838 < _zz_dataOut_payload_0_2841);
  assign _zz_dataOut_payload_0_3219 = (_zz_dataOut_payload_0_3218 ? _zz_dataOut_payload_0_2838 : _zz_dataOut_payload_0_2841);
  assign _zz_dataOut_payload_0_3220 = (_zz_dataOut_payload_0_3218 ? _zz_dataOut_payload_0_2841 : _zz_dataOut_payload_0_2838);
  assign _zz_dataOut_payload_0_3221 = (_zz_dataOut_payload_0_2839 < _zz_dataOut_payload_0_2840);
  assign _zz_dataOut_payload_0_3222 = (_zz_dataOut_payload_0_3221 ? _zz_dataOut_payload_0_2839 : _zz_dataOut_payload_0_2840);
  assign _zz_dataOut_payload_0_3223 = (_zz_dataOut_payload_0_3221 ? _zz_dataOut_payload_0_2840 : _zz_dataOut_payload_0_2839);
  assign _zz_dataOut_payload_0_3224 = (_zz_dataOut_payload_0_3201 < _zz_dataOut_payload_0_3213);
  assign _zz_dataOut_payload_0_3225 = (_zz_dataOut_payload_0_3224 ? _zz_dataOut_payload_0_3201 : _zz_dataOut_payload_0_3213);
  assign _zz_dataOut_payload_0_3226 = (_zz_dataOut_payload_0_3224 ? _zz_dataOut_payload_0_3213 : _zz_dataOut_payload_0_3201);
  assign _zz_dataOut_payload_0_3227 = (_zz_dataOut_payload_0_3204 < _zz_dataOut_payload_0_3216);
  assign _zz_dataOut_payload_0_3228 = (_zz_dataOut_payload_0_3227 ? _zz_dataOut_payload_0_3204 : _zz_dataOut_payload_0_3216);
  assign _zz_dataOut_payload_0_3229 = (_zz_dataOut_payload_0_3227 ? _zz_dataOut_payload_0_3216 : _zz_dataOut_payload_0_3204);
  assign _zz_dataOut_payload_0_3230 = (_zz_dataOut_payload_0_3207 < _zz_dataOut_payload_0_3219);
  assign _zz_dataOut_payload_0_3231 = (_zz_dataOut_payload_0_3230 ? _zz_dataOut_payload_0_3207 : _zz_dataOut_payload_0_3219);
  assign _zz_dataOut_payload_0_3232 = (_zz_dataOut_payload_0_3230 ? _zz_dataOut_payload_0_3219 : _zz_dataOut_payload_0_3207);
  assign _zz_dataOut_payload_0_3233 = (_zz_dataOut_payload_0_3210 < _zz_dataOut_payload_0_3222);
  assign _zz_dataOut_payload_0_3234 = (_zz_dataOut_payload_0_3233 ? _zz_dataOut_payload_0_3210 : _zz_dataOut_payload_0_3222);
  assign _zz_dataOut_payload_0_3235 = (_zz_dataOut_payload_0_3233 ? _zz_dataOut_payload_0_3222 : _zz_dataOut_payload_0_3210);
  assign _zz_dataOut_payload_0_3236 = (_zz_dataOut_payload_0_3225 < _zz_dataOut_payload_0_3231);
  assign _zz_dataOut_payload_0_3237 = (_zz_dataOut_payload_0_3236 ? _zz_dataOut_payload_0_3225 : _zz_dataOut_payload_0_3231);
  assign _zz_dataOut_payload_0_3238 = (_zz_dataOut_payload_0_3236 ? _zz_dataOut_payload_0_3231 : _zz_dataOut_payload_0_3225);
  assign _zz_dataOut_payload_0_3239 = (_zz_dataOut_payload_0_3228 < _zz_dataOut_payload_0_3234);
  assign _zz_dataOut_payload_0_3240 = (_zz_dataOut_payload_0_3239 ? _zz_dataOut_payload_0_3228 : _zz_dataOut_payload_0_3234);
  assign _zz_dataOut_payload_0_3241 = (_zz_dataOut_payload_0_3239 ? _zz_dataOut_payload_0_3234 : _zz_dataOut_payload_0_3228);
  assign _zz_dataOut_payload_0_3242 = (_zz_dataOut_payload_0_3237 < _zz_dataOut_payload_0_3240);
  assign _zz_dataOut_payload_0_3243 = (_zz_dataOut_payload_0_3238 < _zz_dataOut_payload_0_3241);
  assign _zz_dataOut_payload_0_3248 = (_zz_dataOut_payload_0_3226 < _zz_dataOut_payload_0_3232);
  assign _zz_dataOut_payload_0_3249 = (_zz_dataOut_payload_0_3248 ? _zz_dataOut_payload_0_3226 : _zz_dataOut_payload_0_3232);
  assign _zz_dataOut_payload_0_3250 = (_zz_dataOut_payload_0_3248 ? _zz_dataOut_payload_0_3232 : _zz_dataOut_payload_0_3226);
  assign _zz_dataOut_payload_0_3251 = (_zz_dataOut_payload_0_3229 < _zz_dataOut_payload_0_3235);
  assign _zz_dataOut_payload_0_3252 = (_zz_dataOut_payload_0_3251 ? _zz_dataOut_payload_0_3229 : _zz_dataOut_payload_0_3235);
  assign _zz_dataOut_payload_0_3253 = (_zz_dataOut_payload_0_3251 ? _zz_dataOut_payload_0_3235 : _zz_dataOut_payload_0_3229);
  assign _zz_dataOut_payload_0_3254 = (_zz_dataOut_payload_0_3249 < _zz_dataOut_payload_0_3252);
  assign _zz_dataOut_payload_0_3255 = (_zz_dataOut_payload_0_3250 < _zz_dataOut_payload_0_3253);
  assign _zz_dataOut_payload_0_3268 = (_zz_dataOut_payload_0_3223 < _zz_dataOut_payload_0_3211);
  assign _zz_dataOut_payload_0_3269 = (_zz_dataOut_payload_0_3268 ? _zz_dataOut_payload_0_3223 : _zz_dataOut_payload_0_3211);
  assign _zz_dataOut_payload_0_3270 = (_zz_dataOut_payload_0_3268 ? _zz_dataOut_payload_0_3211 : _zz_dataOut_payload_0_3223);
  assign _zz_dataOut_payload_0_3271 = (_zz_dataOut_payload_0_3220 < _zz_dataOut_payload_0_3208);
  assign _zz_dataOut_payload_0_3272 = (_zz_dataOut_payload_0_3271 ? _zz_dataOut_payload_0_3220 : _zz_dataOut_payload_0_3208);
  assign _zz_dataOut_payload_0_3273 = (_zz_dataOut_payload_0_3271 ? _zz_dataOut_payload_0_3208 : _zz_dataOut_payload_0_3220);
  assign _zz_dataOut_payload_0_3274 = (_zz_dataOut_payload_0_3217 < _zz_dataOut_payload_0_3205);
  assign _zz_dataOut_payload_0_3275 = (_zz_dataOut_payload_0_3274 ? _zz_dataOut_payload_0_3217 : _zz_dataOut_payload_0_3205);
  assign _zz_dataOut_payload_0_3276 = (_zz_dataOut_payload_0_3274 ? _zz_dataOut_payload_0_3205 : _zz_dataOut_payload_0_3217);
  assign _zz_dataOut_payload_0_3277 = (_zz_dataOut_payload_0_3214 < _zz_dataOut_payload_0_3202);
  assign _zz_dataOut_payload_0_3278 = (_zz_dataOut_payload_0_3277 ? _zz_dataOut_payload_0_3214 : _zz_dataOut_payload_0_3202);
  assign _zz_dataOut_payload_0_3279 = (_zz_dataOut_payload_0_3277 ? _zz_dataOut_payload_0_3202 : _zz_dataOut_payload_0_3214);
  assign _zz_dataOut_payload_0_3280 = (_zz_dataOut_payload_0_3269 < _zz_dataOut_payload_0_3275);
  assign _zz_dataOut_payload_0_3281 = (_zz_dataOut_payload_0_3280 ? _zz_dataOut_payload_0_3269 : _zz_dataOut_payload_0_3275);
  assign _zz_dataOut_payload_0_3282 = (_zz_dataOut_payload_0_3280 ? _zz_dataOut_payload_0_3275 : _zz_dataOut_payload_0_3269);
  assign _zz_dataOut_payload_0_3283 = (_zz_dataOut_payload_0_3272 < _zz_dataOut_payload_0_3278);
  assign _zz_dataOut_payload_0_3284 = (_zz_dataOut_payload_0_3283 ? _zz_dataOut_payload_0_3272 : _zz_dataOut_payload_0_3278);
  assign _zz_dataOut_payload_0_3285 = (_zz_dataOut_payload_0_3283 ? _zz_dataOut_payload_0_3278 : _zz_dataOut_payload_0_3272);
  assign _zz_dataOut_payload_0_3286 = (_zz_dataOut_payload_0_3281 < _zz_dataOut_payload_0_3284);
  assign _zz_dataOut_payload_0_3287 = (_zz_dataOut_payload_0_3282 < _zz_dataOut_payload_0_3285);
  assign _zz_dataOut_payload_0_3292 = (_zz_dataOut_payload_0_3270 < _zz_dataOut_payload_0_3276);
  assign _zz_dataOut_payload_0_3293 = (_zz_dataOut_payload_0_3292 ? _zz_dataOut_payload_0_3270 : _zz_dataOut_payload_0_3276);
  assign _zz_dataOut_payload_0_3294 = (_zz_dataOut_payload_0_3292 ? _zz_dataOut_payload_0_3276 : _zz_dataOut_payload_0_3270);
  assign _zz_dataOut_payload_0_3295 = (_zz_dataOut_payload_0_3273 < _zz_dataOut_payload_0_3279);
  assign _zz_dataOut_payload_0_3296 = (_zz_dataOut_payload_0_3295 ? _zz_dataOut_payload_0_3273 : _zz_dataOut_payload_0_3279);
  assign _zz_dataOut_payload_0_3297 = (_zz_dataOut_payload_0_3295 ? _zz_dataOut_payload_0_3279 : _zz_dataOut_payload_0_3273);
  assign _zz_dataOut_payload_0_3298 = (_zz_dataOut_payload_0_3293 < _zz_dataOut_payload_0_3296);
  assign _zz_dataOut_payload_0_3299 = (_zz_dataOut_payload_0_3294 < _zz_dataOut_payload_0_3297);
  assign _zz_dataOut_payload_0_3328 = (_zz_dataOut_payload_0_2848 < _zz_dataOut_payload_0_2863);
  assign _zz_dataOut_payload_0_3329 = (_zz_dataOut_payload_0_3328 ? _zz_dataOut_payload_0_2848 : _zz_dataOut_payload_0_2863);
  assign _zz_dataOut_payload_0_3330 = (_zz_dataOut_payload_0_3328 ? _zz_dataOut_payload_0_2863 : _zz_dataOut_payload_0_2848);
  assign _zz_dataOut_payload_0_3331 = (_zz_dataOut_payload_0_2849 < _zz_dataOut_payload_0_2862);
  assign _zz_dataOut_payload_0_3332 = (_zz_dataOut_payload_0_3331 ? _zz_dataOut_payload_0_2849 : _zz_dataOut_payload_0_2862);
  assign _zz_dataOut_payload_0_3333 = (_zz_dataOut_payload_0_3331 ? _zz_dataOut_payload_0_2862 : _zz_dataOut_payload_0_2849);
  assign _zz_dataOut_payload_0_3334 = (_zz_dataOut_payload_0_2850 < _zz_dataOut_payload_0_2861);
  assign _zz_dataOut_payload_0_3335 = (_zz_dataOut_payload_0_3334 ? _zz_dataOut_payload_0_2850 : _zz_dataOut_payload_0_2861);
  assign _zz_dataOut_payload_0_3336 = (_zz_dataOut_payload_0_3334 ? _zz_dataOut_payload_0_2861 : _zz_dataOut_payload_0_2850);
  assign _zz_dataOut_payload_0_3337 = (_zz_dataOut_payload_0_2851 < _zz_dataOut_payload_0_2860);
  assign _zz_dataOut_payload_0_3338 = (_zz_dataOut_payload_0_3337 ? _zz_dataOut_payload_0_2851 : _zz_dataOut_payload_0_2860);
  assign _zz_dataOut_payload_0_3339 = (_zz_dataOut_payload_0_3337 ? _zz_dataOut_payload_0_2860 : _zz_dataOut_payload_0_2851);
  assign _zz_dataOut_payload_0_3340 = (_zz_dataOut_payload_0_2852 < _zz_dataOut_payload_0_2859);
  assign _zz_dataOut_payload_0_3341 = (_zz_dataOut_payload_0_3340 ? _zz_dataOut_payload_0_2852 : _zz_dataOut_payload_0_2859);
  assign _zz_dataOut_payload_0_3342 = (_zz_dataOut_payload_0_3340 ? _zz_dataOut_payload_0_2859 : _zz_dataOut_payload_0_2852);
  assign _zz_dataOut_payload_0_3343 = (_zz_dataOut_payload_0_2853 < _zz_dataOut_payload_0_2858);
  assign _zz_dataOut_payload_0_3344 = (_zz_dataOut_payload_0_3343 ? _zz_dataOut_payload_0_2853 : _zz_dataOut_payload_0_2858);
  assign _zz_dataOut_payload_0_3345 = (_zz_dataOut_payload_0_3343 ? _zz_dataOut_payload_0_2858 : _zz_dataOut_payload_0_2853);
  assign _zz_dataOut_payload_0_3346 = (_zz_dataOut_payload_0_2854 < _zz_dataOut_payload_0_2857);
  assign _zz_dataOut_payload_0_3347 = (_zz_dataOut_payload_0_3346 ? _zz_dataOut_payload_0_2854 : _zz_dataOut_payload_0_2857);
  assign _zz_dataOut_payload_0_3348 = (_zz_dataOut_payload_0_3346 ? _zz_dataOut_payload_0_2857 : _zz_dataOut_payload_0_2854);
  assign _zz_dataOut_payload_0_3349 = (_zz_dataOut_payload_0_2855 < _zz_dataOut_payload_0_2856);
  assign _zz_dataOut_payload_0_3350 = (_zz_dataOut_payload_0_3349 ? _zz_dataOut_payload_0_2855 : _zz_dataOut_payload_0_2856);
  assign _zz_dataOut_payload_0_3351 = (_zz_dataOut_payload_0_3349 ? _zz_dataOut_payload_0_2856 : _zz_dataOut_payload_0_2855);
  assign _zz_dataOut_payload_0_3352 = (_zz_dataOut_payload_0_3329 < _zz_dataOut_payload_0_3341);
  assign _zz_dataOut_payload_0_3353 = (_zz_dataOut_payload_0_3352 ? _zz_dataOut_payload_0_3329 : _zz_dataOut_payload_0_3341);
  assign _zz_dataOut_payload_0_3354 = (_zz_dataOut_payload_0_3352 ? _zz_dataOut_payload_0_3341 : _zz_dataOut_payload_0_3329);
  assign _zz_dataOut_payload_0_3355 = (_zz_dataOut_payload_0_3332 < _zz_dataOut_payload_0_3344);
  assign _zz_dataOut_payload_0_3356 = (_zz_dataOut_payload_0_3355 ? _zz_dataOut_payload_0_3332 : _zz_dataOut_payload_0_3344);
  assign _zz_dataOut_payload_0_3357 = (_zz_dataOut_payload_0_3355 ? _zz_dataOut_payload_0_3344 : _zz_dataOut_payload_0_3332);
  assign _zz_dataOut_payload_0_3358 = (_zz_dataOut_payload_0_3335 < _zz_dataOut_payload_0_3347);
  assign _zz_dataOut_payload_0_3359 = (_zz_dataOut_payload_0_3358 ? _zz_dataOut_payload_0_3335 : _zz_dataOut_payload_0_3347);
  assign _zz_dataOut_payload_0_3360 = (_zz_dataOut_payload_0_3358 ? _zz_dataOut_payload_0_3347 : _zz_dataOut_payload_0_3335);
  assign _zz_dataOut_payload_0_3361 = (_zz_dataOut_payload_0_3338 < _zz_dataOut_payload_0_3350);
  assign _zz_dataOut_payload_0_3362 = (_zz_dataOut_payload_0_3361 ? _zz_dataOut_payload_0_3338 : _zz_dataOut_payload_0_3350);
  assign _zz_dataOut_payload_0_3363 = (_zz_dataOut_payload_0_3361 ? _zz_dataOut_payload_0_3350 : _zz_dataOut_payload_0_3338);
  assign _zz_dataOut_payload_0_3364 = (_zz_dataOut_payload_0_3353 < _zz_dataOut_payload_0_3359);
  assign _zz_dataOut_payload_0_3365 = (_zz_dataOut_payload_0_3364 ? _zz_dataOut_payload_0_3353 : _zz_dataOut_payload_0_3359);
  assign _zz_dataOut_payload_0_3366 = (_zz_dataOut_payload_0_3364 ? _zz_dataOut_payload_0_3359 : _zz_dataOut_payload_0_3353);
  assign _zz_dataOut_payload_0_3367 = (_zz_dataOut_payload_0_3356 < _zz_dataOut_payload_0_3362);
  assign _zz_dataOut_payload_0_3368 = (_zz_dataOut_payload_0_3367 ? _zz_dataOut_payload_0_3356 : _zz_dataOut_payload_0_3362);
  assign _zz_dataOut_payload_0_3369 = (_zz_dataOut_payload_0_3367 ? _zz_dataOut_payload_0_3362 : _zz_dataOut_payload_0_3356);
  assign _zz_dataOut_payload_0_3370 = (_zz_dataOut_payload_0_3365 < _zz_dataOut_payload_0_3368);
  assign _zz_dataOut_payload_0_3371 = (_zz_dataOut_payload_0_3366 < _zz_dataOut_payload_0_3369);
  assign _zz_dataOut_payload_0_3376 = (_zz_dataOut_payload_0_3354 < _zz_dataOut_payload_0_3360);
  assign _zz_dataOut_payload_0_3377 = (_zz_dataOut_payload_0_3376 ? _zz_dataOut_payload_0_3354 : _zz_dataOut_payload_0_3360);
  assign _zz_dataOut_payload_0_3378 = (_zz_dataOut_payload_0_3376 ? _zz_dataOut_payload_0_3360 : _zz_dataOut_payload_0_3354);
  assign _zz_dataOut_payload_0_3379 = (_zz_dataOut_payload_0_3357 < _zz_dataOut_payload_0_3363);
  assign _zz_dataOut_payload_0_3380 = (_zz_dataOut_payload_0_3379 ? _zz_dataOut_payload_0_3357 : _zz_dataOut_payload_0_3363);
  assign _zz_dataOut_payload_0_3381 = (_zz_dataOut_payload_0_3379 ? _zz_dataOut_payload_0_3363 : _zz_dataOut_payload_0_3357);
  assign _zz_dataOut_payload_0_3382 = (_zz_dataOut_payload_0_3377 < _zz_dataOut_payload_0_3380);
  assign _zz_dataOut_payload_0_3383 = (_zz_dataOut_payload_0_3378 < _zz_dataOut_payload_0_3381);
  assign _zz_dataOut_payload_0_3396 = (_zz_dataOut_payload_0_3351 < _zz_dataOut_payload_0_3339);
  assign _zz_dataOut_payload_0_3397 = (_zz_dataOut_payload_0_3396 ? _zz_dataOut_payload_0_3351 : _zz_dataOut_payload_0_3339);
  assign _zz_dataOut_payload_0_3398 = (_zz_dataOut_payload_0_3396 ? _zz_dataOut_payload_0_3339 : _zz_dataOut_payload_0_3351);
  assign _zz_dataOut_payload_0_3399 = (_zz_dataOut_payload_0_3348 < _zz_dataOut_payload_0_3336);
  assign _zz_dataOut_payload_0_3400 = (_zz_dataOut_payload_0_3399 ? _zz_dataOut_payload_0_3348 : _zz_dataOut_payload_0_3336);
  assign _zz_dataOut_payload_0_3401 = (_zz_dataOut_payload_0_3399 ? _zz_dataOut_payload_0_3336 : _zz_dataOut_payload_0_3348);
  assign _zz_dataOut_payload_0_3402 = (_zz_dataOut_payload_0_3345 < _zz_dataOut_payload_0_3333);
  assign _zz_dataOut_payload_0_3403 = (_zz_dataOut_payload_0_3402 ? _zz_dataOut_payload_0_3345 : _zz_dataOut_payload_0_3333);
  assign _zz_dataOut_payload_0_3404 = (_zz_dataOut_payload_0_3402 ? _zz_dataOut_payload_0_3333 : _zz_dataOut_payload_0_3345);
  assign _zz_dataOut_payload_0_3405 = (_zz_dataOut_payload_0_3342 < _zz_dataOut_payload_0_3330);
  assign _zz_dataOut_payload_0_3406 = (_zz_dataOut_payload_0_3405 ? _zz_dataOut_payload_0_3342 : _zz_dataOut_payload_0_3330);
  assign _zz_dataOut_payload_0_3407 = (_zz_dataOut_payload_0_3405 ? _zz_dataOut_payload_0_3330 : _zz_dataOut_payload_0_3342);
  assign _zz_dataOut_payload_0_3408 = (_zz_dataOut_payload_0_3397 < _zz_dataOut_payload_0_3403);
  assign _zz_dataOut_payload_0_3409 = (_zz_dataOut_payload_0_3408 ? _zz_dataOut_payload_0_3397 : _zz_dataOut_payload_0_3403);
  assign _zz_dataOut_payload_0_3410 = (_zz_dataOut_payload_0_3408 ? _zz_dataOut_payload_0_3403 : _zz_dataOut_payload_0_3397);
  assign _zz_dataOut_payload_0_3411 = (_zz_dataOut_payload_0_3400 < _zz_dataOut_payload_0_3406);
  assign _zz_dataOut_payload_0_3412 = (_zz_dataOut_payload_0_3411 ? _zz_dataOut_payload_0_3400 : _zz_dataOut_payload_0_3406);
  assign _zz_dataOut_payload_0_3413 = (_zz_dataOut_payload_0_3411 ? _zz_dataOut_payload_0_3406 : _zz_dataOut_payload_0_3400);
  assign _zz_dataOut_payload_0_3414 = (_zz_dataOut_payload_0_3409 < _zz_dataOut_payload_0_3412);
  assign _zz_dataOut_payload_0_3415 = (_zz_dataOut_payload_0_3410 < _zz_dataOut_payload_0_3413);
  assign _zz_dataOut_payload_0_3420 = (_zz_dataOut_payload_0_3398 < _zz_dataOut_payload_0_3404);
  assign _zz_dataOut_payload_0_3421 = (_zz_dataOut_payload_0_3420 ? _zz_dataOut_payload_0_3398 : _zz_dataOut_payload_0_3404);
  assign _zz_dataOut_payload_0_3422 = (_zz_dataOut_payload_0_3420 ? _zz_dataOut_payload_0_3404 : _zz_dataOut_payload_0_3398);
  assign _zz_dataOut_payload_0_3423 = (_zz_dataOut_payload_0_3401 < _zz_dataOut_payload_0_3407);
  assign _zz_dataOut_payload_0_3424 = (_zz_dataOut_payload_0_3423 ? _zz_dataOut_payload_0_3401 : _zz_dataOut_payload_0_3407);
  assign _zz_dataOut_payload_0_3425 = (_zz_dataOut_payload_0_3423 ? _zz_dataOut_payload_0_3407 : _zz_dataOut_payload_0_3401);
  assign _zz_dataOut_payload_0_3426 = (_zz_dataOut_payload_0_3421 < _zz_dataOut_payload_0_3424);
  assign _zz_dataOut_payload_0_3427 = (_zz_dataOut_payload_0_3422 < _zz_dataOut_payload_0_3425);
  assign _zz_dataOut_payload_0_3456 = (_zz_dataOut_payload_0_2864 < _zz_dataOut_payload_0_2879);
  assign _zz_dataOut_payload_0_3457 = (_zz_dataOut_payload_0_3456 ? _zz_dataOut_payload_0_2864 : _zz_dataOut_payload_0_2879);
  assign _zz_dataOut_payload_0_3458 = (_zz_dataOut_payload_0_3456 ? _zz_dataOut_payload_0_2879 : _zz_dataOut_payload_0_2864);
  assign _zz_dataOut_payload_0_3459 = (_zz_dataOut_payload_0_2865 < _zz_dataOut_payload_0_2878);
  assign _zz_dataOut_payload_0_3460 = (_zz_dataOut_payload_0_3459 ? _zz_dataOut_payload_0_2865 : _zz_dataOut_payload_0_2878);
  assign _zz_dataOut_payload_0_3461 = (_zz_dataOut_payload_0_3459 ? _zz_dataOut_payload_0_2878 : _zz_dataOut_payload_0_2865);
  assign _zz_dataOut_payload_0_3462 = (_zz_dataOut_payload_0_2866 < _zz_dataOut_payload_0_2877);
  assign _zz_dataOut_payload_0_3463 = (_zz_dataOut_payload_0_3462 ? _zz_dataOut_payload_0_2866 : _zz_dataOut_payload_0_2877);
  assign _zz_dataOut_payload_0_3464 = (_zz_dataOut_payload_0_3462 ? _zz_dataOut_payload_0_2877 : _zz_dataOut_payload_0_2866);
  assign _zz_dataOut_payload_0_3465 = (_zz_dataOut_payload_0_2867 < _zz_dataOut_payload_0_2876);
  assign _zz_dataOut_payload_0_3466 = (_zz_dataOut_payload_0_3465 ? _zz_dataOut_payload_0_2867 : _zz_dataOut_payload_0_2876);
  assign _zz_dataOut_payload_0_3467 = (_zz_dataOut_payload_0_3465 ? _zz_dataOut_payload_0_2876 : _zz_dataOut_payload_0_2867);
  assign _zz_dataOut_payload_0_3468 = (_zz_dataOut_payload_0_2868 < _zz_dataOut_payload_0_2875);
  assign _zz_dataOut_payload_0_3469 = (_zz_dataOut_payload_0_3468 ? _zz_dataOut_payload_0_2868 : _zz_dataOut_payload_0_2875);
  assign _zz_dataOut_payload_0_3470 = (_zz_dataOut_payload_0_3468 ? _zz_dataOut_payload_0_2875 : _zz_dataOut_payload_0_2868);
  assign _zz_dataOut_payload_0_3471 = (_zz_dataOut_payload_0_2869 < _zz_dataOut_payload_0_2874);
  assign _zz_dataOut_payload_0_3472 = (_zz_dataOut_payload_0_3471 ? _zz_dataOut_payload_0_2869 : _zz_dataOut_payload_0_2874);
  assign _zz_dataOut_payload_0_3473 = (_zz_dataOut_payload_0_3471 ? _zz_dataOut_payload_0_2874 : _zz_dataOut_payload_0_2869);
  assign _zz_dataOut_payload_0_3474 = (_zz_dataOut_payload_0_2870 < _zz_dataOut_payload_0_2873);
  assign _zz_dataOut_payload_0_3475 = (_zz_dataOut_payload_0_3474 ? _zz_dataOut_payload_0_2870 : _zz_dataOut_payload_0_2873);
  assign _zz_dataOut_payload_0_3476 = (_zz_dataOut_payload_0_3474 ? _zz_dataOut_payload_0_2873 : _zz_dataOut_payload_0_2870);
  assign _zz_dataOut_payload_0_3477 = (_zz_dataOut_payload_0_2871 < _zz_dataOut_payload_0_2872);
  assign _zz_dataOut_payload_0_3478 = (_zz_dataOut_payload_0_3477 ? _zz_dataOut_payload_0_2871 : _zz_dataOut_payload_0_2872);
  assign _zz_dataOut_payload_0_3479 = (_zz_dataOut_payload_0_3477 ? _zz_dataOut_payload_0_2872 : _zz_dataOut_payload_0_2871);
  assign _zz_dataOut_payload_0_3480 = (_zz_dataOut_payload_0_3457 < _zz_dataOut_payload_0_3469);
  assign _zz_dataOut_payload_0_3481 = (_zz_dataOut_payload_0_3480 ? _zz_dataOut_payload_0_3457 : _zz_dataOut_payload_0_3469);
  assign _zz_dataOut_payload_0_3482 = (_zz_dataOut_payload_0_3480 ? _zz_dataOut_payload_0_3469 : _zz_dataOut_payload_0_3457);
  assign _zz_dataOut_payload_0_3483 = (_zz_dataOut_payload_0_3460 < _zz_dataOut_payload_0_3472);
  assign _zz_dataOut_payload_0_3484 = (_zz_dataOut_payload_0_3483 ? _zz_dataOut_payload_0_3460 : _zz_dataOut_payload_0_3472);
  assign _zz_dataOut_payload_0_3485 = (_zz_dataOut_payload_0_3483 ? _zz_dataOut_payload_0_3472 : _zz_dataOut_payload_0_3460);
  assign _zz_dataOut_payload_0_3486 = (_zz_dataOut_payload_0_3463 < _zz_dataOut_payload_0_3475);
  assign _zz_dataOut_payload_0_3487 = (_zz_dataOut_payload_0_3486 ? _zz_dataOut_payload_0_3463 : _zz_dataOut_payload_0_3475);
  assign _zz_dataOut_payload_0_3488 = (_zz_dataOut_payload_0_3486 ? _zz_dataOut_payload_0_3475 : _zz_dataOut_payload_0_3463);
  assign _zz_dataOut_payload_0_3489 = (_zz_dataOut_payload_0_3466 < _zz_dataOut_payload_0_3478);
  assign _zz_dataOut_payload_0_3490 = (_zz_dataOut_payload_0_3489 ? _zz_dataOut_payload_0_3466 : _zz_dataOut_payload_0_3478);
  assign _zz_dataOut_payload_0_3491 = (_zz_dataOut_payload_0_3489 ? _zz_dataOut_payload_0_3478 : _zz_dataOut_payload_0_3466);
  assign _zz_dataOut_payload_0_3492 = (_zz_dataOut_payload_0_3481 < _zz_dataOut_payload_0_3487);
  assign _zz_dataOut_payload_0_3493 = (_zz_dataOut_payload_0_3492 ? _zz_dataOut_payload_0_3481 : _zz_dataOut_payload_0_3487);
  assign _zz_dataOut_payload_0_3494 = (_zz_dataOut_payload_0_3492 ? _zz_dataOut_payload_0_3487 : _zz_dataOut_payload_0_3481);
  assign _zz_dataOut_payload_0_3495 = (_zz_dataOut_payload_0_3484 < _zz_dataOut_payload_0_3490);
  assign _zz_dataOut_payload_0_3496 = (_zz_dataOut_payload_0_3495 ? _zz_dataOut_payload_0_3484 : _zz_dataOut_payload_0_3490);
  assign _zz_dataOut_payload_0_3497 = (_zz_dataOut_payload_0_3495 ? _zz_dataOut_payload_0_3490 : _zz_dataOut_payload_0_3484);
  assign _zz_dataOut_payload_0_3498 = (_zz_dataOut_payload_0_3493 < _zz_dataOut_payload_0_3496);
  assign _zz_dataOut_payload_0_3499 = (_zz_dataOut_payload_0_3494 < _zz_dataOut_payload_0_3497);
  assign _zz_dataOut_payload_0_3504 = (_zz_dataOut_payload_0_3482 < _zz_dataOut_payload_0_3488);
  assign _zz_dataOut_payload_0_3505 = (_zz_dataOut_payload_0_3504 ? _zz_dataOut_payload_0_3482 : _zz_dataOut_payload_0_3488);
  assign _zz_dataOut_payload_0_3506 = (_zz_dataOut_payload_0_3504 ? _zz_dataOut_payload_0_3488 : _zz_dataOut_payload_0_3482);
  assign _zz_dataOut_payload_0_3507 = (_zz_dataOut_payload_0_3485 < _zz_dataOut_payload_0_3491);
  assign _zz_dataOut_payload_0_3508 = (_zz_dataOut_payload_0_3507 ? _zz_dataOut_payload_0_3485 : _zz_dataOut_payload_0_3491);
  assign _zz_dataOut_payload_0_3509 = (_zz_dataOut_payload_0_3507 ? _zz_dataOut_payload_0_3491 : _zz_dataOut_payload_0_3485);
  assign _zz_dataOut_payload_0_3510 = (_zz_dataOut_payload_0_3505 < _zz_dataOut_payload_0_3508);
  assign _zz_dataOut_payload_0_3511 = (_zz_dataOut_payload_0_3506 < _zz_dataOut_payload_0_3509);
  assign _zz_dataOut_payload_0_3524 = (_zz_dataOut_payload_0_3479 < _zz_dataOut_payload_0_3467);
  assign _zz_dataOut_payload_0_3525 = (_zz_dataOut_payload_0_3524 ? _zz_dataOut_payload_0_3479 : _zz_dataOut_payload_0_3467);
  assign _zz_dataOut_payload_0_3526 = (_zz_dataOut_payload_0_3524 ? _zz_dataOut_payload_0_3467 : _zz_dataOut_payload_0_3479);
  assign _zz_dataOut_payload_0_3527 = (_zz_dataOut_payload_0_3476 < _zz_dataOut_payload_0_3464);
  assign _zz_dataOut_payload_0_3528 = (_zz_dataOut_payload_0_3527 ? _zz_dataOut_payload_0_3476 : _zz_dataOut_payload_0_3464);
  assign _zz_dataOut_payload_0_3529 = (_zz_dataOut_payload_0_3527 ? _zz_dataOut_payload_0_3464 : _zz_dataOut_payload_0_3476);
  assign _zz_dataOut_payload_0_3530 = (_zz_dataOut_payload_0_3473 < _zz_dataOut_payload_0_3461);
  assign _zz_dataOut_payload_0_3531 = (_zz_dataOut_payload_0_3530 ? _zz_dataOut_payload_0_3473 : _zz_dataOut_payload_0_3461);
  assign _zz_dataOut_payload_0_3532 = (_zz_dataOut_payload_0_3530 ? _zz_dataOut_payload_0_3461 : _zz_dataOut_payload_0_3473);
  assign _zz_dataOut_payload_0_3533 = (_zz_dataOut_payload_0_3470 < _zz_dataOut_payload_0_3458);
  assign _zz_dataOut_payload_0_3534 = (_zz_dataOut_payload_0_3533 ? _zz_dataOut_payload_0_3470 : _zz_dataOut_payload_0_3458);
  assign _zz_dataOut_payload_0_3535 = (_zz_dataOut_payload_0_3533 ? _zz_dataOut_payload_0_3458 : _zz_dataOut_payload_0_3470);
  assign _zz_dataOut_payload_0_3536 = (_zz_dataOut_payload_0_3525 < _zz_dataOut_payload_0_3531);
  assign _zz_dataOut_payload_0_3537 = (_zz_dataOut_payload_0_3536 ? _zz_dataOut_payload_0_3525 : _zz_dataOut_payload_0_3531);
  assign _zz_dataOut_payload_0_3538 = (_zz_dataOut_payload_0_3536 ? _zz_dataOut_payload_0_3531 : _zz_dataOut_payload_0_3525);
  assign _zz_dataOut_payload_0_3539 = (_zz_dataOut_payload_0_3528 < _zz_dataOut_payload_0_3534);
  assign _zz_dataOut_payload_0_3540 = (_zz_dataOut_payload_0_3539 ? _zz_dataOut_payload_0_3528 : _zz_dataOut_payload_0_3534);
  assign _zz_dataOut_payload_0_3541 = (_zz_dataOut_payload_0_3539 ? _zz_dataOut_payload_0_3534 : _zz_dataOut_payload_0_3528);
  assign _zz_dataOut_payload_0_3542 = (_zz_dataOut_payload_0_3537 < _zz_dataOut_payload_0_3540);
  assign _zz_dataOut_payload_0_3543 = (_zz_dataOut_payload_0_3538 < _zz_dataOut_payload_0_3541);
  assign _zz_dataOut_payload_0_3548 = (_zz_dataOut_payload_0_3526 < _zz_dataOut_payload_0_3532);
  assign _zz_dataOut_payload_0_3549 = (_zz_dataOut_payload_0_3548 ? _zz_dataOut_payload_0_3526 : _zz_dataOut_payload_0_3532);
  assign _zz_dataOut_payload_0_3550 = (_zz_dataOut_payload_0_3548 ? _zz_dataOut_payload_0_3532 : _zz_dataOut_payload_0_3526);
  assign _zz_dataOut_payload_0_3551 = (_zz_dataOut_payload_0_3529 < _zz_dataOut_payload_0_3535);
  assign _zz_dataOut_payload_0_3552 = (_zz_dataOut_payload_0_3551 ? _zz_dataOut_payload_0_3529 : _zz_dataOut_payload_0_3535);
  assign _zz_dataOut_payload_0_3553 = (_zz_dataOut_payload_0_3551 ? _zz_dataOut_payload_0_3535 : _zz_dataOut_payload_0_3529);
  assign _zz_dataOut_payload_0_3554 = (_zz_dataOut_payload_0_3549 < _zz_dataOut_payload_0_3552);
  assign _zz_dataOut_payload_0_3555 = (_zz_dataOut_payload_0_3550 < _zz_dataOut_payload_0_3553);
  assign _zz_dataOut_payload_0_3584 = (_zz_dataOut_payload_0_2880 < _zz_dataOut_payload_0_2895);
  assign _zz_dataOut_payload_0_3585 = (_zz_dataOut_payload_0_3584 ? _zz_dataOut_payload_0_2880 : _zz_dataOut_payload_0_2895);
  assign _zz_dataOut_payload_0_3586 = (_zz_dataOut_payload_0_3584 ? _zz_dataOut_payload_0_2895 : _zz_dataOut_payload_0_2880);
  assign _zz_dataOut_payload_0_3587 = (_zz_dataOut_payload_0_2881 < _zz_dataOut_payload_0_2894);
  assign _zz_dataOut_payload_0_3588 = (_zz_dataOut_payload_0_3587 ? _zz_dataOut_payload_0_2881 : _zz_dataOut_payload_0_2894);
  assign _zz_dataOut_payload_0_3589 = (_zz_dataOut_payload_0_3587 ? _zz_dataOut_payload_0_2894 : _zz_dataOut_payload_0_2881);
  assign _zz_dataOut_payload_0_3590 = (_zz_dataOut_payload_0_2882 < _zz_dataOut_payload_0_2893);
  assign _zz_dataOut_payload_0_3591 = (_zz_dataOut_payload_0_3590 ? _zz_dataOut_payload_0_2882 : _zz_dataOut_payload_0_2893);
  assign _zz_dataOut_payload_0_3592 = (_zz_dataOut_payload_0_3590 ? _zz_dataOut_payload_0_2893 : _zz_dataOut_payload_0_2882);
  assign _zz_dataOut_payload_0_3593 = (_zz_dataOut_payload_0_2883 < _zz_dataOut_payload_0_2892);
  assign _zz_dataOut_payload_0_3594 = (_zz_dataOut_payload_0_3593 ? _zz_dataOut_payload_0_2883 : _zz_dataOut_payload_0_2892);
  assign _zz_dataOut_payload_0_3595 = (_zz_dataOut_payload_0_3593 ? _zz_dataOut_payload_0_2892 : _zz_dataOut_payload_0_2883);
  assign _zz_dataOut_payload_0_3596 = (_zz_dataOut_payload_0_2884 < _zz_dataOut_payload_0_2891);
  assign _zz_dataOut_payload_0_3597 = (_zz_dataOut_payload_0_3596 ? _zz_dataOut_payload_0_2884 : _zz_dataOut_payload_0_2891);
  assign _zz_dataOut_payload_0_3598 = (_zz_dataOut_payload_0_3596 ? _zz_dataOut_payload_0_2891 : _zz_dataOut_payload_0_2884);
  assign _zz_dataOut_payload_0_3599 = (_zz_dataOut_payload_0_2885 < _zz_dataOut_payload_0_2890);
  assign _zz_dataOut_payload_0_3600 = (_zz_dataOut_payload_0_3599 ? _zz_dataOut_payload_0_2885 : _zz_dataOut_payload_0_2890);
  assign _zz_dataOut_payload_0_3601 = (_zz_dataOut_payload_0_3599 ? _zz_dataOut_payload_0_2890 : _zz_dataOut_payload_0_2885);
  assign _zz_dataOut_payload_0_3602 = (_zz_dataOut_payload_0_2886 < _zz_dataOut_payload_0_2889);
  assign _zz_dataOut_payload_0_3603 = (_zz_dataOut_payload_0_3602 ? _zz_dataOut_payload_0_2886 : _zz_dataOut_payload_0_2889);
  assign _zz_dataOut_payload_0_3604 = (_zz_dataOut_payload_0_3602 ? _zz_dataOut_payload_0_2889 : _zz_dataOut_payload_0_2886);
  assign _zz_dataOut_payload_0_3605 = (_zz_dataOut_payload_0_2887 < _zz_dataOut_payload_0_2888);
  assign _zz_dataOut_payload_0_3606 = (_zz_dataOut_payload_0_3605 ? _zz_dataOut_payload_0_2887 : _zz_dataOut_payload_0_2888);
  assign _zz_dataOut_payload_0_3607 = (_zz_dataOut_payload_0_3605 ? _zz_dataOut_payload_0_2888 : _zz_dataOut_payload_0_2887);
  assign _zz_dataOut_payload_0_3608 = (_zz_dataOut_payload_0_3585 < _zz_dataOut_payload_0_3597);
  assign _zz_dataOut_payload_0_3609 = (_zz_dataOut_payload_0_3608 ? _zz_dataOut_payload_0_3585 : _zz_dataOut_payload_0_3597);
  assign _zz_dataOut_payload_0_3610 = (_zz_dataOut_payload_0_3608 ? _zz_dataOut_payload_0_3597 : _zz_dataOut_payload_0_3585);
  assign _zz_dataOut_payload_0_3611 = (_zz_dataOut_payload_0_3588 < _zz_dataOut_payload_0_3600);
  assign _zz_dataOut_payload_0_3612 = (_zz_dataOut_payload_0_3611 ? _zz_dataOut_payload_0_3588 : _zz_dataOut_payload_0_3600);
  assign _zz_dataOut_payload_0_3613 = (_zz_dataOut_payload_0_3611 ? _zz_dataOut_payload_0_3600 : _zz_dataOut_payload_0_3588);
  assign _zz_dataOut_payload_0_3614 = (_zz_dataOut_payload_0_3591 < _zz_dataOut_payload_0_3603);
  assign _zz_dataOut_payload_0_3615 = (_zz_dataOut_payload_0_3614 ? _zz_dataOut_payload_0_3591 : _zz_dataOut_payload_0_3603);
  assign _zz_dataOut_payload_0_3616 = (_zz_dataOut_payload_0_3614 ? _zz_dataOut_payload_0_3603 : _zz_dataOut_payload_0_3591);
  assign _zz_dataOut_payload_0_3617 = (_zz_dataOut_payload_0_3594 < _zz_dataOut_payload_0_3606);
  assign _zz_dataOut_payload_0_3618 = (_zz_dataOut_payload_0_3617 ? _zz_dataOut_payload_0_3594 : _zz_dataOut_payload_0_3606);
  assign _zz_dataOut_payload_0_3619 = (_zz_dataOut_payload_0_3617 ? _zz_dataOut_payload_0_3606 : _zz_dataOut_payload_0_3594);
  assign _zz_dataOut_payload_0_3620 = (_zz_dataOut_payload_0_3609 < _zz_dataOut_payload_0_3615);
  assign _zz_dataOut_payload_0_3621 = (_zz_dataOut_payload_0_3620 ? _zz_dataOut_payload_0_3609 : _zz_dataOut_payload_0_3615);
  assign _zz_dataOut_payload_0_3622 = (_zz_dataOut_payload_0_3620 ? _zz_dataOut_payload_0_3615 : _zz_dataOut_payload_0_3609);
  assign _zz_dataOut_payload_0_3623 = (_zz_dataOut_payload_0_3612 < _zz_dataOut_payload_0_3618);
  assign _zz_dataOut_payload_0_3624 = (_zz_dataOut_payload_0_3623 ? _zz_dataOut_payload_0_3612 : _zz_dataOut_payload_0_3618);
  assign _zz_dataOut_payload_0_3625 = (_zz_dataOut_payload_0_3623 ? _zz_dataOut_payload_0_3618 : _zz_dataOut_payload_0_3612);
  assign _zz_dataOut_payload_0_3626 = (_zz_dataOut_payload_0_3621 < _zz_dataOut_payload_0_3624);
  assign _zz_dataOut_payload_0_3627 = (_zz_dataOut_payload_0_3622 < _zz_dataOut_payload_0_3625);
  assign _zz_dataOut_payload_0_3632 = (_zz_dataOut_payload_0_3610 < _zz_dataOut_payload_0_3616);
  assign _zz_dataOut_payload_0_3633 = (_zz_dataOut_payload_0_3632 ? _zz_dataOut_payload_0_3610 : _zz_dataOut_payload_0_3616);
  assign _zz_dataOut_payload_0_3634 = (_zz_dataOut_payload_0_3632 ? _zz_dataOut_payload_0_3616 : _zz_dataOut_payload_0_3610);
  assign _zz_dataOut_payload_0_3635 = (_zz_dataOut_payload_0_3613 < _zz_dataOut_payload_0_3619);
  assign _zz_dataOut_payload_0_3636 = (_zz_dataOut_payload_0_3635 ? _zz_dataOut_payload_0_3613 : _zz_dataOut_payload_0_3619);
  assign _zz_dataOut_payload_0_3637 = (_zz_dataOut_payload_0_3635 ? _zz_dataOut_payload_0_3619 : _zz_dataOut_payload_0_3613);
  assign _zz_dataOut_payload_0_3638 = (_zz_dataOut_payload_0_3633 < _zz_dataOut_payload_0_3636);
  assign _zz_dataOut_payload_0_3639 = (_zz_dataOut_payload_0_3634 < _zz_dataOut_payload_0_3637);
  assign _zz_dataOut_payload_0_3652 = (_zz_dataOut_payload_0_3607 < _zz_dataOut_payload_0_3595);
  assign _zz_dataOut_payload_0_3653 = (_zz_dataOut_payload_0_3652 ? _zz_dataOut_payload_0_3607 : _zz_dataOut_payload_0_3595);
  assign _zz_dataOut_payload_0_3654 = (_zz_dataOut_payload_0_3652 ? _zz_dataOut_payload_0_3595 : _zz_dataOut_payload_0_3607);
  assign _zz_dataOut_payload_0_3655 = (_zz_dataOut_payload_0_3604 < _zz_dataOut_payload_0_3592);
  assign _zz_dataOut_payload_0_3656 = (_zz_dataOut_payload_0_3655 ? _zz_dataOut_payload_0_3604 : _zz_dataOut_payload_0_3592);
  assign _zz_dataOut_payload_0_3657 = (_zz_dataOut_payload_0_3655 ? _zz_dataOut_payload_0_3592 : _zz_dataOut_payload_0_3604);
  assign _zz_dataOut_payload_0_3658 = (_zz_dataOut_payload_0_3601 < _zz_dataOut_payload_0_3589);
  assign _zz_dataOut_payload_0_3659 = (_zz_dataOut_payload_0_3658 ? _zz_dataOut_payload_0_3601 : _zz_dataOut_payload_0_3589);
  assign _zz_dataOut_payload_0_3660 = (_zz_dataOut_payload_0_3658 ? _zz_dataOut_payload_0_3589 : _zz_dataOut_payload_0_3601);
  assign _zz_dataOut_payload_0_3661 = (_zz_dataOut_payload_0_3598 < _zz_dataOut_payload_0_3586);
  assign _zz_dataOut_payload_0_3662 = (_zz_dataOut_payload_0_3661 ? _zz_dataOut_payload_0_3598 : _zz_dataOut_payload_0_3586);
  assign _zz_dataOut_payload_0_3663 = (_zz_dataOut_payload_0_3661 ? _zz_dataOut_payload_0_3586 : _zz_dataOut_payload_0_3598);
  assign _zz_dataOut_payload_0_3664 = (_zz_dataOut_payload_0_3653 < _zz_dataOut_payload_0_3659);
  assign _zz_dataOut_payload_0_3665 = (_zz_dataOut_payload_0_3664 ? _zz_dataOut_payload_0_3653 : _zz_dataOut_payload_0_3659);
  assign _zz_dataOut_payload_0_3666 = (_zz_dataOut_payload_0_3664 ? _zz_dataOut_payload_0_3659 : _zz_dataOut_payload_0_3653);
  assign _zz_dataOut_payload_0_3667 = (_zz_dataOut_payload_0_3656 < _zz_dataOut_payload_0_3662);
  assign _zz_dataOut_payload_0_3668 = (_zz_dataOut_payload_0_3667 ? _zz_dataOut_payload_0_3656 : _zz_dataOut_payload_0_3662);
  assign _zz_dataOut_payload_0_3669 = (_zz_dataOut_payload_0_3667 ? _zz_dataOut_payload_0_3662 : _zz_dataOut_payload_0_3656);
  assign _zz_dataOut_payload_0_3670 = (_zz_dataOut_payload_0_3665 < _zz_dataOut_payload_0_3668);
  assign _zz_dataOut_payload_0_3671 = (_zz_dataOut_payload_0_3666 < _zz_dataOut_payload_0_3669);
  assign _zz_dataOut_payload_0_3676 = (_zz_dataOut_payload_0_3654 < _zz_dataOut_payload_0_3660);
  assign _zz_dataOut_payload_0_3677 = (_zz_dataOut_payload_0_3676 ? _zz_dataOut_payload_0_3654 : _zz_dataOut_payload_0_3660);
  assign _zz_dataOut_payload_0_3678 = (_zz_dataOut_payload_0_3676 ? _zz_dataOut_payload_0_3660 : _zz_dataOut_payload_0_3654);
  assign _zz_dataOut_payload_0_3679 = (_zz_dataOut_payload_0_3657 < _zz_dataOut_payload_0_3663);
  assign _zz_dataOut_payload_0_3680 = (_zz_dataOut_payload_0_3679 ? _zz_dataOut_payload_0_3657 : _zz_dataOut_payload_0_3663);
  assign _zz_dataOut_payload_0_3681 = (_zz_dataOut_payload_0_3679 ? _zz_dataOut_payload_0_3663 : _zz_dataOut_payload_0_3657);
  assign _zz_dataOut_payload_0_3682 = (_zz_dataOut_payload_0_3677 < _zz_dataOut_payload_0_3680);
  assign _zz_dataOut_payload_0_3683 = (_zz_dataOut_payload_0_3678 < _zz_dataOut_payload_0_3681);
  assign _zz_dataOut_payload_0_3712 = (_zz_dataOut_payload_0_2896 < _zz_dataOut_payload_0_2911);
  assign _zz_dataOut_payload_0_3713 = (_zz_dataOut_payload_0_3712 ? _zz_dataOut_payload_0_2896 : _zz_dataOut_payload_0_2911);
  assign _zz_dataOut_payload_0_3714 = (_zz_dataOut_payload_0_3712 ? _zz_dataOut_payload_0_2911 : _zz_dataOut_payload_0_2896);
  assign _zz_dataOut_payload_0_3715 = (_zz_dataOut_payload_0_2897 < _zz_dataOut_payload_0_2910);
  assign _zz_dataOut_payload_0_3716 = (_zz_dataOut_payload_0_3715 ? _zz_dataOut_payload_0_2897 : _zz_dataOut_payload_0_2910);
  assign _zz_dataOut_payload_0_3717 = (_zz_dataOut_payload_0_3715 ? _zz_dataOut_payload_0_2910 : _zz_dataOut_payload_0_2897);
  assign _zz_dataOut_payload_0_3718 = (_zz_dataOut_payload_0_2898 < _zz_dataOut_payload_0_2909);
  assign _zz_dataOut_payload_0_3719 = (_zz_dataOut_payload_0_3718 ? _zz_dataOut_payload_0_2898 : _zz_dataOut_payload_0_2909);
  assign _zz_dataOut_payload_0_3720 = (_zz_dataOut_payload_0_3718 ? _zz_dataOut_payload_0_2909 : _zz_dataOut_payload_0_2898);
  assign _zz_dataOut_payload_0_3721 = (_zz_dataOut_payload_0_2899 < _zz_dataOut_payload_0_2908);
  assign _zz_dataOut_payload_0_3722 = (_zz_dataOut_payload_0_3721 ? _zz_dataOut_payload_0_2899 : _zz_dataOut_payload_0_2908);
  assign _zz_dataOut_payload_0_3723 = (_zz_dataOut_payload_0_3721 ? _zz_dataOut_payload_0_2908 : _zz_dataOut_payload_0_2899);
  assign _zz_dataOut_payload_0_3724 = (_zz_dataOut_payload_0_2900 < _zz_dataOut_payload_0_2907);
  assign _zz_dataOut_payload_0_3725 = (_zz_dataOut_payload_0_3724 ? _zz_dataOut_payload_0_2900 : _zz_dataOut_payload_0_2907);
  assign _zz_dataOut_payload_0_3726 = (_zz_dataOut_payload_0_3724 ? _zz_dataOut_payload_0_2907 : _zz_dataOut_payload_0_2900);
  assign _zz_dataOut_payload_0_3727 = (_zz_dataOut_payload_0_2901 < _zz_dataOut_payload_0_2906);
  assign _zz_dataOut_payload_0_3728 = (_zz_dataOut_payload_0_3727 ? _zz_dataOut_payload_0_2901 : _zz_dataOut_payload_0_2906);
  assign _zz_dataOut_payload_0_3729 = (_zz_dataOut_payload_0_3727 ? _zz_dataOut_payload_0_2906 : _zz_dataOut_payload_0_2901);
  assign _zz_dataOut_payload_0_3730 = (_zz_dataOut_payload_0_2902 < _zz_dataOut_payload_0_2905);
  assign _zz_dataOut_payload_0_3731 = (_zz_dataOut_payload_0_3730 ? _zz_dataOut_payload_0_2902 : _zz_dataOut_payload_0_2905);
  assign _zz_dataOut_payload_0_3732 = (_zz_dataOut_payload_0_3730 ? _zz_dataOut_payload_0_2905 : _zz_dataOut_payload_0_2902);
  assign _zz_dataOut_payload_0_3733 = (_zz_dataOut_payload_0_2903 < _zz_dataOut_payload_0_2904);
  assign _zz_dataOut_payload_0_3734 = (_zz_dataOut_payload_0_3733 ? _zz_dataOut_payload_0_2903 : _zz_dataOut_payload_0_2904);
  assign _zz_dataOut_payload_0_3735 = (_zz_dataOut_payload_0_3733 ? _zz_dataOut_payload_0_2904 : _zz_dataOut_payload_0_2903);
  assign _zz_dataOut_payload_0_3736 = (_zz_dataOut_payload_0_3713 < _zz_dataOut_payload_0_3725);
  assign _zz_dataOut_payload_0_3737 = (_zz_dataOut_payload_0_3736 ? _zz_dataOut_payload_0_3713 : _zz_dataOut_payload_0_3725);
  assign _zz_dataOut_payload_0_3738 = (_zz_dataOut_payload_0_3736 ? _zz_dataOut_payload_0_3725 : _zz_dataOut_payload_0_3713);
  assign _zz_dataOut_payload_0_3739 = (_zz_dataOut_payload_0_3716 < _zz_dataOut_payload_0_3728);
  assign _zz_dataOut_payload_0_3740 = (_zz_dataOut_payload_0_3739 ? _zz_dataOut_payload_0_3716 : _zz_dataOut_payload_0_3728);
  assign _zz_dataOut_payload_0_3741 = (_zz_dataOut_payload_0_3739 ? _zz_dataOut_payload_0_3728 : _zz_dataOut_payload_0_3716);
  assign _zz_dataOut_payload_0_3742 = (_zz_dataOut_payload_0_3719 < _zz_dataOut_payload_0_3731);
  assign _zz_dataOut_payload_0_3743 = (_zz_dataOut_payload_0_3742 ? _zz_dataOut_payload_0_3719 : _zz_dataOut_payload_0_3731);
  assign _zz_dataOut_payload_0_3744 = (_zz_dataOut_payload_0_3742 ? _zz_dataOut_payload_0_3731 : _zz_dataOut_payload_0_3719);
  assign _zz_dataOut_payload_0_3745 = (_zz_dataOut_payload_0_3722 < _zz_dataOut_payload_0_3734);
  assign _zz_dataOut_payload_0_3746 = (_zz_dataOut_payload_0_3745 ? _zz_dataOut_payload_0_3722 : _zz_dataOut_payload_0_3734);
  assign _zz_dataOut_payload_0_3747 = (_zz_dataOut_payload_0_3745 ? _zz_dataOut_payload_0_3734 : _zz_dataOut_payload_0_3722);
  assign _zz_dataOut_payload_0_3748 = (_zz_dataOut_payload_0_3737 < _zz_dataOut_payload_0_3743);
  assign _zz_dataOut_payload_0_3749 = (_zz_dataOut_payload_0_3748 ? _zz_dataOut_payload_0_3737 : _zz_dataOut_payload_0_3743);
  assign _zz_dataOut_payload_0_3750 = (_zz_dataOut_payload_0_3748 ? _zz_dataOut_payload_0_3743 : _zz_dataOut_payload_0_3737);
  assign _zz_dataOut_payload_0_3751 = (_zz_dataOut_payload_0_3740 < _zz_dataOut_payload_0_3746);
  assign _zz_dataOut_payload_0_3752 = (_zz_dataOut_payload_0_3751 ? _zz_dataOut_payload_0_3740 : _zz_dataOut_payload_0_3746);
  assign _zz_dataOut_payload_0_3753 = (_zz_dataOut_payload_0_3751 ? _zz_dataOut_payload_0_3746 : _zz_dataOut_payload_0_3740);
  assign _zz_dataOut_payload_0_3754 = (_zz_dataOut_payload_0_3749 < _zz_dataOut_payload_0_3752);
  assign _zz_dataOut_payload_0_3755 = (_zz_dataOut_payload_0_3750 < _zz_dataOut_payload_0_3753);
  assign _zz_dataOut_payload_0_3760 = (_zz_dataOut_payload_0_3738 < _zz_dataOut_payload_0_3744);
  assign _zz_dataOut_payload_0_3761 = (_zz_dataOut_payload_0_3760 ? _zz_dataOut_payload_0_3738 : _zz_dataOut_payload_0_3744);
  assign _zz_dataOut_payload_0_3762 = (_zz_dataOut_payload_0_3760 ? _zz_dataOut_payload_0_3744 : _zz_dataOut_payload_0_3738);
  assign _zz_dataOut_payload_0_3763 = (_zz_dataOut_payload_0_3741 < _zz_dataOut_payload_0_3747);
  assign _zz_dataOut_payload_0_3764 = (_zz_dataOut_payload_0_3763 ? _zz_dataOut_payload_0_3741 : _zz_dataOut_payload_0_3747);
  assign _zz_dataOut_payload_0_3765 = (_zz_dataOut_payload_0_3763 ? _zz_dataOut_payload_0_3747 : _zz_dataOut_payload_0_3741);
  assign _zz_dataOut_payload_0_3766 = (_zz_dataOut_payload_0_3761 < _zz_dataOut_payload_0_3764);
  assign _zz_dataOut_payload_0_3767 = (_zz_dataOut_payload_0_3762 < _zz_dataOut_payload_0_3765);
  assign _zz_dataOut_payload_0_3780 = (_zz_dataOut_payload_0_3735 < _zz_dataOut_payload_0_3723);
  assign _zz_dataOut_payload_0_3781 = (_zz_dataOut_payload_0_3780 ? _zz_dataOut_payload_0_3735 : _zz_dataOut_payload_0_3723);
  assign _zz_dataOut_payload_0_3782 = (_zz_dataOut_payload_0_3780 ? _zz_dataOut_payload_0_3723 : _zz_dataOut_payload_0_3735);
  assign _zz_dataOut_payload_0_3783 = (_zz_dataOut_payload_0_3732 < _zz_dataOut_payload_0_3720);
  assign _zz_dataOut_payload_0_3784 = (_zz_dataOut_payload_0_3783 ? _zz_dataOut_payload_0_3732 : _zz_dataOut_payload_0_3720);
  assign _zz_dataOut_payload_0_3785 = (_zz_dataOut_payload_0_3783 ? _zz_dataOut_payload_0_3720 : _zz_dataOut_payload_0_3732);
  assign _zz_dataOut_payload_0_3786 = (_zz_dataOut_payload_0_3729 < _zz_dataOut_payload_0_3717);
  assign _zz_dataOut_payload_0_3787 = (_zz_dataOut_payload_0_3786 ? _zz_dataOut_payload_0_3729 : _zz_dataOut_payload_0_3717);
  assign _zz_dataOut_payload_0_3788 = (_zz_dataOut_payload_0_3786 ? _zz_dataOut_payload_0_3717 : _zz_dataOut_payload_0_3729);
  assign _zz_dataOut_payload_0_3789 = (_zz_dataOut_payload_0_3726 < _zz_dataOut_payload_0_3714);
  assign _zz_dataOut_payload_0_3790 = (_zz_dataOut_payload_0_3789 ? _zz_dataOut_payload_0_3726 : _zz_dataOut_payload_0_3714);
  assign _zz_dataOut_payload_0_3791 = (_zz_dataOut_payload_0_3789 ? _zz_dataOut_payload_0_3714 : _zz_dataOut_payload_0_3726);
  assign _zz_dataOut_payload_0_3792 = (_zz_dataOut_payload_0_3781 < _zz_dataOut_payload_0_3787);
  assign _zz_dataOut_payload_0_3793 = (_zz_dataOut_payload_0_3792 ? _zz_dataOut_payload_0_3781 : _zz_dataOut_payload_0_3787);
  assign _zz_dataOut_payload_0_3794 = (_zz_dataOut_payload_0_3792 ? _zz_dataOut_payload_0_3787 : _zz_dataOut_payload_0_3781);
  assign _zz_dataOut_payload_0_3795 = (_zz_dataOut_payload_0_3784 < _zz_dataOut_payload_0_3790);
  assign _zz_dataOut_payload_0_3796 = (_zz_dataOut_payload_0_3795 ? _zz_dataOut_payload_0_3784 : _zz_dataOut_payload_0_3790);
  assign _zz_dataOut_payload_0_3797 = (_zz_dataOut_payload_0_3795 ? _zz_dataOut_payload_0_3790 : _zz_dataOut_payload_0_3784);
  assign _zz_dataOut_payload_0_3798 = (_zz_dataOut_payload_0_3793 < _zz_dataOut_payload_0_3796);
  assign _zz_dataOut_payload_0_3799 = (_zz_dataOut_payload_0_3794 < _zz_dataOut_payload_0_3797);
  assign _zz_dataOut_payload_0_3804 = (_zz_dataOut_payload_0_3782 < _zz_dataOut_payload_0_3788);
  assign _zz_dataOut_payload_0_3805 = (_zz_dataOut_payload_0_3804 ? _zz_dataOut_payload_0_3782 : _zz_dataOut_payload_0_3788);
  assign _zz_dataOut_payload_0_3806 = (_zz_dataOut_payload_0_3804 ? _zz_dataOut_payload_0_3788 : _zz_dataOut_payload_0_3782);
  assign _zz_dataOut_payload_0_3807 = (_zz_dataOut_payload_0_3785 < _zz_dataOut_payload_0_3791);
  assign _zz_dataOut_payload_0_3808 = (_zz_dataOut_payload_0_3807 ? _zz_dataOut_payload_0_3785 : _zz_dataOut_payload_0_3791);
  assign _zz_dataOut_payload_0_3809 = (_zz_dataOut_payload_0_3807 ? _zz_dataOut_payload_0_3791 : _zz_dataOut_payload_0_3785);
  assign _zz_dataOut_payload_0_3810 = (_zz_dataOut_payload_0_3805 < _zz_dataOut_payload_0_3808);
  assign _zz_dataOut_payload_0_3811 = (_zz_dataOut_payload_0_3806 < _zz_dataOut_payload_0_3809);
  assign _zz_dataOut_payload_0_3840 = (_zz_dataOut_payload_0_2912 < _zz_dataOut_payload_0_2927);
  assign _zz_dataOut_payload_0_3841 = (_zz_dataOut_payload_0_3840 ? _zz_dataOut_payload_0_2912 : _zz_dataOut_payload_0_2927);
  assign _zz_dataOut_payload_0_3842 = (_zz_dataOut_payload_0_3840 ? _zz_dataOut_payload_0_2927 : _zz_dataOut_payload_0_2912);
  assign _zz_dataOut_payload_0_3843 = (_zz_dataOut_payload_0_2913 < _zz_dataOut_payload_0_2926);
  assign _zz_dataOut_payload_0_3844 = (_zz_dataOut_payload_0_3843 ? _zz_dataOut_payload_0_2913 : _zz_dataOut_payload_0_2926);
  assign _zz_dataOut_payload_0_3845 = (_zz_dataOut_payload_0_3843 ? _zz_dataOut_payload_0_2926 : _zz_dataOut_payload_0_2913);
  assign _zz_dataOut_payload_0_3846 = (_zz_dataOut_payload_0_2914 < _zz_dataOut_payload_0_2925);
  assign _zz_dataOut_payload_0_3847 = (_zz_dataOut_payload_0_3846 ? _zz_dataOut_payload_0_2914 : _zz_dataOut_payload_0_2925);
  assign _zz_dataOut_payload_0_3848 = (_zz_dataOut_payload_0_3846 ? _zz_dataOut_payload_0_2925 : _zz_dataOut_payload_0_2914);
  assign _zz_dataOut_payload_0_3849 = (_zz_dataOut_payload_0_2915 < _zz_dataOut_payload_0_2924);
  assign _zz_dataOut_payload_0_3850 = (_zz_dataOut_payload_0_3849 ? _zz_dataOut_payload_0_2915 : _zz_dataOut_payload_0_2924);
  assign _zz_dataOut_payload_0_3851 = (_zz_dataOut_payload_0_3849 ? _zz_dataOut_payload_0_2924 : _zz_dataOut_payload_0_2915);
  assign _zz_dataOut_payload_0_3852 = (_zz_dataOut_payload_0_2916 < _zz_dataOut_payload_0_2923);
  assign _zz_dataOut_payload_0_3853 = (_zz_dataOut_payload_0_3852 ? _zz_dataOut_payload_0_2916 : _zz_dataOut_payload_0_2923);
  assign _zz_dataOut_payload_0_3854 = (_zz_dataOut_payload_0_3852 ? _zz_dataOut_payload_0_2923 : _zz_dataOut_payload_0_2916);
  assign _zz_dataOut_payload_0_3855 = (_zz_dataOut_payload_0_2917 < _zz_dataOut_payload_0_2922);
  assign _zz_dataOut_payload_0_3856 = (_zz_dataOut_payload_0_3855 ? _zz_dataOut_payload_0_2917 : _zz_dataOut_payload_0_2922);
  assign _zz_dataOut_payload_0_3857 = (_zz_dataOut_payload_0_3855 ? _zz_dataOut_payload_0_2922 : _zz_dataOut_payload_0_2917);
  assign _zz_dataOut_payload_0_3858 = (_zz_dataOut_payload_0_2918 < _zz_dataOut_payload_0_2921);
  assign _zz_dataOut_payload_0_3859 = (_zz_dataOut_payload_0_3858 ? _zz_dataOut_payload_0_2918 : _zz_dataOut_payload_0_2921);
  assign _zz_dataOut_payload_0_3860 = (_zz_dataOut_payload_0_3858 ? _zz_dataOut_payload_0_2921 : _zz_dataOut_payload_0_2918);
  assign _zz_dataOut_payload_0_3861 = (_zz_dataOut_payload_0_2919 < _zz_dataOut_payload_0_2920);
  assign _zz_dataOut_payload_0_3862 = (_zz_dataOut_payload_0_3861 ? _zz_dataOut_payload_0_2919 : _zz_dataOut_payload_0_2920);
  assign _zz_dataOut_payload_0_3863 = (_zz_dataOut_payload_0_3861 ? _zz_dataOut_payload_0_2920 : _zz_dataOut_payload_0_2919);
  assign _zz_dataOut_payload_0_3864 = (_zz_dataOut_payload_0_3841 < _zz_dataOut_payload_0_3853);
  assign _zz_dataOut_payload_0_3865 = (_zz_dataOut_payload_0_3864 ? _zz_dataOut_payload_0_3841 : _zz_dataOut_payload_0_3853);
  assign _zz_dataOut_payload_0_3866 = (_zz_dataOut_payload_0_3864 ? _zz_dataOut_payload_0_3853 : _zz_dataOut_payload_0_3841);
  assign _zz_dataOut_payload_0_3867 = (_zz_dataOut_payload_0_3844 < _zz_dataOut_payload_0_3856);
  assign _zz_dataOut_payload_0_3868 = (_zz_dataOut_payload_0_3867 ? _zz_dataOut_payload_0_3844 : _zz_dataOut_payload_0_3856);
  assign _zz_dataOut_payload_0_3869 = (_zz_dataOut_payload_0_3867 ? _zz_dataOut_payload_0_3856 : _zz_dataOut_payload_0_3844);
  assign _zz_dataOut_payload_0_3870 = (_zz_dataOut_payload_0_3847 < _zz_dataOut_payload_0_3859);
  assign _zz_dataOut_payload_0_3871 = (_zz_dataOut_payload_0_3870 ? _zz_dataOut_payload_0_3847 : _zz_dataOut_payload_0_3859);
  assign _zz_dataOut_payload_0_3872 = (_zz_dataOut_payload_0_3870 ? _zz_dataOut_payload_0_3859 : _zz_dataOut_payload_0_3847);
  assign _zz_dataOut_payload_0_3873 = (_zz_dataOut_payload_0_3850 < _zz_dataOut_payload_0_3862);
  assign _zz_dataOut_payload_0_3874 = (_zz_dataOut_payload_0_3873 ? _zz_dataOut_payload_0_3850 : _zz_dataOut_payload_0_3862);
  assign _zz_dataOut_payload_0_3875 = (_zz_dataOut_payload_0_3873 ? _zz_dataOut_payload_0_3862 : _zz_dataOut_payload_0_3850);
  assign _zz_dataOut_payload_0_3876 = (_zz_dataOut_payload_0_3865 < _zz_dataOut_payload_0_3871);
  assign _zz_dataOut_payload_0_3877 = (_zz_dataOut_payload_0_3876 ? _zz_dataOut_payload_0_3865 : _zz_dataOut_payload_0_3871);
  assign _zz_dataOut_payload_0_3878 = (_zz_dataOut_payload_0_3876 ? _zz_dataOut_payload_0_3871 : _zz_dataOut_payload_0_3865);
  assign _zz_dataOut_payload_0_3879 = (_zz_dataOut_payload_0_3868 < _zz_dataOut_payload_0_3874);
  assign _zz_dataOut_payload_0_3880 = (_zz_dataOut_payload_0_3879 ? _zz_dataOut_payload_0_3868 : _zz_dataOut_payload_0_3874);
  assign _zz_dataOut_payload_0_3881 = (_zz_dataOut_payload_0_3879 ? _zz_dataOut_payload_0_3874 : _zz_dataOut_payload_0_3868);
  assign _zz_dataOut_payload_0_3882 = (_zz_dataOut_payload_0_3877 < _zz_dataOut_payload_0_3880);
  assign _zz_dataOut_payload_0_3883 = (_zz_dataOut_payload_0_3878 < _zz_dataOut_payload_0_3881);
  assign _zz_dataOut_payload_0_3888 = (_zz_dataOut_payload_0_3866 < _zz_dataOut_payload_0_3872);
  assign _zz_dataOut_payload_0_3889 = (_zz_dataOut_payload_0_3888 ? _zz_dataOut_payload_0_3866 : _zz_dataOut_payload_0_3872);
  assign _zz_dataOut_payload_0_3890 = (_zz_dataOut_payload_0_3888 ? _zz_dataOut_payload_0_3872 : _zz_dataOut_payload_0_3866);
  assign _zz_dataOut_payload_0_3891 = (_zz_dataOut_payload_0_3869 < _zz_dataOut_payload_0_3875);
  assign _zz_dataOut_payload_0_3892 = (_zz_dataOut_payload_0_3891 ? _zz_dataOut_payload_0_3869 : _zz_dataOut_payload_0_3875);
  assign _zz_dataOut_payload_0_3893 = (_zz_dataOut_payload_0_3891 ? _zz_dataOut_payload_0_3875 : _zz_dataOut_payload_0_3869);
  assign _zz_dataOut_payload_0_3894 = (_zz_dataOut_payload_0_3889 < _zz_dataOut_payload_0_3892);
  assign _zz_dataOut_payload_0_3895 = (_zz_dataOut_payload_0_3890 < _zz_dataOut_payload_0_3893);
  assign _zz_dataOut_payload_0_3908 = (_zz_dataOut_payload_0_3863 < _zz_dataOut_payload_0_3851);
  assign _zz_dataOut_payload_0_3909 = (_zz_dataOut_payload_0_3908 ? _zz_dataOut_payload_0_3863 : _zz_dataOut_payload_0_3851);
  assign _zz_dataOut_payload_0_3910 = (_zz_dataOut_payload_0_3908 ? _zz_dataOut_payload_0_3851 : _zz_dataOut_payload_0_3863);
  assign _zz_dataOut_payload_0_3911 = (_zz_dataOut_payload_0_3860 < _zz_dataOut_payload_0_3848);
  assign _zz_dataOut_payload_0_3912 = (_zz_dataOut_payload_0_3911 ? _zz_dataOut_payload_0_3860 : _zz_dataOut_payload_0_3848);
  assign _zz_dataOut_payload_0_3913 = (_zz_dataOut_payload_0_3911 ? _zz_dataOut_payload_0_3848 : _zz_dataOut_payload_0_3860);
  assign _zz_dataOut_payload_0_3914 = (_zz_dataOut_payload_0_3857 < _zz_dataOut_payload_0_3845);
  assign _zz_dataOut_payload_0_3915 = (_zz_dataOut_payload_0_3914 ? _zz_dataOut_payload_0_3857 : _zz_dataOut_payload_0_3845);
  assign _zz_dataOut_payload_0_3916 = (_zz_dataOut_payload_0_3914 ? _zz_dataOut_payload_0_3845 : _zz_dataOut_payload_0_3857);
  assign _zz_dataOut_payload_0_3917 = (_zz_dataOut_payload_0_3854 < _zz_dataOut_payload_0_3842);
  assign _zz_dataOut_payload_0_3918 = (_zz_dataOut_payload_0_3917 ? _zz_dataOut_payload_0_3854 : _zz_dataOut_payload_0_3842);
  assign _zz_dataOut_payload_0_3919 = (_zz_dataOut_payload_0_3917 ? _zz_dataOut_payload_0_3842 : _zz_dataOut_payload_0_3854);
  assign _zz_dataOut_payload_0_3920 = (_zz_dataOut_payload_0_3909 < _zz_dataOut_payload_0_3915);
  assign _zz_dataOut_payload_0_3921 = (_zz_dataOut_payload_0_3920 ? _zz_dataOut_payload_0_3909 : _zz_dataOut_payload_0_3915);
  assign _zz_dataOut_payload_0_3922 = (_zz_dataOut_payload_0_3920 ? _zz_dataOut_payload_0_3915 : _zz_dataOut_payload_0_3909);
  assign _zz_dataOut_payload_0_3923 = (_zz_dataOut_payload_0_3912 < _zz_dataOut_payload_0_3918);
  assign _zz_dataOut_payload_0_3924 = (_zz_dataOut_payload_0_3923 ? _zz_dataOut_payload_0_3912 : _zz_dataOut_payload_0_3918);
  assign _zz_dataOut_payload_0_3925 = (_zz_dataOut_payload_0_3923 ? _zz_dataOut_payload_0_3918 : _zz_dataOut_payload_0_3912);
  assign _zz_dataOut_payload_0_3926 = (_zz_dataOut_payload_0_3921 < _zz_dataOut_payload_0_3924);
  assign _zz_dataOut_payload_0_3927 = (_zz_dataOut_payload_0_3922 < _zz_dataOut_payload_0_3925);
  assign _zz_dataOut_payload_0_3932 = (_zz_dataOut_payload_0_3910 < _zz_dataOut_payload_0_3916);
  assign _zz_dataOut_payload_0_3933 = (_zz_dataOut_payload_0_3932 ? _zz_dataOut_payload_0_3910 : _zz_dataOut_payload_0_3916);
  assign _zz_dataOut_payload_0_3934 = (_zz_dataOut_payload_0_3932 ? _zz_dataOut_payload_0_3916 : _zz_dataOut_payload_0_3910);
  assign _zz_dataOut_payload_0_3935 = (_zz_dataOut_payload_0_3913 < _zz_dataOut_payload_0_3919);
  assign _zz_dataOut_payload_0_3936 = (_zz_dataOut_payload_0_3935 ? _zz_dataOut_payload_0_3913 : _zz_dataOut_payload_0_3919);
  assign _zz_dataOut_payload_0_3937 = (_zz_dataOut_payload_0_3935 ? _zz_dataOut_payload_0_3919 : _zz_dataOut_payload_0_3913);
  assign _zz_dataOut_payload_0_3938 = (_zz_dataOut_payload_0_3933 < _zz_dataOut_payload_0_3936);
  assign _zz_dataOut_payload_0_3939 = (_zz_dataOut_payload_0_3934 < _zz_dataOut_payload_0_3937);
  assign _zz_dataOut_payload_0_3968 = (_zz_dataOut_payload_0_2928 < _zz_dataOut_payload_0_2943);
  assign _zz_dataOut_payload_0_3969 = (_zz_dataOut_payload_0_3968 ? _zz_dataOut_payload_0_2928 : _zz_dataOut_payload_0_2943);
  assign _zz_dataOut_payload_0_3970 = (_zz_dataOut_payload_0_3968 ? _zz_dataOut_payload_0_2943 : _zz_dataOut_payload_0_2928);
  assign _zz_dataOut_payload_0_3971 = (_zz_dataOut_payload_0_2929 < _zz_dataOut_payload_0_2942);
  assign _zz_dataOut_payload_0_3972 = (_zz_dataOut_payload_0_3971 ? _zz_dataOut_payload_0_2929 : _zz_dataOut_payload_0_2942);
  assign _zz_dataOut_payload_0_3973 = (_zz_dataOut_payload_0_3971 ? _zz_dataOut_payload_0_2942 : _zz_dataOut_payload_0_2929);
  assign _zz_dataOut_payload_0_3974 = (_zz_dataOut_payload_0_2930 < _zz_dataOut_payload_0_2941);
  assign _zz_dataOut_payload_0_3975 = (_zz_dataOut_payload_0_3974 ? _zz_dataOut_payload_0_2930 : _zz_dataOut_payload_0_2941);
  assign _zz_dataOut_payload_0_3976 = (_zz_dataOut_payload_0_3974 ? _zz_dataOut_payload_0_2941 : _zz_dataOut_payload_0_2930);
  assign _zz_dataOut_payload_0_3977 = (_zz_dataOut_payload_0_2931 < _zz_dataOut_payload_0_2940);
  assign _zz_dataOut_payload_0_3978 = (_zz_dataOut_payload_0_3977 ? _zz_dataOut_payload_0_2931 : _zz_dataOut_payload_0_2940);
  assign _zz_dataOut_payload_0_3979 = (_zz_dataOut_payload_0_3977 ? _zz_dataOut_payload_0_2940 : _zz_dataOut_payload_0_2931);
  assign _zz_dataOut_payload_0_3980 = (_zz_dataOut_payload_0_2932 < _zz_dataOut_payload_0_2939);
  assign _zz_dataOut_payload_0_3981 = (_zz_dataOut_payload_0_3980 ? _zz_dataOut_payload_0_2932 : _zz_dataOut_payload_0_2939);
  assign _zz_dataOut_payload_0_3982 = (_zz_dataOut_payload_0_3980 ? _zz_dataOut_payload_0_2939 : _zz_dataOut_payload_0_2932);
  assign _zz_dataOut_payload_0_3983 = (_zz_dataOut_payload_0_2933 < _zz_dataOut_payload_0_2938);
  assign _zz_dataOut_payload_0_3984 = (_zz_dataOut_payload_0_3983 ? _zz_dataOut_payload_0_2933 : _zz_dataOut_payload_0_2938);
  assign _zz_dataOut_payload_0_3985 = (_zz_dataOut_payload_0_3983 ? _zz_dataOut_payload_0_2938 : _zz_dataOut_payload_0_2933);
  assign _zz_dataOut_payload_0_3986 = (_zz_dataOut_payload_0_2934 < _zz_dataOut_payload_0_2937);
  assign _zz_dataOut_payload_0_3987 = (_zz_dataOut_payload_0_3986 ? _zz_dataOut_payload_0_2934 : _zz_dataOut_payload_0_2937);
  assign _zz_dataOut_payload_0_3988 = (_zz_dataOut_payload_0_3986 ? _zz_dataOut_payload_0_2937 : _zz_dataOut_payload_0_2934);
  assign _zz_dataOut_payload_0_3989 = (_zz_dataOut_payload_0_2935 < _zz_dataOut_payload_0_2936);
  assign _zz_dataOut_payload_0_3990 = (_zz_dataOut_payload_0_3989 ? _zz_dataOut_payload_0_2935 : _zz_dataOut_payload_0_2936);
  assign _zz_dataOut_payload_0_3991 = (_zz_dataOut_payload_0_3989 ? _zz_dataOut_payload_0_2936 : _zz_dataOut_payload_0_2935);
  assign _zz_dataOut_payload_0_3992 = (_zz_dataOut_payload_0_3969 < _zz_dataOut_payload_0_3981);
  assign _zz_dataOut_payload_0_3993 = (_zz_dataOut_payload_0_3992 ? _zz_dataOut_payload_0_3969 : _zz_dataOut_payload_0_3981);
  assign _zz_dataOut_payload_0_3994 = (_zz_dataOut_payload_0_3992 ? _zz_dataOut_payload_0_3981 : _zz_dataOut_payload_0_3969);
  assign _zz_dataOut_payload_0_3995 = (_zz_dataOut_payload_0_3972 < _zz_dataOut_payload_0_3984);
  assign _zz_dataOut_payload_0_3996 = (_zz_dataOut_payload_0_3995 ? _zz_dataOut_payload_0_3972 : _zz_dataOut_payload_0_3984);
  assign _zz_dataOut_payload_0_3997 = (_zz_dataOut_payload_0_3995 ? _zz_dataOut_payload_0_3984 : _zz_dataOut_payload_0_3972);
  assign _zz_dataOut_payload_0_3998 = (_zz_dataOut_payload_0_3975 < _zz_dataOut_payload_0_3987);
  assign _zz_dataOut_payload_0_3999 = (_zz_dataOut_payload_0_3998 ? _zz_dataOut_payload_0_3975 : _zz_dataOut_payload_0_3987);
  assign _zz_dataOut_payload_0_4000 = (_zz_dataOut_payload_0_3998 ? _zz_dataOut_payload_0_3987 : _zz_dataOut_payload_0_3975);
  assign _zz_dataOut_payload_0_4001 = (_zz_dataOut_payload_0_3978 < _zz_dataOut_payload_0_3990);
  assign _zz_dataOut_payload_0_4002 = (_zz_dataOut_payload_0_4001 ? _zz_dataOut_payload_0_3978 : _zz_dataOut_payload_0_3990);
  assign _zz_dataOut_payload_0_4003 = (_zz_dataOut_payload_0_4001 ? _zz_dataOut_payload_0_3990 : _zz_dataOut_payload_0_3978);
  assign _zz_dataOut_payload_0_4004 = (_zz_dataOut_payload_0_3993 < _zz_dataOut_payload_0_3999);
  assign _zz_dataOut_payload_0_4005 = (_zz_dataOut_payload_0_4004 ? _zz_dataOut_payload_0_3993 : _zz_dataOut_payload_0_3999);
  assign _zz_dataOut_payload_0_4006 = (_zz_dataOut_payload_0_4004 ? _zz_dataOut_payload_0_3999 : _zz_dataOut_payload_0_3993);
  assign _zz_dataOut_payload_0_4007 = (_zz_dataOut_payload_0_3996 < _zz_dataOut_payload_0_4002);
  assign _zz_dataOut_payload_0_4008 = (_zz_dataOut_payload_0_4007 ? _zz_dataOut_payload_0_3996 : _zz_dataOut_payload_0_4002);
  assign _zz_dataOut_payload_0_4009 = (_zz_dataOut_payload_0_4007 ? _zz_dataOut_payload_0_4002 : _zz_dataOut_payload_0_3996);
  assign _zz_dataOut_payload_0_4010 = (_zz_dataOut_payload_0_4005 < _zz_dataOut_payload_0_4008);
  assign _zz_dataOut_payload_0_4011 = (_zz_dataOut_payload_0_4006 < _zz_dataOut_payload_0_4009);
  assign _zz_dataOut_payload_0_4016 = (_zz_dataOut_payload_0_3994 < _zz_dataOut_payload_0_4000);
  assign _zz_dataOut_payload_0_4017 = (_zz_dataOut_payload_0_4016 ? _zz_dataOut_payload_0_3994 : _zz_dataOut_payload_0_4000);
  assign _zz_dataOut_payload_0_4018 = (_zz_dataOut_payload_0_4016 ? _zz_dataOut_payload_0_4000 : _zz_dataOut_payload_0_3994);
  assign _zz_dataOut_payload_0_4019 = (_zz_dataOut_payload_0_3997 < _zz_dataOut_payload_0_4003);
  assign _zz_dataOut_payload_0_4020 = (_zz_dataOut_payload_0_4019 ? _zz_dataOut_payload_0_3997 : _zz_dataOut_payload_0_4003);
  assign _zz_dataOut_payload_0_4021 = (_zz_dataOut_payload_0_4019 ? _zz_dataOut_payload_0_4003 : _zz_dataOut_payload_0_3997);
  assign _zz_dataOut_payload_0_4022 = (_zz_dataOut_payload_0_4017 < _zz_dataOut_payload_0_4020);
  assign _zz_dataOut_payload_0_4023 = (_zz_dataOut_payload_0_4018 < _zz_dataOut_payload_0_4021);
  assign _zz_dataOut_payload_0_4036 = (_zz_dataOut_payload_0_3991 < _zz_dataOut_payload_0_3979);
  assign _zz_dataOut_payload_0_4037 = (_zz_dataOut_payload_0_4036 ? _zz_dataOut_payload_0_3991 : _zz_dataOut_payload_0_3979);
  assign _zz_dataOut_payload_0_4038 = (_zz_dataOut_payload_0_4036 ? _zz_dataOut_payload_0_3979 : _zz_dataOut_payload_0_3991);
  assign _zz_dataOut_payload_0_4039 = (_zz_dataOut_payload_0_3988 < _zz_dataOut_payload_0_3976);
  assign _zz_dataOut_payload_0_4040 = (_zz_dataOut_payload_0_4039 ? _zz_dataOut_payload_0_3988 : _zz_dataOut_payload_0_3976);
  assign _zz_dataOut_payload_0_4041 = (_zz_dataOut_payload_0_4039 ? _zz_dataOut_payload_0_3976 : _zz_dataOut_payload_0_3988);
  assign _zz_dataOut_payload_0_4042 = (_zz_dataOut_payload_0_3985 < _zz_dataOut_payload_0_3973);
  assign _zz_dataOut_payload_0_4043 = (_zz_dataOut_payload_0_4042 ? _zz_dataOut_payload_0_3985 : _zz_dataOut_payload_0_3973);
  assign _zz_dataOut_payload_0_4044 = (_zz_dataOut_payload_0_4042 ? _zz_dataOut_payload_0_3973 : _zz_dataOut_payload_0_3985);
  assign _zz_dataOut_payload_0_4045 = (_zz_dataOut_payload_0_3982 < _zz_dataOut_payload_0_3970);
  assign _zz_dataOut_payload_0_4046 = (_zz_dataOut_payload_0_4045 ? _zz_dataOut_payload_0_3982 : _zz_dataOut_payload_0_3970);
  assign _zz_dataOut_payload_0_4047 = (_zz_dataOut_payload_0_4045 ? _zz_dataOut_payload_0_3970 : _zz_dataOut_payload_0_3982);
  assign _zz_dataOut_payload_0_4048 = (_zz_dataOut_payload_0_4037 < _zz_dataOut_payload_0_4043);
  assign _zz_dataOut_payload_0_4049 = (_zz_dataOut_payload_0_4048 ? _zz_dataOut_payload_0_4037 : _zz_dataOut_payload_0_4043);
  assign _zz_dataOut_payload_0_4050 = (_zz_dataOut_payload_0_4048 ? _zz_dataOut_payload_0_4043 : _zz_dataOut_payload_0_4037);
  assign _zz_dataOut_payload_0_4051 = (_zz_dataOut_payload_0_4040 < _zz_dataOut_payload_0_4046);
  assign _zz_dataOut_payload_0_4052 = (_zz_dataOut_payload_0_4051 ? _zz_dataOut_payload_0_4040 : _zz_dataOut_payload_0_4046);
  assign _zz_dataOut_payload_0_4053 = (_zz_dataOut_payload_0_4051 ? _zz_dataOut_payload_0_4046 : _zz_dataOut_payload_0_4040);
  assign _zz_dataOut_payload_0_4054 = (_zz_dataOut_payload_0_4049 < _zz_dataOut_payload_0_4052);
  assign _zz_dataOut_payload_0_4055 = (_zz_dataOut_payload_0_4050 < _zz_dataOut_payload_0_4053);
  assign _zz_dataOut_payload_0_4060 = (_zz_dataOut_payload_0_4038 < _zz_dataOut_payload_0_4044);
  assign _zz_dataOut_payload_0_4061 = (_zz_dataOut_payload_0_4060 ? _zz_dataOut_payload_0_4038 : _zz_dataOut_payload_0_4044);
  assign _zz_dataOut_payload_0_4062 = (_zz_dataOut_payload_0_4060 ? _zz_dataOut_payload_0_4044 : _zz_dataOut_payload_0_4038);
  assign _zz_dataOut_payload_0_4063 = (_zz_dataOut_payload_0_4041 < _zz_dataOut_payload_0_4047);
  assign _zz_dataOut_payload_0_4064 = (_zz_dataOut_payload_0_4063 ? _zz_dataOut_payload_0_4041 : _zz_dataOut_payload_0_4047);
  assign _zz_dataOut_payload_0_4065 = (_zz_dataOut_payload_0_4063 ? _zz_dataOut_payload_0_4047 : _zz_dataOut_payload_0_4041);
  assign _zz_dataOut_payload_0_4066 = (_zz_dataOut_payload_0_4061 < _zz_dataOut_payload_0_4064);
  assign _zz_dataOut_payload_0_4067 = (_zz_dataOut_payload_0_4062 < _zz_dataOut_payload_0_4065);
  assign _zz_dataOut_payload_0_4096 = (_zz_dataOut_payload_0_2944 < _zz_dataOut_payload_0_2959);
  assign _zz_dataOut_payload_0_4097 = (_zz_dataOut_payload_0_4096 ? _zz_dataOut_payload_0_2944 : _zz_dataOut_payload_0_2959);
  assign _zz_dataOut_payload_0_4098 = (_zz_dataOut_payload_0_4096 ? _zz_dataOut_payload_0_2959 : _zz_dataOut_payload_0_2944);
  assign _zz_dataOut_payload_0_4099 = (_zz_dataOut_payload_0_2945 < _zz_dataOut_payload_0_2958);
  assign _zz_dataOut_payload_0_4100 = (_zz_dataOut_payload_0_4099 ? _zz_dataOut_payload_0_2945 : _zz_dataOut_payload_0_2958);
  assign _zz_dataOut_payload_0_4101 = (_zz_dataOut_payload_0_4099 ? _zz_dataOut_payload_0_2958 : _zz_dataOut_payload_0_2945);
  assign _zz_dataOut_payload_0_4102 = (_zz_dataOut_payload_0_2946 < _zz_dataOut_payload_0_2957);
  assign _zz_dataOut_payload_0_4103 = (_zz_dataOut_payload_0_4102 ? _zz_dataOut_payload_0_2946 : _zz_dataOut_payload_0_2957);
  assign _zz_dataOut_payload_0_4104 = (_zz_dataOut_payload_0_4102 ? _zz_dataOut_payload_0_2957 : _zz_dataOut_payload_0_2946);
  assign _zz_dataOut_payload_0_4105 = (_zz_dataOut_payload_0_2947 < _zz_dataOut_payload_0_2956);
  assign _zz_dataOut_payload_0_4106 = (_zz_dataOut_payload_0_4105 ? _zz_dataOut_payload_0_2947 : _zz_dataOut_payload_0_2956);
  assign _zz_dataOut_payload_0_4107 = (_zz_dataOut_payload_0_4105 ? _zz_dataOut_payload_0_2956 : _zz_dataOut_payload_0_2947);
  assign _zz_dataOut_payload_0_4108 = (_zz_dataOut_payload_0_2948 < _zz_dataOut_payload_0_2955);
  assign _zz_dataOut_payload_0_4109 = (_zz_dataOut_payload_0_4108 ? _zz_dataOut_payload_0_2948 : _zz_dataOut_payload_0_2955);
  assign _zz_dataOut_payload_0_4110 = (_zz_dataOut_payload_0_4108 ? _zz_dataOut_payload_0_2955 : _zz_dataOut_payload_0_2948);
  assign _zz_dataOut_payload_0_4111 = (_zz_dataOut_payload_0_2949 < _zz_dataOut_payload_0_2954);
  assign _zz_dataOut_payload_0_4112 = (_zz_dataOut_payload_0_4111 ? _zz_dataOut_payload_0_2949 : _zz_dataOut_payload_0_2954);
  assign _zz_dataOut_payload_0_4113 = (_zz_dataOut_payload_0_4111 ? _zz_dataOut_payload_0_2954 : _zz_dataOut_payload_0_2949);
  assign _zz_dataOut_payload_0_4114 = (_zz_dataOut_payload_0_2950 < _zz_dataOut_payload_0_2953);
  assign _zz_dataOut_payload_0_4115 = (_zz_dataOut_payload_0_4114 ? _zz_dataOut_payload_0_2950 : _zz_dataOut_payload_0_2953);
  assign _zz_dataOut_payload_0_4116 = (_zz_dataOut_payload_0_4114 ? _zz_dataOut_payload_0_2953 : _zz_dataOut_payload_0_2950);
  assign _zz_dataOut_payload_0_4117 = (_zz_dataOut_payload_0_2951 < _zz_dataOut_payload_0_2952);
  assign _zz_dataOut_payload_0_4118 = (_zz_dataOut_payload_0_4117 ? _zz_dataOut_payload_0_2951 : _zz_dataOut_payload_0_2952);
  assign _zz_dataOut_payload_0_4119 = (_zz_dataOut_payload_0_4117 ? _zz_dataOut_payload_0_2952 : _zz_dataOut_payload_0_2951);
  assign _zz_dataOut_payload_0_4120 = (_zz_dataOut_payload_0_4097 < _zz_dataOut_payload_0_4109);
  assign _zz_dataOut_payload_0_4121 = (_zz_dataOut_payload_0_4120 ? _zz_dataOut_payload_0_4097 : _zz_dataOut_payload_0_4109);
  assign _zz_dataOut_payload_0_4122 = (_zz_dataOut_payload_0_4120 ? _zz_dataOut_payload_0_4109 : _zz_dataOut_payload_0_4097);
  assign _zz_dataOut_payload_0_4123 = (_zz_dataOut_payload_0_4100 < _zz_dataOut_payload_0_4112);
  assign _zz_dataOut_payload_0_4124 = (_zz_dataOut_payload_0_4123 ? _zz_dataOut_payload_0_4100 : _zz_dataOut_payload_0_4112);
  assign _zz_dataOut_payload_0_4125 = (_zz_dataOut_payload_0_4123 ? _zz_dataOut_payload_0_4112 : _zz_dataOut_payload_0_4100);
  assign _zz_dataOut_payload_0_4126 = (_zz_dataOut_payload_0_4103 < _zz_dataOut_payload_0_4115);
  assign _zz_dataOut_payload_0_4127 = (_zz_dataOut_payload_0_4126 ? _zz_dataOut_payload_0_4103 : _zz_dataOut_payload_0_4115);
  assign _zz_dataOut_payload_0_4128 = (_zz_dataOut_payload_0_4126 ? _zz_dataOut_payload_0_4115 : _zz_dataOut_payload_0_4103);
  assign _zz_dataOut_payload_0_4129 = (_zz_dataOut_payload_0_4106 < _zz_dataOut_payload_0_4118);
  assign _zz_dataOut_payload_0_4130 = (_zz_dataOut_payload_0_4129 ? _zz_dataOut_payload_0_4106 : _zz_dataOut_payload_0_4118);
  assign _zz_dataOut_payload_0_4131 = (_zz_dataOut_payload_0_4129 ? _zz_dataOut_payload_0_4118 : _zz_dataOut_payload_0_4106);
  assign _zz_dataOut_payload_0_4132 = (_zz_dataOut_payload_0_4121 < _zz_dataOut_payload_0_4127);
  assign _zz_dataOut_payload_0_4133 = (_zz_dataOut_payload_0_4132 ? _zz_dataOut_payload_0_4121 : _zz_dataOut_payload_0_4127);
  assign _zz_dataOut_payload_0_4134 = (_zz_dataOut_payload_0_4132 ? _zz_dataOut_payload_0_4127 : _zz_dataOut_payload_0_4121);
  assign _zz_dataOut_payload_0_4135 = (_zz_dataOut_payload_0_4124 < _zz_dataOut_payload_0_4130);
  assign _zz_dataOut_payload_0_4136 = (_zz_dataOut_payload_0_4135 ? _zz_dataOut_payload_0_4124 : _zz_dataOut_payload_0_4130);
  assign _zz_dataOut_payload_0_4137 = (_zz_dataOut_payload_0_4135 ? _zz_dataOut_payload_0_4130 : _zz_dataOut_payload_0_4124);
  assign _zz_dataOut_payload_0_4138 = (_zz_dataOut_payload_0_4133 < _zz_dataOut_payload_0_4136);
  assign _zz_dataOut_payload_0_4139 = (_zz_dataOut_payload_0_4134 < _zz_dataOut_payload_0_4137);
  assign _zz_dataOut_payload_0_4144 = (_zz_dataOut_payload_0_4122 < _zz_dataOut_payload_0_4128);
  assign _zz_dataOut_payload_0_4145 = (_zz_dataOut_payload_0_4144 ? _zz_dataOut_payload_0_4122 : _zz_dataOut_payload_0_4128);
  assign _zz_dataOut_payload_0_4146 = (_zz_dataOut_payload_0_4144 ? _zz_dataOut_payload_0_4128 : _zz_dataOut_payload_0_4122);
  assign _zz_dataOut_payload_0_4147 = (_zz_dataOut_payload_0_4125 < _zz_dataOut_payload_0_4131);
  assign _zz_dataOut_payload_0_4148 = (_zz_dataOut_payload_0_4147 ? _zz_dataOut_payload_0_4125 : _zz_dataOut_payload_0_4131);
  assign _zz_dataOut_payload_0_4149 = (_zz_dataOut_payload_0_4147 ? _zz_dataOut_payload_0_4131 : _zz_dataOut_payload_0_4125);
  assign _zz_dataOut_payload_0_4150 = (_zz_dataOut_payload_0_4145 < _zz_dataOut_payload_0_4148);
  assign _zz_dataOut_payload_0_4151 = (_zz_dataOut_payload_0_4146 < _zz_dataOut_payload_0_4149);
  assign _zz_dataOut_payload_0_4164 = (_zz_dataOut_payload_0_4119 < _zz_dataOut_payload_0_4107);
  assign _zz_dataOut_payload_0_4165 = (_zz_dataOut_payload_0_4164 ? _zz_dataOut_payload_0_4119 : _zz_dataOut_payload_0_4107);
  assign _zz_dataOut_payload_0_4166 = (_zz_dataOut_payload_0_4164 ? _zz_dataOut_payload_0_4107 : _zz_dataOut_payload_0_4119);
  assign _zz_dataOut_payload_0_4167 = (_zz_dataOut_payload_0_4116 < _zz_dataOut_payload_0_4104);
  assign _zz_dataOut_payload_0_4168 = (_zz_dataOut_payload_0_4167 ? _zz_dataOut_payload_0_4116 : _zz_dataOut_payload_0_4104);
  assign _zz_dataOut_payload_0_4169 = (_zz_dataOut_payload_0_4167 ? _zz_dataOut_payload_0_4104 : _zz_dataOut_payload_0_4116);
  assign _zz_dataOut_payload_0_4170 = (_zz_dataOut_payload_0_4113 < _zz_dataOut_payload_0_4101);
  assign _zz_dataOut_payload_0_4171 = (_zz_dataOut_payload_0_4170 ? _zz_dataOut_payload_0_4113 : _zz_dataOut_payload_0_4101);
  assign _zz_dataOut_payload_0_4172 = (_zz_dataOut_payload_0_4170 ? _zz_dataOut_payload_0_4101 : _zz_dataOut_payload_0_4113);
  assign _zz_dataOut_payload_0_4173 = (_zz_dataOut_payload_0_4110 < _zz_dataOut_payload_0_4098);
  assign _zz_dataOut_payload_0_4174 = (_zz_dataOut_payload_0_4173 ? _zz_dataOut_payload_0_4110 : _zz_dataOut_payload_0_4098);
  assign _zz_dataOut_payload_0_4175 = (_zz_dataOut_payload_0_4173 ? _zz_dataOut_payload_0_4098 : _zz_dataOut_payload_0_4110);
  assign _zz_dataOut_payload_0_4176 = (_zz_dataOut_payload_0_4165 < _zz_dataOut_payload_0_4171);
  assign _zz_dataOut_payload_0_4177 = (_zz_dataOut_payload_0_4176 ? _zz_dataOut_payload_0_4165 : _zz_dataOut_payload_0_4171);
  assign _zz_dataOut_payload_0_4178 = (_zz_dataOut_payload_0_4176 ? _zz_dataOut_payload_0_4171 : _zz_dataOut_payload_0_4165);
  assign _zz_dataOut_payload_0_4179 = (_zz_dataOut_payload_0_4168 < _zz_dataOut_payload_0_4174);
  assign _zz_dataOut_payload_0_4180 = (_zz_dataOut_payload_0_4179 ? _zz_dataOut_payload_0_4168 : _zz_dataOut_payload_0_4174);
  assign _zz_dataOut_payload_0_4181 = (_zz_dataOut_payload_0_4179 ? _zz_dataOut_payload_0_4174 : _zz_dataOut_payload_0_4168);
  assign _zz_dataOut_payload_0_4182 = (_zz_dataOut_payload_0_4177 < _zz_dataOut_payload_0_4180);
  assign _zz_dataOut_payload_0_4183 = (_zz_dataOut_payload_0_4178 < _zz_dataOut_payload_0_4181);
  assign _zz_dataOut_payload_0_4188 = (_zz_dataOut_payload_0_4166 < _zz_dataOut_payload_0_4172);
  assign _zz_dataOut_payload_0_4189 = (_zz_dataOut_payload_0_4188 ? _zz_dataOut_payload_0_4166 : _zz_dataOut_payload_0_4172);
  assign _zz_dataOut_payload_0_4190 = (_zz_dataOut_payload_0_4188 ? _zz_dataOut_payload_0_4172 : _zz_dataOut_payload_0_4166);
  assign _zz_dataOut_payload_0_4191 = (_zz_dataOut_payload_0_4169 < _zz_dataOut_payload_0_4175);
  assign _zz_dataOut_payload_0_4192 = (_zz_dataOut_payload_0_4191 ? _zz_dataOut_payload_0_4169 : _zz_dataOut_payload_0_4175);
  assign _zz_dataOut_payload_0_4193 = (_zz_dataOut_payload_0_4191 ? _zz_dataOut_payload_0_4175 : _zz_dataOut_payload_0_4169);
  assign _zz_dataOut_payload_0_4194 = (_zz_dataOut_payload_0_4189 < _zz_dataOut_payload_0_4192);
  assign _zz_dataOut_payload_0_4195 = (_zz_dataOut_payload_0_4190 < _zz_dataOut_payload_0_4193);
  assign _zz_dataOut_payload_0_4224 = (_zz_dataOut_payload_0_2960 < _zz_dataOut_payload_0_2975);
  assign _zz_dataOut_payload_0_4225 = (_zz_dataOut_payload_0_4224 ? _zz_dataOut_payload_0_2960 : _zz_dataOut_payload_0_2975);
  assign _zz_dataOut_payload_0_4226 = (_zz_dataOut_payload_0_4224 ? _zz_dataOut_payload_0_2975 : _zz_dataOut_payload_0_2960);
  assign _zz_dataOut_payload_0_4227 = (_zz_dataOut_payload_0_2961 < _zz_dataOut_payload_0_2974);
  assign _zz_dataOut_payload_0_4228 = (_zz_dataOut_payload_0_4227 ? _zz_dataOut_payload_0_2961 : _zz_dataOut_payload_0_2974);
  assign _zz_dataOut_payload_0_4229 = (_zz_dataOut_payload_0_4227 ? _zz_dataOut_payload_0_2974 : _zz_dataOut_payload_0_2961);
  assign _zz_dataOut_payload_0_4230 = (_zz_dataOut_payload_0_2962 < _zz_dataOut_payload_0_2973);
  assign _zz_dataOut_payload_0_4231 = (_zz_dataOut_payload_0_4230 ? _zz_dataOut_payload_0_2962 : _zz_dataOut_payload_0_2973);
  assign _zz_dataOut_payload_0_4232 = (_zz_dataOut_payload_0_4230 ? _zz_dataOut_payload_0_2973 : _zz_dataOut_payload_0_2962);
  assign _zz_dataOut_payload_0_4233 = (_zz_dataOut_payload_0_2963 < _zz_dataOut_payload_0_2972);
  assign _zz_dataOut_payload_0_4234 = (_zz_dataOut_payload_0_4233 ? _zz_dataOut_payload_0_2963 : _zz_dataOut_payload_0_2972);
  assign _zz_dataOut_payload_0_4235 = (_zz_dataOut_payload_0_4233 ? _zz_dataOut_payload_0_2972 : _zz_dataOut_payload_0_2963);
  assign _zz_dataOut_payload_0_4236 = (_zz_dataOut_payload_0_2964 < _zz_dataOut_payload_0_2971);
  assign _zz_dataOut_payload_0_4237 = (_zz_dataOut_payload_0_4236 ? _zz_dataOut_payload_0_2964 : _zz_dataOut_payload_0_2971);
  assign _zz_dataOut_payload_0_4238 = (_zz_dataOut_payload_0_4236 ? _zz_dataOut_payload_0_2971 : _zz_dataOut_payload_0_2964);
  assign _zz_dataOut_payload_0_4239 = (_zz_dataOut_payload_0_2965 < _zz_dataOut_payload_0_2970);
  assign _zz_dataOut_payload_0_4240 = (_zz_dataOut_payload_0_4239 ? _zz_dataOut_payload_0_2965 : _zz_dataOut_payload_0_2970);
  assign _zz_dataOut_payload_0_4241 = (_zz_dataOut_payload_0_4239 ? _zz_dataOut_payload_0_2970 : _zz_dataOut_payload_0_2965);
  assign _zz_dataOut_payload_0_4242 = (_zz_dataOut_payload_0_2966 < _zz_dataOut_payload_0_2969);
  assign _zz_dataOut_payload_0_4243 = (_zz_dataOut_payload_0_4242 ? _zz_dataOut_payload_0_2966 : _zz_dataOut_payload_0_2969);
  assign _zz_dataOut_payload_0_4244 = (_zz_dataOut_payload_0_4242 ? _zz_dataOut_payload_0_2969 : _zz_dataOut_payload_0_2966);
  assign _zz_dataOut_payload_0_4245 = (_zz_dataOut_payload_0_2967 < _zz_dataOut_payload_0_2968);
  assign _zz_dataOut_payload_0_4246 = (_zz_dataOut_payload_0_4245 ? _zz_dataOut_payload_0_2967 : _zz_dataOut_payload_0_2968);
  assign _zz_dataOut_payload_0_4247 = (_zz_dataOut_payload_0_4245 ? _zz_dataOut_payload_0_2968 : _zz_dataOut_payload_0_2967);
  assign _zz_dataOut_payload_0_4248 = (_zz_dataOut_payload_0_4225 < _zz_dataOut_payload_0_4237);
  assign _zz_dataOut_payload_0_4249 = (_zz_dataOut_payload_0_4248 ? _zz_dataOut_payload_0_4225 : _zz_dataOut_payload_0_4237);
  assign _zz_dataOut_payload_0_4250 = (_zz_dataOut_payload_0_4248 ? _zz_dataOut_payload_0_4237 : _zz_dataOut_payload_0_4225);
  assign _zz_dataOut_payload_0_4251 = (_zz_dataOut_payload_0_4228 < _zz_dataOut_payload_0_4240);
  assign _zz_dataOut_payload_0_4252 = (_zz_dataOut_payload_0_4251 ? _zz_dataOut_payload_0_4228 : _zz_dataOut_payload_0_4240);
  assign _zz_dataOut_payload_0_4253 = (_zz_dataOut_payload_0_4251 ? _zz_dataOut_payload_0_4240 : _zz_dataOut_payload_0_4228);
  assign _zz_dataOut_payload_0_4254 = (_zz_dataOut_payload_0_4231 < _zz_dataOut_payload_0_4243);
  assign _zz_dataOut_payload_0_4255 = (_zz_dataOut_payload_0_4254 ? _zz_dataOut_payload_0_4231 : _zz_dataOut_payload_0_4243);
  assign _zz_dataOut_payload_0_4256 = (_zz_dataOut_payload_0_4254 ? _zz_dataOut_payload_0_4243 : _zz_dataOut_payload_0_4231);
  assign _zz_dataOut_payload_0_4257 = (_zz_dataOut_payload_0_4234 < _zz_dataOut_payload_0_4246);
  assign _zz_dataOut_payload_0_4258 = (_zz_dataOut_payload_0_4257 ? _zz_dataOut_payload_0_4234 : _zz_dataOut_payload_0_4246);
  assign _zz_dataOut_payload_0_4259 = (_zz_dataOut_payload_0_4257 ? _zz_dataOut_payload_0_4246 : _zz_dataOut_payload_0_4234);
  assign _zz_dataOut_payload_0_4260 = (_zz_dataOut_payload_0_4249 < _zz_dataOut_payload_0_4255);
  assign _zz_dataOut_payload_0_4261 = (_zz_dataOut_payload_0_4260 ? _zz_dataOut_payload_0_4249 : _zz_dataOut_payload_0_4255);
  assign _zz_dataOut_payload_0_4262 = (_zz_dataOut_payload_0_4260 ? _zz_dataOut_payload_0_4255 : _zz_dataOut_payload_0_4249);
  assign _zz_dataOut_payload_0_4263 = (_zz_dataOut_payload_0_4252 < _zz_dataOut_payload_0_4258);
  assign _zz_dataOut_payload_0_4264 = (_zz_dataOut_payload_0_4263 ? _zz_dataOut_payload_0_4252 : _zz_dataOut_payload_0_4258);
  assign _zz_dataOut_payload_0_4265 = (_zz_dataOut_payload_0_4263 ? _zz_dataOut_payload_0_4258 : _zz_dataOut_payload_0_4252);
  assign _zz_dataOut_payload_0_4266 = (_zz_dataOut_payload_0_4261 < _zz_dataOut_payload_0_4264);
  assign _zz_dataOut_payload_0_4267 = (_zz_dataOut_payload_0_4262 < _zz_dataOut_payload_0_4265);
  assign _zz_dataOut_payload_0_4272 = (_zz_dataOut_payload_0_4250 < _zz_dataOut_payload_0_4256);
  assign _zz_dataOut_payload_0_4273 = (_zz_dataOut_payload_0_4272 ? _zz_dataOut_payload_0_4250 : _zz_dataOut_payload_0_4256);
  assign _zz_dataOut_payload_0_4274 = (_zz_dataOut_payload_0_4272 ? _zz_dataOut_payload_0_4256 : _zz_dataOut_payload_0_4250);
  assign _zz_dataOut_payload_0_4275 = (_zz_dataOut_payload_0_4253 < _zz_dataOut_payload_0_4259);
  assign _zz_dataOut_payload_0_4276 = (_zz_dataOut_payload_0_4275 ? _zz_dataOut_payload_0_4253 : _zz_dataOut_payload_0_4259);
  assign _zz_dataOut_payload_0_4277 = (_zz_dataOut_payload_0_4275 ? _zz_dataOut_payload_0_4259 : _zz_dataOut_payload_0_4253);
  assign _zz_dataOut_payload_0_4278 = (_zz_dataOut_payload_0_4273 < _zz_dataOut_payload_0_4276);
  assign _zz_dataOut_payload_0_4279 = (_zz_dataOut_payload_0_4274 < _zz_dataOut_payload_0_4277);
  assign _zz_dataOut_payload_0_4292 = (_zz_dataOut_payload_0_4247 < _zz_dataOut_payload_0_4235);
  assign _zz_dataOut_payload_0_4293 = (_zz_dataOut_payload_0_4292 ? _zz_dataOut_payload_0_4247 : _zz_dataOut_payload_0_4235);
  assign _zz_dataOut_payload_0_4294 = (_zz_dataOut_payload_0_4292 ? _zz_dataOut_payload_0_4235 : _zz_dataOut_payload_0_4247);
  assign _zz_dataOut_payload_0_4295 = (_zz_dataOut_payload_0_4244 < _zz_dataOut_payload_0_4232);
  assign _zz_dataOut_payload_0_4296 = (_zz_dataOut_payload_0_4295 ? _zz_dataOut_payload_0_4244 : _zz_dataOut_payload_0_4232);
  assign _zz_dataOut_payload_0_4297 = (_zz_dataOut_payload_0_4295 ? _zz_dataOut_payload_0_4232 : _zz_dataOut_payload_0_4244);
  assign _zz_dataOut_payload_0_4298 = (_zz_dataOut_payload_0_4241 < _zz_dataOut_payload_0_4229);
  assign _zz_dataOut_payload_0_4299 = (_zz_dataOut_payload_0_4298 ? _zz_dataOut_payload_0_4241 : _zz_dataOut_payload_0_4229);
  assign _zz_dataOut_payload_0_4300 = (_zz_dataOut_payload_0_4298 ? _zz_dataOut_payload_0_4229 : _zz_dataOut_payload_0_4241);
  assign _zz_dataOut_payload_0_4301 = (_zz_dataOut_payload_0_4238 < _zz_dataOut_payload_0_4226);
  assign _zz_dataOut_payload_0_4302 = (_zz_dataOut_payload_0_4301 ? _zz_dataOut_payload_0_4238 : _zz_dataOut_payload_0_4226);
  assign _zz_dataOut_payload_0_4303 = (_zz_dataOut_payload_0_4301 ? _zz_dataOut_payload_0_4226 : _zz_dataOut_payload_0_4238);
  assign _zz_dataOut_payload_0_4304 = (_zz_dataOut_payload_0_4293 < _zz_dataOut_payload_0_4299);
  assign _zz_dataOut_payload_0_4305 = (_zz_dataOut_payload_0_4304 ? _zz_dataOut_payload_0_4293 : _zz_dataOut_payload_0_4299);
  assign _zz_dataOut_payload_0_4306 = (_zz_dataOut_payload_0_4304 ? _zz_dataOut_payload_0_4299 : _zz_dataOut_payload_0_4293);
  assign _zz_dataOut_payload_0_4307 = (_zz_dataOut_payload_0_4296 < _zz_dataOut_payload_0_4302);
  assign _zz_dataOut_payload_0_4308 = (_zz_dataOut_payload_0_4307 ? _zz_dataOut_payload_0_4296 : _zz_dataOut_payload_0_4302);
  assign _zz_dataOut_payload_0_4309 = (_zz_dataOut_payload_0_4307 ? _zz_dataOut_payload_0_4302 : _zz_dataOut_payload_0_4296);
  assign _zz_dataOut_payload_0_4310 = (_zz_dataOut_payload_0_4305 < _zz_dataOut_payload_0_4308);
  assign _zz_dataOut_payload_0_4311 = (_zz_dataOut_payload_0_4306 < _zz_dataOut_payload_0_4309);
  assign _zz_dataOut_payload_0_4316 = (_zz_dataOut_payload_0_4294 < _zz_dataOut_payload_0_4300);
  assign _zz_dataOut_payload_0_4317 = (_zz_dataOut_payload_0_4316 ? _zz_dataOut_payload_0_4294 : _zz_dataOut_payload_0_4300);
  assign _zz_dataOut_payload_0_4318 = (_zz_dataOut_payload_0_4316 ? _zz_dataOut_payload_0_4300 : _zz_dataOut_payload_0_4294);
  assign _zz_dataOut_payload_0_4319 = (_zz_dataOut_payload_0_4297 < _zz_dataOut_payload_0_4303);
  assign _zz_dataOut_payload_0_4320 = (_zz_dataOut_payload_0_4319 ? _zz_dataOut_payload_0_4297 : _zz_dataOut_payload_0_4303);
  assign _zz_dataOut_payload_0_4321 = (_zz_dataOut_payload_0_4319 ? _zz_dataOut_payload_0_4303 : _zz_dataOut_payload_0_4297);
  assign _zz_dataOut_payload_0_4322 = (_zz_dataOut_payload_0_4317 < _zz_dataOut_payload_0_4320);
  assign _zz_dataOut_payload_0_4323 = (_zz_dataOut_payload_0_4318 < _zz_dataOut_payload_0_4321);
  assign _zz_dataOut_payload_0_4352 = (_zz_dataOut_payload_0_2976 < _zz_dataOut_payload_0_2991);
  assign _zz_dataOut_payload_0_4353 = (_zz_dataOut_payload_0_4352 ? _zz_dataOut_payload_0_2976 : _zz_dataOut_payload_0_2991);
  assign _zz_dataOut_payload_0_4354 = (_zz_dataOut_payload_0_4352 ? _zz_dataOut_payload_0_2991 : _zz_dataOut_payload_0_2976);
  assign _zz_dataOut_payload_0_4355 = (_zz_dataOut_payload_0_2977 < _zz_dataOut_payload_0_2990);
  assign _zz_dataOut_payload_0_4356 = (_zz_dataOut_payload_0_4355 ? _zz_dataOut_payload_0_2977 : _zz_dataOut_payload_0_2990);
  assign _zz_dataOut_payload_0_4357 = (_zz_dataOut_payload_0_4355 ? _zz_dataOut_payload_0_2990 : _zz_dataOut_payload_0_2977);
  assign _zz_dataOut_payload_0_4358 = (_zz_dataOut_payload_0_2978 < _zz_dataOut_payload_0_2989);
  assign _zz_dataOut_payload_0_4359 = (_zz_dataOut_payload_0_4358 ? _zz_dataOut_payload_0_2978 : _zz_dataOut_payload_0_2989);
  assign _zz_dataOut_payload_0_4360 = (_zz_dataOut_payload_0_4358 ? _zz_dataOut_payload_0_2989 : _zz_dataOut_payload_0_2978);
  assign _zz_dataOut_payload_0_4361 = (_zz_dataOut_payload_0_2979 < _zz_dataOut_payload_0_2988);
  assign _zz_dataOut_payload_0_4362 = (_zz_dataOut_payload_0_4361 ? _zz_dataOut_payload_0_2979 : _zz_dataOut_payload_0_2988);
  assign _zz_dataOut_payload_0_4363 = (_zz_dataOut_payload_0_4361 ? _zz_dataOut_payload_0_2988 : _zz_dataOut_payload_0_2979);
  assign _zz_dataOut_payload_0_4364 = (_zz_dataOut_payload_0_2980 < _zz_dataOut_payload_0_2987);
  assign _zz_dataOut_payload_0_4365 = (_zz_dataOut_payload_0_4364 ? _zz_dataOut_payload_0_2980 : _zz_dataOut_payload_0_2987);
  assign _zz_dataOut_payload_0_4366 = (_zz_dataOut_payload_0_4364 ? _zz_dataOut_payload_0_2987 : _zz_dataOut_payload_0_2980);
  assign _zz_dataOut_payload_0_4367 = (_zz_dataOut_payload_0_2981 < _zz_dataOut_payload_0_2986);
  assign _zz_dataOut_payload_0_4368 = (_zz_dataOut_payload_0_4367 ? _zz_dataOut_payload_0_2981 : _zz_dataOut_payload_0_2986);
  assign _zz_dataOut_payload_0_4369 = (_zz_dataOut_payload_0_4367 ? _zz_dataOut_payload_0_2986 : _zz_dataOut_payload_0_2981);
  assign _zz_dataOut_payload_0_4370 = (_zz_dataOut_payload_0_2982 < _zz_dataOut_payload_0_2985);
  assign _zz_dataOut_payload_0_4371 = (_zz_dataOut_payload_0_4370 ? _zz_dataOut_payload_0_2982 : _zz_dataOut_payload_0_2985);
  assign _zz_dataOut_payload_0_4372 = (_zz_dataOut_payload_0_4370 ? _zz_dataOut_payload_0_2985 : _zz_dataOut_payload_0_2982);
  assign _zz_dataOut_payload_0_4373 = (_zz_dataOut_payload_0_2983 < _zz_dataOut_payload_0_2984);
  assign _zz_dataOut_payload_0_4374 = (_zz_dataOut_payload_0_4373 ? _zz_dataOut_payload_0_2983 : _zz_dataOut_payload_0_2984);
  assign _zz_dataOut_payload_0_4375 = (_zz_dataOut_payload_0_4373 ? _zz_dataOut_payload_0_2984 : _zz_dataOut_payload_0_2983);
  assign _zz_dataOut_payload_0_4376 = (_zz_dataOut_payload_0_4353 < _zz_dataOut_payload_0_4365);
  assign _zz_dataOut_payload_0_4377 = (_zz_dataOut_payload_0_4376 ? _zz_dataOut_payload_0_4353 : _zz_dataOut_payload_0_4365);
  assign _zz_dataOut_payload_0_4378 = (_zz_dataOut_payload_0_4376 ? _zz_dataOut_payload_0_4365 : _zz_dataOut_payload_0_4353);
  assign _zz_dataOut_payload_0_4379 = (_zz_dataOut_payload_0_4356 < _zz_dataOut_payload_0_4368);
  assign _zz_dataOut_payload_0_4380 = (_zz_dataOut_payload_0_4379 ? _zz_dataOut_payload_0_4356 : _zz_dataOut_payload_0_4368);
  assign _zz_dataOut_payload_0_4381 = (_zz_dataOut_payload_0_4379 ? _zz_dataOut_payload_0_4368 : _zz_dataOut_payload_0_4356);
  assign _zz_dataOut_payload_0_4382 = (_zz_dataOut_payload_0_4359 < _zz_dataOut_payload_0_4371);
  assign _zz_dataOut_payload_0_4383 = (_zz_dataOut_payload_0_4382 ? _zz_dataOut_payload_0_4359 : _zz_dataOut_payload_0_4371);
  assign _zz_dataOut_payload_0_4384 = (_zz_dataOut_payload_0_4382 ? _zz_dataOut_payload_0_4371 : _zz_dataOut_payload_0_4359);
  assign _zz_dataOut_payload_0_4385 = (_zz_dataOut_payload_0_4362 < _zz_dataOut_payload_0_4374);
  assign _zz_dataOut_payload_0_4386 = (_zz_dataOut_payload_0_4385 ? _zz_dataOut_payload_0_4362 : _zz_dataOut_payload_0_4374);
  assign _zz_dataOut_payload_0_4387 = (_zz_dataOut_payload_0_4385 ? _zz_dataOut_payload_0_4374 : _zz_dataOut_payload_0_4362);
  assign _zz_dataOut_payload_0_4388 = (_zz_dataOut_payload_0_4377 < _zz_dataOut_payload_0_4383);
  assign _zz_dataOut_payload_0_4389 = (_zz_dataOut_payload_0_4388 ? _zz_dataOut_payload_0_4377 : _zz_dataOut_payload_0_4383);
  assign _zz_dataOut_payload_0_4390 = (_zz_dataOut_payload_0_4388 ? _zz_dataOut_payload_0_4383 : _zz_dataOut_payload_0_4377);
  assign _zz_dataOut_payload_0_4391 = (_zz_dataOut_payload_0_4380 < _zz_dataOut_payload_0_4386);
  assign _zz_dataOut_payload_0_4392 = (_zz_dataOut_payload_0_4391 ? _zz_dataOut_payload_0_4380 : _zz_dataOut_payload_0_4386);
  assign _zz_dataOut_payload_0_4393 = (_zz_dataOut_payload_0_4391 ? _zz_dataOut_payload_0_4386 : _zz_dataOut_payload_0_4380);
  assign _zz_dataOut_payload_0_4394 = (_zz_dataOut_payload_0_4389 < _zz_dataOut_payload_0_4392);
  assign _zz_dataOut_payload_0_4395 = (_zz_dataOut_payload_0_4390 < _zz_dataOut_payload_0_4393);
  assign _zz_dataOut_payload_0_4400 = (_zz_dataOut_payload_0_4378 < _zz_dataOut_payload_0_4384);
  assign _zz_dataOut_payload_0_4401 = (_zz_dataOut_payload_0_4400 ? _zz_dataOut_payload_0_4378 : _zz_dataOut_payload_0_4384);
  assign _zz_dataOut_payload_0_4402 = (_zz_dataOut_payload_0_4400 ? _zz_dataOut_payload_0_4384 : _zz_dataOut_payload_0_4378);
  assign _zz_dataOut_payload_0_4403 = (_zz_dataOut_payload_0_4381 < _zz_dataOut_payload_0_4387);
  assign _zz_dataOut_payload_0_4404 = (_zz_dataOut_payload_0_4403 ? _zz_dataOut_payload_0_4381 : _zz_dataOut_payload_0_4387);
  assign _zz_dataOut_payload_0_4405 = (_zz_dataOut_payload_0_4403 ? _zz_dataOut_payload_0_4387 : _zz_dataOut_payload_0_4381);
  assign _zz_dataOut_payload_0_4406 = (_zz_dataOut_payload_0_4401 < _zz_dataOut_payload_0_4404);
  assign _zz_dataOut_payload_0_4407 = (_zz_dataOut_payload_0_4402 < _zz_dataOut_payload_0_4405);
  assign _zz_dataOut_payload_0_4420 = (_zz_dataOut_payload_0_4375 < _zz_dataOut_payload_0_4363);
  assign _zz_dataOut_payload_0_4421 = (_zz_dataOut_payload_0_4420 ? _zz_dataOut_payload_0_4375 : _zz_dataOut_payload_0_4363);
  assign _zz_dataOut_payload_0_4422 = (_zz_dataOut_payload_0_4420 ? _zz_dataOut_payload_0_4363 : _zz_dataOut_payload_0_4375);
  assign _zz_dataOut_payload_0_4423 = (_zz_dataOut_payload_0_4372 < _zz_dataOut_payload_0_4360);
  assign _zz_dataOut_payload_0_4424 = (_zz_dataOut_payload_0_4423 ? _zz_dataOut_payload_0_4372 : _zz_dataOut_payload_0_4360);
  assign _zz_dataOut_payload_0_4425 = (_zz_dataOut_payload_0_4423 ? _zz_dataOut_payload_0_4360 : _zz_dataOut_payload_0_4372);
  assign _zz_dataOut_payload_0_4426 = (_zz_dataOut_payload_0_4369 < _zz_dataOut_payload_0_4357);
  assign _zz_dataOut_payload_0_4427 = (_zz_dataOut_payload_0_4426 ? _zz_dataOut_payload_0_4369 : _zz_dataOut_payload_0_4357);
  assign _zz_dataOut_payload_0_4428 = (_zz_dataOut_payload_0_4426 ? _zz_dataOut_payload_0_4357 : _zz_dataOut_payload_0_4369);
  assign _zz_dataOut_payload_0_4429 = (_zz_dataOut_payload_0_4366 < _zz_dataOut_payload_0_4354);
  assign _zz_dataOut_payload_0_4430 = (_zz_dataOut_payload_0_4429 ? _zz_dataOut_payload_0_4366 : _zz_dataOut_payload_0_4354);
  assign _zz_dataOut_payload_0_4431 = (_zz_dataOut_payload_0_4429 ? _zz_dataOut_payload_0_4354 : _zz_dataOut_payload_0_4366);
  assign _zz_dataOut_payload_0_4432 = (_zz_dataOut_payload_0_4421 < _zz_dataOut_payload_0_4427);
  assign _zz_dataOut_payload_0_4433 = (_zz_dataOut_payload_0_4432 ? _zz_dataOut_payload_0_4421 : _zz_dataOut_payload_0_4427);
  assign _zz_dataOut_payload_0_4434 = (_zz_dataOut_payload_0_4432 ? _zz_dataOut_payload_0_4427 : _zz_dataOut_payload_0_4421);
  assign _zz_dataOut_payload_0_4435 = (_zz_dataOut_payload_0_4424 < _zz_dataOut_payload_0_4430);
  assign _zz_dataOut_payload_0_4436 = (_zz_dataOut_payload_0_4435 ? _zz_dataOut_payload_0_4424 : _zz_dataOut_payload_0_4430);
  assign _zz_dataOut_payload_0_4437 = (_zz_dataOut_payload_0_4435 ? _zz_dataOut_payload_0_4430 : _zz_dataOut_payload_0_4424);
  assign _zz_dataOut_payload_0_4438 = (_zz_dataOut_payload_0_4433 < _zz_dataOut_payload_0_4436);
  assign _zz_dataOut_payload_0_4439 = (_zz_dataOut_payload_0_4434 < _zz_dataOut_payload_0_4437);
  assign _zz_dataOut_payload_0_4444 = (_zz_dataOut_payload_0_4422 < _zz_dataOut_payload_0_4428);
  assign _zz_dataOut_payload_0_4445 = (_zz_dataOut_payload_0_4444 ? _zz_dataOut_payload_0_4422 : _zz_dataOut_payload_0_4428);
  assign _zz_dataOut_payload_0_4446 = (_zz_dataOut_payload_0_4444 ? _zz_dataOut_payload_0_4428 : _zz_dataOut_payload_0_4422);
  assign _zz_dataOut_payload_0_4447 = (_zz_dataOut_payload_0_4425 < _zz_dataOut_payload_0_4431);
  assign _zz_dataOut_payload_0_4448 = (_zz_dataOut_payload_0_4447 ? _zz_dataOut_payload_0_4425 : _zz_dataOut_payload_0_4431);
  assign _zz_dataOut_payload_0_4449 = (_zz_dataOut_payload_0_4447 ? _zz_dataOut_payload_0_4431 : _zz_dataOut_payload_0_4425);
  assign _zz_dataOut_payload_0_4450 = (_zz_dataOut_payload_0_4445 < _zz_dataOut_payload_0_4448);
  assign _zz_dataOut_payload_0_4451 = (_zz_dataOut_payload_0_4446 < _zz_dataOut_payload_0_4449);
  assign _zz_dataOut_payload_0_4480 = (_zz_dataOut_payload_0_2992 < _zz_dataOut_payload_0_3007);
  assign _zz_dataOut_payload_0_4481 = (_zz_dataOut_payload_0_4480 ? _zz_dataOut_payload_0_2992 : _zz_dataOut_payload_0_3007);
  assign _zz_dataOut_payload_0_4482 = (_zz_dataOut_payload_0_4480 ? _zz_dataOut_payload_0_3007 : _zz_dataOut_payload_0_2992);
  assign _zz_dataOut_payload_0_4483 = (_zz_dataOut_payload_0_2993 < _zz_dataOut_payload_0_3006);
  assign _zz_dataOut_payload_0_4484 = (_zz_dataOut_payload_0_4483 ? _zz_dataOut_payload_0_2993 : _zz_dataOut_payload_0_3006);
  assign _zz_dataOut_payload_0_4485 = (_zz_dataOut_payload_0_4483 ? _zz_dataOut_payload_0_3006 : _zz_dataOut_payload_0_2993);
  assign _zz_dataOut_payload_0_4486 = (_zz_dataOut_payload_0_2994 < _zz_dataOut_payload_0_3005);
  assign _zz_dataOut_payload_0_4487 = (_zz_dataOut_payload_0_4486 ? _zz_dataOut_payload_0_2994 : _zz_dataOut_payload_0_3005);
  assign _zz_dataOut_payload_0_4488 = (_zz_dataOut_payload_0_4486 ? _zz_dataOut_payload_0_3005 : _zz_dataOut_payload_0_2994);
  assign _zz_dataOut_payload_0_4489 = (_zz_dataOut_payload_0_2995 < _zz_dataOut_payload_0_3004);
  assign _zz_dataOut_payload_0_4490 = (_zz_dataOut_payload_0_4489 ? _zz_dataOut_payload_0_2995 : _zz_dataOut_payload_0_3004);
  assign _zz_dataOut_payload_0_4491 = (_zz_dataOut_payload_0_4489 ? _zz_dataOut_payload_0_3004 : _zz_dataOut_payload_0_2995);
  assign _zz_dataOut_payload_0_4492 = (_zz_dataOut_payload_0_2996 < _zz_dataOut_payload_0_3003);
  assign _zz_dataOut_payload_0_4493 = (_zz_dataOut_payload_0_4492 ? _zz_dataOut_payload_0_2996 : _zz_dataOut_payload_0_3003);
  assign _zz_dataOut_payload_0_4494 = (_zz_dataOut_payload_0_4492 ? _zz_dataOut_payload_0_3003 : _zz_dataOut_payload_0_2996);
  assign _zz_dataOut_payload_0_4495 = (_zz_dataOut_payload_0_2997 < _zz_dataOut_payload_0_3002);
  assign _zz_dataOut_payload_0_4496 = (_zz_dataOut_payload_0_4495 ? _zz_dataOut_payload_0_2997 : _zz_dataOut_payload_0_3002);
  assign _zz_dataOut_payload_0_4497 = (_zz_dataOut_payload_0_4495 ? _zz_dataOut_payload_0_3002 : _zz_dataOut_payload_0_2997);
  assign _zz_dataOut_payload_0_4498 = (_zz_dataOut_payload_0_2998 < _zz_dataOut_payload_0_3001);
  assign _zz_dataOut_payload_0_4499 = (_zz_dataOut_payload_0_4498 ? _zz_dataOut_payload_0_2998 : _zz_dataOut_payload_0_3001);
  assign _zz_dataOut_payload_0_4500 = (_zz_dataOut_payload_0_4498 ? _zz_dataOut_payload_0_3001 : _zz_dataOut_payload_0_2998);
  assign _zz_dataOut_payload_0_4501 = (_zz_dataOut_payload_0_2999 < _zz_dataOut_payload_0_3000);
  assign _zz_dataOut_payload_0_4502 = (_zz_dataOut_payload_0_4501 ? _zz_dataOut_payload_0_2999 : _zz_dataOut_payload_0_3000);
  assign _zz_dataOut_payload_0_4503 = (_zz_dataOut_payload_0_4501 ? _zz_dataOut_payload_0_3000 : _zz_dataOut_payload_0_2999);
  assign _zz_dataOut_payload_0_4504 = (_zz_dataOut_payload_0_4481 < _zz_dataOut_payload_0_4493);
  assign _zz_dataOut_payload_0_4505 = (_zz_dataOut_payload_0_4504 ? _zz_dataOut_payload_0_4481 : _zz_dataOut_payload_0_4493);
  assign _zz_dataOut_payload_0_4506 = (_zz_dataOut_payload_0_4504 ? _zz_dataOut_payload_0_4493 : _zz_dataOut_payload_0_4481);
  assign _zz_dataOut_payload_0_4507 = (_zz_dataOut_payload_0_4484 < _zz_dataOut_payload_0_4496);
  assign _zz_dataOut_payload_0_4508 = (_zz_dataOut_payload_0_4507 ? _zz_dataOut_payload_0_4484 : _zz_dataOut_payload_0_4496);
  assign _zz_dataOut_payload_0_4509 = (_zz_dataOut_payload_0_4507 ? _zz_dataOut_payload_0_4496 : _zz_dataOut_payload_0_4484);
  assign _zz_dataOut_payload_0_4510 = (_zz_dataOut_payload_0_4487 < _zz_dataOut_payload_0_4499);
  assign _zz_dataOut_payload_0_4511 = (_zz_dataOut_payload_0_4510 ? _zz_dataOut_payload_0_4487 : _zz_dataOut_payload_0_4499);
  assign _zz_dataOut_payload_0_4512 = (_zz_dataOut_payload_0_4510 ? _zz_dataOut_payload_0_4499 : _zz_dataOut_payload_0_4487);
  assign _zz_dataOut_payload_0_4513 = (_zz_dataOut_payload_0_4490 < _zz_dataOut_payload_0_4502);
  assign _zz_dataOut_payload_0_4514 = (_zz_dataOut_payload_0_4513 ? _zz_dataOut_payload_0_4490 : _zz_dataOut_payload_0_4502);
  assign _zz_dataOut_payload_0_4515 = (_zz_dataOut_payload_0_4513 ? _zz_dataOut_payload_0_4502 : _zz_dataOut_payload_0_4490);
  assign _zz_dataOut_payload_0_4516 = (_zz_dataOut_payload_0_4505 < _zz_dataOut_payload_0_4511);
  assign _zz_dataOut_payload_0_4517 = (_zz_dataOut_payload_0_4516 ? _zz_dataOut_payload_0_4505 : _zz_dataOut_payload_0_4511);
  assign _zz_dataOut_payload_0_4518 = (_zz_dataOut_payload_0_4516 ? _zz_dataOut_payload_0_4511 : _zz_dataOut_payload_0_4505);
  assign _zz_dataOut_payload_0_4519 = (_zz_dataOut_payload_0_4508 < _zz_dataOut_payload_0_4514);
  assign _zz_dataOut_payload_0_4520 = (_zz_dataOut_payload_0_4519 ? _zz_dataOut_payload_0_4508 : _zz_dataOut_payload_0_4514);
  assign _zz_dataOut_payload_0_4521 = (_zz_dataOut_payload_0_4519 ? _zz_dataOut_payload_0_4514 : _zz_dataOut_payload_0_4508);
  assign _zz_dataOut_payload_0_4522 = (_zz_dataOut_payload_0_4517 < _zz_dataOut_payload_0_4520);
  assign _zz_dataOut_payload_0_4523 = (_zz_dataOut_payload_0_4518 < _zz_dataOut_payload_0_4521);
  assign _zz_dataOut_payload_0_4528 = (_zz_dataOut_payload_0_4506 < _zz_dataOut_payload_0_4512);
  assign _zz_dataOut_payload_0_4529 = (_zz_dataOut_payload_0_4528 ? _zz_dataOut_payload_0_4506 : _zz_dataOut_payload_0_4512);
  assign _zz_dataOut_payload_0_4530 = (_zz_dataOut_payload_0_4528 ? _zz_dataOut_payload_0_4512 : _zz_dataOut_payload_0_4506);
  assign _zz_dataOut_payload_0_4531 = (_zz_dataOut_payload_0_4509 < _zz_dataOut_payload_0_4515);
  assign _zz_dataOut_payload_0_4532 = (_zz_dataOut_payload_0_4531 ? _zz_dataOut_payload_0_4509 : _zz_dataOut_payload_0_4515);
  assign _zz_dataOut_payload_0_4533 = (_zz_dataOut_payload_0_4531 ? _zz_dataOut_payload_0_4515 : _zz_dataOut_payload_0_4509);
  assign _zz_dataOut_payload_0_4534 = (_zz_dataOut_payload_0_4529 < _zz_dataOut_payload_0_4532);
  assign _zz_dataOut_payload_0_4535 = (_zz_dataOut_payload_0_4530 < _zz_dataOut_payload_0_4533);
  assign _zz_dataOut_payload_0_4548 = (_zz_dataOut_payload_0_4503 < _zz_dataOut_payload_0_4491);
  assign _zz_dataOut_payload_0_4549 = (_zz_dataOut_payload_0_4548 ? _zz_dataOut_payload_0_4503 : _zz_dataOut_payload_0_4491);
  assign _zz_dataOut_payload_0_4550 = (_zz_dataOut_payload_0_4548 ? _zz_dataOut_payload_0_4491 : _zz_dataOut_payload_0_4503);
  assign _zz_dataOut_payload_0_4551 = (_zz_dataOut_payload_0_4500 < _zz_dataOut_payload_0_4488);
  assign _zz_dataOut_payload_0_4552 = (_zz_dataOut_payload_0_4551 ? _zz_dataOut_payload_0_4500 : _zz_dataOut_payload_0_4488);
  assign _zz_dataOut_payload_0_4553 = (_zz_dataOut_payload_0_4551 ? _zz_dataOut_payload_0_4488 : _zz_dataOut_payload_0_4500);
  assign _zz_dataOut_payload_0_4554 = (_zz_dataOut_payload_0_4497 < _zz_dataOut_payload_0_4485);
  assign _zz_dataOut_payload_0_4555 = (_zz_dataOut_payload_0_4554 ? _zz_dataOut_payload_0_4497 : _zz_dataOut_payload_0_4485);
  assign _zz_dataOut_payload_0_4556 = (_zz_dataOut_payload_0_4554 ? _zz_dataOut_payload_0_4485 : _zz_dataOut_payload_0_4497);
  assign _zz_dataOut_payload_0_4557 = (_zz_dataOut_payload_0_4494 < _zz_dataOut_payload_0_4482);
  assign _zz_dataOut_payload_0_4558 = (_zz_dataOut_payload_0_4557 ? _zz_dataOut_payload_0_4494 : _zz_dataOut_payload_0_4482);
  assign _zz_dataOut_payload_0_4559 = (_zz_dataOut_payload_0_4557 ? _zz_dataOut_payload_0_4482 : _zz_dataOut_payload_0_4494);
  assign _zz_dataOut_payload_0_4560 = (_zz_dataOut_payload_0_4549 < _zz_dataOut_payload_0_4555);
  assign _zz_dataOut_payload_0_4561 = (_zz_dataOut_payload_0_4560 ? _zz_dataOut_payload_0_4549 : _zz_dataOut_payload_0_4555);
  assign _zz_dataOut_payload_0_4562 = (_zz_dataOut_payload_0_4560 ? _zz_dataOut_payload_0_4555 : _zz_dataOut_payload_0_4549);
  assign _zz_dataOut_payload_0_4563 = (_zz_dataOut_payload_0_4552 < _zz_dataOut_payload_0_4558);
  assign _zz_dataOut_payload_0_4564 = (_zz_dataOut_payload_0_4563 ? _zz_dataOut_payload_0_4552 : _zz_dataOut_payload_0_4558);
  assign _zz_dataOut_payload_0_4565 = (_zz_dataOut_payload_0_4563 ? _zz_dataOut_payload_0_4558 : _zz_dataOut_payload_0_4552);
  assign _zz_dataOut_payload_0_4566 = (_zz_dataOut_payload_0_4561 < _zz_dataOut_payload_0_4564);
  assign _zz_dataOut_payload_0_4567 = (_zz_dataOut_payload_0_4562 < _zz_dataOut_payload_0_4565);
  assign _zz_dataOut_payload_0_4572 = (_zz_dataOut_payload_0_4550 < _zz_dataOut_payload_0_4556);
  assign _zz_dataOut_payload_0_4573 = (_zz_dataOut_payload_0_4572 ? _zz_dataOut_payload_0_4550 : _zz_dataOut_payload_0_4556);
  assign _zz_dataOut_payload_0_4574 = (_zz_dataOut_payload_0_4572 ? _zz_dataOut_payload_0_4556 : _zz_dataOut_payload_0_4550);
  assign _zz_dataOut_payload_0_4575 = (_zz_dataOut_payload_0_4553 < _zz_dataOut_payload_0_4559);
  assign _zz_dataOut_payload_0_4576 = (_zz_dataOut_payload_0_4575 ? _zz_dataOut_payload_0_4553 : _zz_dataOut_payload_0_4559);
  assign _zz_dataOut_payload_0_4577 = (_zz_dataOut_payload_0_4575 ? _zz_dataOut_payload_0_4559 : _zz_dataOut_payload_0_4553);
  assign _zz_dataOut_payload_0_4578 = (_zz_dataOut_payload_0_4573 < _zz_dataOut_payload_0_4576);
  assign _zz_dataOut_payload_0_4579 = (_zz_dataOut_payload_0_4574 < _zz_dataOut_payload_0_4577);
  assign _zz_dataOut_payload_0_4608 = (_zz_dataOut_payload_0_3008 < _zz_dataOut_payload_0_3023);
  assign _zz_dataOut_payload_0_4609 = (_zz_dataOut_payload_0_4608 ? _zz_dataOut_payload_0_3008 : _zz_dataOut_payload_0_3023);
  assign _zz_dataOut_payload_0_4610 = (_zz_dataOut_payload_0_4608 ? _zz_dataOut_payload_0_3023 : _zz_dataOut_payload_0_3008);
  assign _zz_dataOut_payload_0_4611 = (_zz_dataOut_payload_0_3009 < _zz_dataOut_payload_0_3022);
  assign _zz_dataOut_payload_0_4612 = (_zz_dataOut_payload_0_4611 ? _zz_dataOut_payload_0_3009 : _zz_dataOut_payload_0_3022);
  assign _zz_dataOut_payload_0_4613 = (_zz_dataOut_payload_0_4611 ? _zz_dataOut_payload_0_3022 : _zz_dataOut_payload_0_3009);
  assign _zz_dataOut_payload_0_4614 = (_zz_dataOut_payload_0_3010 < _zz_dataOut_payload_0_3021);
  assign _zz_dataOut_payload_0_4615 = (_zz_dataOut_payload_0_4614 ? _zz_dataOut_payload_0_3010 : _zz_dataOut_payload_0_3021);
  assign _zz_dataOut_payload_0_4616 = (_zz_dataOut_payload_0_4614 ? _zz_dataOut_payload_0_3021 : _zz_dataOut_payload_0_3010);
  assign _zz_dataOut_payload_0_4617 = (_zz_dataOut_payload_0_3011 < _zz_dataOut_payload_0_3020);
  assign _zz_dataOut_payload_0_4618 = (_zz_dataOut_payload_0_4617 ? _zz_dataOut_payload_0_3011 : _zz_dataOut_payload_0_3020);
  assign _zz_dataOut_payload_0_4619 = (_zz_dataOut_payload_0_4617 ? _zz_dataOut_payload_0_3020 : _zz_dataOut_payload_0_3011);
  assign _zz_dataOut_payload_0_4620 = (_zz_dataOut_payload_0_3012 < _zz_dataOut_payload_0_3019);
  assign _zz_dataOut_payload_0_4621 = (_zz_dataOut_payload_0_4620 ? _zz_dataOut_payload_0_3012 : _zz_dataOut_payload_0_3019);
  assign _zz_dataOut_payload_0_4622 = (_zz_dataOut_payload_0_4620 ? _zz_dataOut_payload_0_3019 : _zz_dataOut_payload_0_3012);
  assign _zz_dataOut_payload_0_4623 = (_zz_dataOut_payload_0_3013 < _zz_dataOut_payload_0_3018);
  assign _zz_dataOut_payload_0_4624 = (_zz_dataOut_payload_0_4623 ? _zz_dataOut_payload_0_3013 : _zz_dataOut_payload_0_3018);
  assign _zz_dataOut_payload_0_4625 = (_zz_dataOut_payload_0_4623 ? _zz_dataOut_payload_0_3018 : _zz_dataOut_payload_0_3013);
  assign _zz_dataOut_payload_0_4626 = (_zz_dataOut_payload_0_3014 < _zz_dataOut_payload_0_3017);
  assign _zz_dataOut_payload_0_4627 = (_zz_dataOut_payload_0_4626 ? _zz_dataOut_payload_0_3014 : _zz_dataOut_payload_0_3017);
  assign _zz_dataOut_payload_0_4628 = (_zz_dataOut_payload_0_4626 ? _zz_dataOut_payload_0_3017 : _zz_dataOut_payload_0_3014);
  assign _zz_dataOut_payload_0_4629 = (_zz_dataOut_payload_0_3015 < _zz_dataOut_payload_0_3016);
  assign _zz_dataOut_payload_0_4630 = (_zz_dataOut_payload_0_4629 ? _zz_dataOut_payload_0_3015 : _zz_dataOut_payload_0_3016);
  assign _zz_dataOut_payload_0_4631 = (_zz_dataOut_payload_0_4629 ? _zz_dataOut_payload_0_3016 : _zz_dataOut_payload_0_3015);
  assign _zz_dataOut_payload_0_4632 = (_zz_dataOut_payload_0_4609 < _zz_dataOut_payload_0_4621);
  assign _zz_dataOut_payload_0_4633 = (_zz_dataOut_payload_0_4632 ? _zz_dataOut_payload_0_4609 : _zz_dataOut_payload_0_4621);
  assign _zz_dataOut_payload_0_4634 = (_zz_dataOut_payload_0_4632 ? _zz_dataOut_payload_0_4621 : _zz_dataOut_payload_0_4609);
  assign _zz_dataOut_payload_0_4635 = (_zz_dataOut_payload_0_4612 < _zz_dataOut_payload_0_4624);
  assign _zz_dataOut_payload_0_4636 = (_zz_dataOut_payload_0_4635 ? _zz_dataOut_payload_0_4612 : _zz_dataOut_payload_0_4624);
  assign _zz_dataOut_payload_0_4637 = (_zz_dataOut_payload_0_4635 ? _zz_dataOut_payload_0_4624 : _zz_dataOut_payload_0_4612);
  assign _zz_dataOut_payload_0_4638 = (_zz_dataOut_payload_0_4615 < _zz_dataOut_payload_0_4627);
  assign _zz_dataOut_payload_0_4639 = (_zz_dataOut_payload_0_4638 ? _zz_dataOut_payload_0_4615 : _zz_dataOut_payload_0_4627);
  assign _zz_dataOut_payload_0_4640 = (_zz_dataOut_payload_0_4638 ? _zz_dataOut_payload_0_4627 : _zz_dataOut_payload_0_4615);
  assign _zz_dataOut_payload_0_4641 = (_zz_dataOut_payload_0_4618 < _zz_dataOut_payload_0_4630);
  assign _zz_dataOut_payload_0_4642 = (_zz_dataOut_payload_0_4641 ? _zz_dataOut_payload_0_4618 : _zz_dataOut_payload_0_4630);
  assign _zz_dataOut_payload_0_4643 = (_zz_dataOut_payload_0_4641 ? _zz_dataOut_payload_0_4630 : _zz_dataOut_payload_0_4618);
  assign _zz_dataOut_payload_0_4644 = (_zz_dataOut_payload_0_4633 < _zz_dataOut_payload_0_4639);
  assign _zz_dataOut_payload_0_4645 = (_zz_dataOut_payload_0_4644 ? _zz_dataOut_payload_0_4633 : _zz_dataOut_payload_0_4639);
  assign _zz_dataOut_payload_0_4646 = (_zz_dataOut_payload_0_4644 ? _zz_dataOut_payload_0_4639 : _zz_dataOut_payload_0_4633);
  assign _zz_dataOut_payload_0_4647 = (_zz_dataOut_payload_0_4636 < _zz_dataOut_payload_0_4642);
  assign _zz_dataOut_payload_0_4648 = (_zz_dataOut_payload_0_4647 ? _zz_dataOut_payload_0_4636 : _zz_dataOut_payload_0_4642);
  assign _zz_dataOut_payload_0_4649 = (_zz_dataOut_payload_0_4647 ? _zz_dataOut_payload_0_4642 : _zz_dataOut_payload_0_4636);
  assign _zz_dataOut_payload_0_4650 = (_zz_dataOut_payload_0_4645 < _zz_dataOut_payload_0_4648);
  assign _zz_dataOut_payload_0_4651 = (_zz_dataOut_payload_0_4646 < _zz_dataOut_payload_0_4649);
  assign _zz_dataOut_payload_0_4656 = (_zz_dataOut_payload_0_4634 < _zz_dataOut_payload_0_4640);
  assign _zz_dataOut_payload_0_4657 = (_zz_dataOut_payload_0_4656 ? _zz_dataOut_payload_0_4634 : _zz_dataOut_payload_0_4640);
  assign _zz_dataOut_payload_0_4658 = (_zz_dataOut_payload_0_4656 ? _zz_dataOut_payload_0_4640 : _zz_dataOut_payload_0_4634);
  assign _zz_dataOut_payload_0_4659 = (_zz_dataOut_payload_0_4637 < _zz_dataOut_payload_0_4643);
  assign _zz_dataOut_payload_0_4660 = (_zz_dataOut_payload_0_4659 ? _zz_dataOut_payload_0_4637 : _zz_dataOut_payload_0_4643);
  assign _zz_dataOut_payload_0_4661 = (_zz_dataOut_payload_0_4659 ? _zz_dataOut_payload_0_4643 : _zz_dataOut_payload_0_4637);
  assign _zz_dataOut_payload_0_4662 = (_zz_dataOut_payload_0_4657 < _zz_dataOut_payload_0_4660);
  assign _zz_dataOut_payload_0_4663 = (_zz_dataOut_payload_0_4658 < _zz_dataOut_payload_0_4661);
  assign _zz_dataOut_payload_0_4676 = (_zz_dataOut_payload_0_4631 < _zz_dataOut_payload_0_4619);
  assign _zz_dataOut_payload_0_4677 = (_zz_dataOut_payload_0_4676 ? _zz_dataOut_payload_0_4631 : _zz_dataOut_payload_0_4619);
  assign _zz_dataOut_payload_0_4678 = (_zz_dataOut_payload_0_4676 ? _zz_dataOut_payload_0_4619 : _zz_dataOut_payload_0_4631);
  assign _zz_dataOut_payload_0_4679 = (_zz_dataOut_payload_0_4628 < _zz_dataOut_payload_0_4616);
  assign _zz_dataOut_payload_0_4680 = (_zz_dataOut_payload_0_4679 ? _zz_dataOut_payload_0_4628 : _zz_dataOut_payload_0_4616);
  assign _zz_dataOut_payload_0_4681 = (_zz_dataOut_payload_0_4679 ? _zz_dataOut_payload_0_4616 : _zz_dataOut_payload_0_4628);
  assign _zz_dataOut_payload_0_4682 = (_zz_dataOut_payload_0_4625 < _zz_dataOut_payload_0_4613);
  assign _zz_dataOut_payload_0_4683 = (_zz_dataOut_payload_0_4682 ? _zz_dataOut_payload_0_4625 : _zz_dataOut_payload_0_4613);
  assign _zz_dataOut_payload_0_4684 = (_zz_dataOut_payload_0_4682 ? _zz_dataOut_payload_0_4613 : _zz_dataOut_payload_0_4625);
  assign _zz_dataOut_payload_0_4685 = (_zz_dataOut_payload_0_4622 < _zz_dataOut_payload_0_4610);
  assign _zz_dataOut_payload_0_4686 = (_zz_dataOut_payload_0_4685 ? _zz_dataOut_payload_0_4622 : _zz_dataOut_payload_0_4610);
  assign _zz_dataOut_payload_0_4687 = (_zz_dataOut_payload_0_4685 ? _zz_dataOut_payload_0_4610 : _zz_dataOut_payload_0_4622);
  assign _zz_dataOut_payload_0_4688 = (_zz_dataOut_payload_0_4677 < _zz_dataOut_payload_0_4683);
  assign _zz_dataOut_payload_0_4689 = (_zz_dataOut_payload_0_4688 ? _zz_dataOut_payload_0_4677 : _zz_dataOut_payload_0_4683);
  assign _zz_dataOut_payload_0_4690 = (_zz_dataOut_payload_0_4688 ? _zz_dataOut_payload_0_4683 : _zz_dataOut_payload_0_4677);
  assign _zz_dataOut_payload_0_4691 = (_zz_dataOut_payload_0_4680 < _zz_dataOut_payload_0_4686);
  assign _zz_dataOut_payload_0_4692 = (_zz_dataOut_payload_0_4691 ? _zz_dataOut_payload_0_4680 : _zz_dataOut_payload_0_4686);
  assign _zz_dataOut_payload_0_4693 = (_zz_dataOut_payload_0_4691 ? _zz_dataOut_payload_0_4686 : _zz_dataOut_payload_0_4680);
  assign _zz_dataOut_payload_0_4694 = (_zz_dataOut_payload_0_4689 < _zz_dataOut_payload_0_4692);
  assign _zz_dataOut_payload_0_4695 = (_zz_dataOut_payload_0_4690 < _zz_dataOut_payload_0_4693);
  assign _zz_dataOut_payload_0_4700 = (_zz_dataOut_payload_0_4678 < _zz_dataOut_payload_0_4684);
  assign _zz_dataOut_payload_0_4701 = (_zz_dataOut_payload_0_4700 ? _zz_dataOut_payload_0_4678 : _zz_dataOut_payload_0_4684);
  assign _zz_dataOut_payload_0_4702 = (_zz_dataOut_payload_0_4700 ? _zz_dataOut_payload_0_4684 : _zz_dataOut_payload_0_4678);
  assign _zz_dataOut_payload_0_4703 = (_zz_dataOut_payload_0_4681 < _zz_dataOut_payload_0_4687);
  assign _zz_dataOut_payload_0_4704 = (_zz_dataOut_payload_0_4703 ? _zz_dataOut_payload_0_4681 : _zz_dataOut_payload_0_4687);
  assign _zz_dataOut_payload_0_4705 = (_zz_dataOut_payload_0_4703 ? _zz_dataOut_payload_0_4687 : _zz_dataOut_payload_0_4681);
  assign _zz_dataOut_payload_0_4706 = (_zz_dataOut_payload_0_4701 < _zz_dataOut_payload_0_4704);
  assign _zz_dataOut_payload_0_4707 = (_zz_dataOut_payload_0_4702 < _zz_dataOut_payload_0_4705);
  assign _zz_dataOut_payload_0_4736 = (_zz_dataOut_payload_0_3024 < _zz_dataOut_payload_0_3039);
  assign _zz_dataOut_payload_0_4737 = (_zz_dataOut_payload_0_4736 ? _zz_dataOut_payload_0_3024 : _zz_dataOut_payload_0_3039);
  assign _zz_dataOut_payload_0_4738 = (_zz_dataOut_payload_0_4736 ? _zz_dataOut_payload_0_3039 : _zz_dataOut_payload_0_3024);
  assign _zz_dataOut_payload_0_4739 = (_zz_dataOut_payload_0_3025 < _zz_dataOut_payload_0_3038);
  assign _zz_dataOut_payload_0_4740 = (_zz_dataOut_payload_0_4739 ? _zz_dataOut_payload_0_3025 : _zz_dataOut_payload_0_3038);
  assign _zz_dataOut_payload_0_4741 = (_zz_dataOut_payload_0_4739 ? _zz_dataOut_payload_0_3038 : _zz_dataOut_payload_0_3025);
  assign _zz_dataOut_payload_0_4742 = (_zz_dataOut_payload_0_3026 < _zz_dataOut_payload_0_3037);
  assign _zz_dataOut_payload_0_4743 = (_zz_dataOut_payload_0_4742 ? _zz_dataOut_payload_0_3026 : _zz_dataOut_payload_0_3037);
  assign _zz_dataOut_payload_0_4744 = (_zz_dataOut_payload_0_4742 ? _zz_dataOut_payload_0_3037 : _zz_dataOut_payload_0_3026);
  assign _zz_dataOut_payload_0_4745 = (_zz_dataOut_payload_0_3027 < _zz_dataOut_payload_0_3036);
  assign _zz_dataOut_payload_0_4746 = (_zz_dataOut_payload_0_4745 ? _zz_dataOut_payload_0_3027 : _zz_dataOut_payload_0_3036);
  assign _zz_dataOut_payload_0_4747 = (_zz_dataOut_payload_0_4745 ? _zz_dataOut_payload_0_3036 : _zz_dataOut_payload_0_3027);
  assign _zz_dataOut_payload_0_4748 = (_zz_dataOut_payload_0_3028 < _zz_dataOut_payload_0_3035);
  assign _zz_dataOut_payload_0_4749 = (_zz_dataOut_payload_0_4748 ? _zz_dataOut_payload_0_3028 : _zz_dataOut_payload_0_3035);
  assign _zz_dataOut_payload_0_4750 = (_zz_dataOut_payload_0_4748 ? _zz_dataOut_payload_0_3035 : _zz_dataOut_payload_0_3028);
  assign _zz_dataOut_payload_0_4751 = (_zz_dataOut_payload_0_3029 < _zz_dataOut_payload_0_3034);
  assign _zz_dataOut_payload_0_4752 = (_zz_dataOut_payload_0_4751 ? _zz_dataOut_payload_0_3029 : _zz_dataOut_payload_0_3034);
  assign _zz_dataOut_payload_0_4753 = (_zz_dataOut_payload_0_4751 ? _zz_dataOut_payload_0_3034 : _zz_dataOut_payload_0_3029);
  assign _zz_dataOut_payload_0_4754 = (_zz_dataOut_payload_0_3030 < _zz_dataOut_payload_0_3033);
  assign _zz_dataOut_payload_0_4755 = (_zz_dataOut_payload_0_4754 ? _zz_dataOut_payload_0_3030 : _zz_dataOut_payload_0_3033);
  assign _zz_dataOut_payload_0_4756 = (_zz_dataOut_payload_0_4754 ? _zz_dataOut_payload_0_3033 : _zz_dataOut_payload_0_3030);
  assign _zz_dataOut_payload_0_4757 = (_zz_dataOut_payload_0_3031 < _zz_dataOut_payload_0_3032);
  assign _zz_dataOut_payload_0_4758 = (_zz_dataOut_payload_0_4757 ? _zz_dataOut_payload_0_3031 : _zz_dataOut_payload_0_3032);
  assign _zz_dataOut_payload_0_4759 = (_zz_dataOut_payload_0_4757 ? _zz_dataOut_payload_0_3032 : _zz_dataOut_payload_0_3031);
  assign _zz_dataOut_payload_0_4760 = (_zz_dataOut_payload_0_4737 < _zz_dataOut_payload_0_4749);
  assign _zz_dataOut_payload_0_4761 = (_zz_dataOut_payload_0_4760 ? _zz_dataOut_payload_0_4737 : _zz_dataOut_payload_0_4749);
  assign _zz_dataOut_payload_0_4762 = (_zz_dataOut_payload_0_4760 ? _zz_dataOut_payload_0_4749 : _zz_dataOut_payload_0_4737);
  assign _zz_dataOut_payload_0_4763 = (_zz_dataOut_payload_0_4740 < _zz_dataOut_payload_0_4752);
  assign _zz_dataOut_payload_0_4764 = (_zz_dataOut_payload_0_4763 ? _zz_dataOut_payload_0_4740 : _zz_dataOut_payload_0_4752);
  assign _zz_dataOut_payload_0_4765 = (_zz_dataOut_payload_0_4763 ? _zz_dataOut_payload_0_4752 : _zz_dataOut_payload_0_4740);
  assign _zz_dataOut_payload_0_4766 = (_zz_dataOut_payload_0_4743 < _zz_dataOut_payload_0_4755);
  assign _zz_dataOut_payload_0_4767 = (_zz_dataOut_payload_0_4766 ? _zz_dataOut_payload_0_4743 : _zz_dataOut_payload_0_4755);
  assign _zz_dataOut_payload_0_4768 = (_zz_dataOut_payload_0_4766 ? _zz_dataOut_payload_0_4755 : _zz_dataOut_payload_0_4743);
  assign _zz_dataOut_payload_0_4769 = (_zz_dataOut_payload_0_4746 < _zz_dataOut_payload_0_4758);
  assign _zz_dataOut_payload_0_4770 = (_zz_dataOut_payload_0_4769 ? _zz_dataOut_payload_0_4746 : _zz_dataOut_payload_0_4758);
  assign _zz_dataOut_payload_0_4771 = (_zz_dataOut_payload_0_4769 ? _zz_dataOut_payload_0_4758 : _zz_dataOut_payload_0_4746);
  assign _zz_dataOut_payload_0_4772 = (_zz_dataOut_payload_0_4761 < _zz_dataOut_payload_0_4767);
  assign _zz_dataOut_payload_0_4773 = (_zz_dataOut_payload_0_4772 ? _zz_dataOut_payload_0_4761 : _zz_dataOut_payload_0_4767);
  assign _zz_dataOut_payload_0_4774 = (_zz_dataOut_payload_0_4772 ? _zz_dataOut_payload_0_4767 : _zz_dataOut_payload_0_4761);
  assign _zz_dataOut_payload_0_4775 = (_zz_dataOut_payload_0_4764 < _zz_dataOut_payload_0_4770);
  assign _zz_dataOut_payload_0_4776 = (_zz_dataOut_payload_0_4775 ? _zz_dataOut_payload_0_4764 : _zz_dataOut_payload_0_4770);
  assign _zz_dataOut_payload_0_4777 = (_zz_dataOut_payload_0_4775 ? _zz_dataOut_payload_0_4770 : _zz_dataOut_payload_0_4764);
  assign _zz_dataOut_payload_0_4778 = (_zz_dataOut_payload_0_4773 < _zz_dataOut_payload_0_4776);
  assign _zz_dataOut_payload_0_4779 = (_zz_dataOut_payload_0_4774 < _zz_dataOut_payload_0_4777);
  assign _zz_dataOut_payload_0_4784 = (_zz_dataOut_payload_0_4762 < _zz_dataOut_payload_0_4768);
  assign _zz_dataOut_payload_0_4785 = (_zz_dataOut_payload_0_4784 ? _zz_dataOut_payload_0_4762 : _zz_dataOut_payload_0_4768);
  assign _zz_dataOut_payload_0_4786 = (_zz_dataOut_payload_0_4784 ? _zz_dataOut_payload_0_4768 : _zz_dataOut_payload_0_4762);
  assign _zz_dataOut_payload_0_4787 = (_zz_dataOut_payload_0_4765 < _zz_dataOut_payload_0_4771);
  assign _zz_dataOut_payload_0_4788 = (_zz_dataOut_payload_0_4787 ? _zz_dataOut_payload_0_4765 : _zz_dataOut_payload_0_4771);
  assign _zz_dataOut_payload_0_4789 = (_zz_dataOut_payload_0_4787 ? _zz_dataOut_payload_0_4771 : _zz_dataOut_payload_0_4765);
  assign _zz_dataOut_payload_0_4790 = (_zz_dataOut_payload_0_4785 < _zz_dataOut_payload_0_4788);
  assign _zz_dataOut_payload_0_4791 = (_zz_dataOut_payload_0_4786 < _zz_dataOut_payload_0_4789);
  assign _zz_dataOut_payload_0_4804 = (_zz_dataOut_payload_0_4759 < _zz_dataOut_payload_0_4747);
  assign _zz_dataOut_payload_0_4805 = (_zz_dataOut_payload_0_4804 ? _zz_dataOut_payload_0_4759 : _zz_dataOut_payload_0_4747);
  assign _zz_dataOut_payload_0_4806 = (_zz_dataOut_payload_0_4804 ? _zz_dataOut_payload_0_4747 : _zz_dataOut_payload_0_4759);
  assign _zz_dataOut_payload_0_4807 = (_zz_dataOut_payload_0_4756 < _zz_dataOut_payload_0_4744);
  assign _zz_dataOut_payload_0_4808 = (_zz_dataOut_payload_0_4807 ? _zz_dataOut_payload_0_4756 : _zz_dataOut_payload_0_4744);
  assign _zz_dataOut_payload_0_4809 = (_zz_dataOut_payload_0_4807 ? _zz_dataOut_payload_0_4744 : _zz_dataOut_payload_0_4756);
  assign _zz_dataOut_payload_0_4810 = (_zz_dataOut_payload_0_4753 < _zz_dataOut_payload_0_4741);
  assign _zz_dataOut_payload_0_4811 = (_zz_dataOut_payload_0_4810 ? _zz_dataOut_payload_0_4753 : _zz_dataOut_payload_0_4741);
  assign _zz_dataOut_payload_0_4812 = (_zz_dataOut_payload_0_4810 ? _zz_dataOut_payload_0_4741 : _zz_dataOut_payload_0_4753);
  assign _zz_dataOut_payload_0_4813 = (_zz_dataOut_payload_0_4750 < _zz_dataOut_payload_0_4738);
  assign _zz_dataOut_payload_0_4814 = (_zz_dataOut_payload_0_4813 ? _zz_dataOut_payload_0_4750 : _zz_dataOut_payload_0_4738);
  assign _zz_dataOut_payload_0_4815 = (_zz_dataOut_payload_0_4813 ? _zz_dataOut_payload_0_4738 : _zz_dataOut_payload_0_4750);
  assign _zz_dataOut_payload_0_4816 = (_zz_dataOut_payload_0_4805 < _zz_dataOut_payload_0_4811);
  assign _zz_dataOut_payload_0_4817 = (_zz_dataOut_payload_0_4816 ? _zz_dataOut_payload_0_4805 : _zz_dataOut_payload_0_4811);
  assign _zz_dataOut_payload_0_4818 = (_zz_dataOut_payload_0_4816 ? _zz_dataOut_payload_0_4811 : _zz_dataOut_payload_0_4805);
  assign _zz_dataOut_payload_0_4819 = (_zz_dataOut_payload_0_4808 < _zz_dataOut_payload_0_4814);
  assign _zz_dataOut_payload_0_4820 = (_zz_dataOut_payload_0_4819 ? _zz_dataOut_payload_0_4808 : _zz_dataOut_payload_0_4814);
  assign _zz_dataOut_payload_0_4821 = (_zz_dataOut_payload_0_4819 ? _zz_dataOut_payload_0_4814 : _zz_dataOut_payload_0_4808);
  assign _zz_dataOut_payload_0_4822 = (_zz_dataOut_payload_0_4817 < _zz_dataOut_payload_0_4820);
  assign _zz_dataOut_payload_0_4823 = (_zz_dataOut_payload_0_4818 < _zz_dataOut_payload_0_4821);
  assign _zz_dataOut_payload_0_4828 = (_zz_dataOut_payload_0_4806 < _zz_dataOut_payload_0_4812);
  assign _zz_dataOut_payload_0_4829 = (_zz_dataOut_payload_0_4828 ? _zz_dataOut_payload_0_4806 : _zz_dataOut_payload_0_4812);
  assign _zz_dataOut_payload_0_4830 = (_zz_dataOut_payload_0_4828 ? _zz_dataOut_payload_0_4812 : _zz_dataOut_payload_0_4806);
  assign _zz_dataOut_payload_0_4831 = (_zz_dataOut_payload_0_4809 < _zz_dataOut_payload_0_4815);
  assign _zz_dataOut_payload_0_4832 = (_zz_dataOut_payload_0_4831 ? _zz_dataOut_payload_0_4809 : _zz_dataOut_payload_0_4815);
  assign _zz_dataOut_payload_0_4833 = (_zz_dataOut_payload_0_4831 ? _zz_dataOut_payload_0_4815 : _zz_dataOut_payload_0_4809);
  assign _zz_dataOut_payload_0_4834 = (_zz_dataOut_payload_0_4829 < _zz_dataOut_payload_0_4832);
  assign _zz_dataOut_payload_0_4835 = (_zz_dataOut_payload_0_4830 < _zz_dataOut_payload_0_4833);
  assign _zz_dataOut_payload_0_4864 = (_zz_dataOut_payload_0_3040 < _zz_dataOut_payload_0_3055);
  assign _zz_dataOut_payload_0_4865 = (_zz_dataOut_payload_0_4864 ? _zz_dataOut_payload_0_3040 : _zz_dataOut_payload_0_3055);
  assign _zz_dataOut_payload_0_4866 = (_zz_dataOut_payload_0_4864 ? _zz_dataOut_payload_0_3055 : _zz_dataOut_payload_0_3040);
  assign _zz_dataOut_payload_0_4867 = (_zz_dataOut_payload_0_3041 < _zz_dataOut_payload_0_3054);
  assign _zz_dataOut_payload_0_4868 = (_zz_dataOut_payload_0_4867 ? _zz_dataOut_payload_0_3041 : _zz_dataOut_payload_0_3054);
  assign _zz_dataOut_payload_0_4869 = (_zz_dataOut_payload_0_4867 ? _zz_dataOut_payload_0_3054 : _zz_dataOut_payload_0_3041);
  assign _zz_dataOut_payload_0_4870 = (_zz_dataOut_payload_0_3042 < _zz_dataOut_payload_0_3053);
  assign _zz_dataOut_payload_0_4871 = (_zz_dataOut_payload_0_4870 ? _zz_dataOut_payload_0_3042 : _zz_dataOut_payload_0_3053);
  assign _zz_dataOut_payload_0_4872 = (_zz_dataOut_payload_0_4870 ? _zz_dataOut_payload_0_3053 : _zz_dataOut_payload_0_3042);
  assign _zz_dataOut_payload_0_4873 = (_zz_dataOut_payload_0_3043 < _zz_dataOut_payload_0_3052);
  assign _zz_dataOut_payload_0_4874 = (_zz_dataOut_payload_0_4873 ? _zz_dataOut_payload_0_3043 : _zz_dataOut_payload_0_3052);
  assign _zz_dataOut_payload_0_4875 = (_zz_dataOut_payload_0_4873 ? _zz_dataOut_payload_0_3052 : _zz_dataOut_payload_0_3043);
  assign _zz_dataOut_payload_0_4876 = (_zz_dataOut_payload_0_3044 < _zz_dataOut_payload_0_3051);
  assign _zz_dataOut_payload_0_4877 = (_zz_dataOut_payload_0_4876 ? _zz_dataOut_payload_0_3044 : _zz_dataOut_payload_0_3051);
  assign _zz_dataOut_payload_0_4878 = (_zz_dataOut_payload_0_4876 ? _zz_dataOut_payload_0_3051 : _zz_dataOut_payload_0_3044);
  assign _zz_dataOut_payload_0_4879 = (_zz_dataOut_payload_0_3045 < _zz_dataOut_payload_0_3050);
  assign _zz_dataOut_payload_0_4880 = (_zz_dataOut_payload_0_4879 ? _zz_dataOut_payload_0_3045 : _zz_dataOut_payload_0_3050);
  assign _zz_dataOut_payload_0_4881 = (_zz_dataOut_payload_0_4879 ? _zz_dataOut_payload_0_3050 : _zz_dataOut_payload_0_3045);
  assign _zz_dataOut_payload_0_4882 = (_zz_dataOut_payload_0_3046 < _zz_dataOut_payload_0_3049);
  assign _zz_dataOut_payload_0_4883 = (_zz_dataOut_payload_0_4882 ? _zz_dataOut_payload_0_3046 : _zz_dataOut_payload_0_3049);
  assign _zz_dataOut_payload_0_4884 = (_zz_dataOut_payload_0_4882 ? _zz_dataOut_payload_0_3049 : _zz_dataOut_payload_0_3046);
  assign _zz_dataOut_payload_0_4885 = (_zz_dataOut_payload_0_3047 < _zz_dataOut_payload_0_3048);
  assign _zz_dataOut_payload_0_4886 = (_zz_dataOut_payload_0_4885 ? _zz_dataOut_payload_0_3047 : _zz_dataOut_payload_0_3048);
  assign _zz_dataOut_payload_0_4887 = (_zz_dataOut_payload_0_4885 ? _zz_dataOut_payload_0_3048 : _zz_dataOut_payload_0_3047);
  assign _zz_dataOut_payload_0_4888 = (_zz_dataOut_payload_0_4865 < _zz_dataOut_payload_0_4877);
  assign _zz_dataOut_payload_0_4889 = (_zz_dataOut_payload_0_4888 ? _zz_dataOut_payload_0_4865 : _zz_dataOut_payload_0_4877);
  assign _zz_dataOut_payload_0_4890 = (_zz_dataOut_payload_0_4888 ? _zz_dataOut_payload_0_4877 : _zz_dataOut_payload_0_4865);
  assign _zz_dataOut_payload_0_4891 = (_zz_dataOut_payload_0_4868 < _zz_dataOut_payload_0_4880);
  assign _zz_dataOut_payload_0_4892 = (_zz_dataOut_payload_0_4891 ? _zz_dataOut_payload_0_4868 : _zz_dataOut_payload_0_4880);
  assign _zz_dataOut_payload_0_4893 = (_zz_dataOut_payload_0_4891 ? _zz_dataOut_payload_0_4880 : _zz_dataOut_payload_0_4868);
  assign _zz_dataOut_payload_0_4894 = (_zz_dataOut_payload_0_4871 < _zz_dataOut_payload_0_4883);
  assign _zz_dataOut_payload_0_4895 = (_zz_dataOut_payload_0_4894 ? _zz_dataOut_payload_0_4871 : _zz_dataOut_payload_0_4883);
  assign _zz_dataOut_payload_0_4896 = (_zz_dataOut_payload_0_4894 ? _zz_dataOut_payload_0_4883 : _zz_dataOut_payload_0_4871);
  assign _zz_dataOut_payload_0_4897 = (_zz_dataOut_payload_0_4874 < _zz_dataOut_payload_0_4886);
  assign _zz_dataOut_payload_0_4898 = (_zz_dataOut_payload_0_4897 ? _zz_dataOut_payload_0_4874 : _zz_dataOut_payload_0_4886);
  assign _zz_dataOut_payload_0_4899 = (_zz_dataOut_payload_0_4897 ? _zz_dataOut_payload_0_4886 : _zz_dataOut_payload_0_4874);
  assign _zz_dataOut_payload_0_4900 = (_zz_dataOut_payload_0_4889 < _zz_dataOut_payload_0_4895);
  assign _zz_dataOut_payload_0_4901 = (_zz_dataOut_payload_0_4900 ? _zz_dataOut_payload_0_4889 : _zz_dataOut_payload_0_4895);
  assign _zz_dataOut_payload_0_4902 = (_zz_dataOut_payload_0_4900 ? _zz_dataOut_payload_0_4895 : _zz_dataOut_payload_0_4889);
  assign _zz_dataOut_payload_0_4903 = (_zz_dataOut_payload_0_4892 < _zz_dataOut_payload_0_4898);
  assign _zz_dataOut_payload_0_4904 = (_zz_dataOut_payload_0_4903 ? _zz_dataOut_payload_0_4892 : _zz_dataOut_payload_0_4898);
  assign _zz_dataOut_payload_0_4905 = (_zz_dataOut_payload_0_4903 ? _zz_dataOut_payload_0_4898 : _zz_dataOut_payload_0_4892);
  assign _zz_dataOut_payload_0_4906 = (_zz_dataOut_payload_0_4901 < _zz_dataOut_payload_0_4904);
  assign _zz_dataOut_payload_0_4907 = (_zz_dataOut_payload_0_4902 < _zz_dataOut_payload_0_4905);
  assign _zz_dataOut_payload_0_4912 = (_zz_dataOut_payload_0_4890 < _zz_dataOut_payload_0_4896);
  assign _zz_dataOut_payload_0_4913 = (_zz_dataOut_payload_0_4912 ? _zz_dataOut_payload_0_4890 : _zz_dataOut_payload_0_4896);
  assign _zz_dataOut_payload_0_4914 = (_zz_dataOut_payload_0_4912 ? _zz_dataOut_payload_0_4896 : _zz_dataOut_payload_0_4890);
  assign _zz_dataOut_payload_0_4915 = (_zz_dataOut_payload_0_4893 < _zz_dataOut_payload_0_4899);
  assign _zz_dataOut_payload_0_4916 = (_zz_dataOut_payload_0_4915 ? _zz_dataOut_payload_0_4893 : _zz_dataOut_payload_0_4899);
  assign _zz_dataOut_payload_0_4917 = (_zz_dataOut_payload_0_4915 ? _zz_dataOut_payload_0_4899 : _zz_dataOut_payload_0_4893);
  assign _zz_dataOut_payload_0_4918 = (_zz_dataOut_payload_0_4913 < _zz_dataOut_payload_0_4916);
  assign _zz_dataOut_payload_0_4919 = (_zz_dataOut_payload_0_4914 < _zz_dataOut_payload_0_4917);
  assign _zz_dataOut_payload_0_4932 = (_zz_dataOut_payload_0_4887 < _zz_dataOut_payload_0_4875);
  assign _zz_dataOut_payload_0_4933 = (_zz_dataOut_payload_0_4932 ? _zz_dataOut_payload_0_4887 : _zz_dataOut_payload_0_4875);
  assign _zz_dataOut_payload_0_4934 = (_zz_dataOut_payload_0_4932 ? _zz_dataOut_payload_0_4875 : _zz_dataOut_payload_0_4887);
  assign _zz_dataOut_payload_0_4935 = (_zz_dataOut_payload_0_4884 < _zz_dataOut_payload_0_4872);
  assign _zz_dataOut_payload_0_4936 = (_zz_dataOut_payload_0_4935 ? _zz_dataOut_payload_0_4884 : _zz_dataOut_payload_0_4872);
  assign _zz_dataOut_payload_0_4937 = (_zz_dataOut_payload_0_4935 ? _zz_dataOut_payload_0_4872 : _zz_dataOut_payload_0_4884);
  assign _zz_dataOut_payload_0_4938 = (_zz_dataOut_payload_0_4881 < _zz_dataOut_payload_0_4869);
  assign _zz_dataOut_payload_0_4939 = (_zz_dataOut_payload_0_4938 ? _zz_dataOut_payload_0_4881 : _zz_dataOut_payload_0_4869);
  assign _zz_dataOut_payload_0_4940 = (_zz_dataOut_payload_0_4938 ? _zz_dataOut_payload_0_4869 : _zz_dataOut_payload_0_4881);
  assign _zz_dataOut_payload_0_4941 = (_zz_dataOut_payload_0_4878 < _zz_dataOut_payload_0_4866);
  assign _zz_dataOut_payload_0_4942 = (_zz_dataOut_payload_0_4941 ? _zz_dataOut_payload_0_4878 : _zz_dataOut_payload_0_4866);
  assign _zz_dataOut_payload_0_4943 = (_zz_dataOut_payload_0_4941 ? _zz_dataOut_payload_0_4866 : _zz_dataOut_payload_0_4878);
  assign _zz_dataOut_payload_0_4944 = (_zz_dataOut_payload_0_4933 < _zz_dataOut_payload_0_4939);
  assign _zz_dataOut_payload_0_4945 = (_zz_dataOut_payload_0_4944 ? _zz_dataOut_payload_0_4933 : _zz_dataOut_payload_0_4939);
  assign _zz_dataOut_payload_0_4946 = (_zz_dataOut_payload_0_4944 ? _zz_dataOut_payload_0_4939 : _zz_dataOut_payload_0_4933);
  assign _zz_dataOut_payload_0_4947 = (_zz_dataOut_payload_0_4936 < _zz_dataOut_payload_0_4942);
  assign _zz_dataOut_payload_0_4948 = (_zz_dataOut_payload_0_4947 ? _zz_dataOut_payload_0_4936 : _zz_dataOut_payload_0_4942);
  assign _zz_dataOut_payload_0_4949 = (_zz_dataOut_payload_0_4947 ? _zz_dataOut_payload_0_4942 : _zz_dataOut_payload_0_4936);
  assign _zz_dataOut_payload_0_4950 = (_zz_dataOut_payload_0_4945 < _zz_dataOut_payload_0_4948);
  assign _zz_dataOut_payload_0_4951 = (_zz_dataOut_payload_0_4946 < _zz_dataOut_payload_0_4949);
  assign _zz_dataOut_payload_0_4956 = (_zz_dataOut_payload_0_4934 < _zz_dataOut_payload_0_4940);
  assign _zz_dataOut_payload_0_4957 = (_zz_dataOut_payload_0_4956 ? _zz_dataOut_payload_0_4934 : _zz_dataOut_payload_0_4940);
  assign _zz_dataOut_payload_0_4958 = (_zz_dataOut_payload_0_4956 ? _zz_dataOut_payload_0_4940 : _zz_dataOut_payload_0_4934);
  assign _zz_dataOut_payload_0_4959 = (_zz_dataOut_payload_0_4937 < _zz_dataOut_payload_0_4943);
  assign _zz_dataOut_payload_0_4960 = (_zz_dataOut_payload_0_4959 ? _zz_dataOut_payload_0_4937 : _zz_dataOut_payload_0_4943);
  assign _zz_dataOut_payload_0_4961 = (_zz_dataOut_payload_0_4959 ? _zz_dataOut_payload_0_4943 : _zz_dataOut_payload_0_4937);
  assign _zz_dataOut_payload_0_4962 = (_zz_dataOut_payload_0_4957 < _zz_dataOut_payload_0_4960);
  assign _zz_dataOut_payload_0_4963 = (_zz_dataOut_payload_0_4958 < _zz_dataOut_payload_0_4961);
  assign _zz_dataOut_payload_0_4992 = (_zz_dataOut_payload_0_3056 < _zz_dataOut_payload_0_3071);
  assign _zz_dataOut_payload_0_4993 = (_zz_dataOut_payload_0_4992 ? _zz_dataOut_payload_0_3056 : _zz_dataOut_payload_0_3071);
  assign _zz_dataOut_payload_0_4994 = (_zz_dataOut_payload_0_4992 ? _zz_dataOut_payload_0_3071 : _zz_dataOut_payload_0_3056);
  assign _zz_dataOut_payload_0_4995 = (_zz_dataOut_payload_0_3057 < _zz_dataOut_payload_0_3070);
  assign _zz_dataOut_payload_0_4996 = (_zz_dataOut_payload_0_4995 ? _zz_dataOut_payload_0_3057 : _zz_dataOut_payload_0_3070);
  assign _zz_dataOut_payload_0_4997 = (_zz_dataOut_payload_0_4995 ? _zz_dataOut_payload_0_3070 : _zz_dataOut_payload_0_3057);
  assign _zz_dataOut_payload_0_4998 = (_zz_dataOut_payload_0_3058 < _zz_dataOut_payload_0_3069);
  assign _zz_dataOut_payload_0_4999 = (_zz_dataOut_payload_0_4998 ? _zz_dataOut_payload_0_3058 : _zz_dataOut_payload_0_3069);
  assign _zz_dataOut_payload_0_5000 = (_zz_dataOut_payload_0_4998 ? _zz_dataOut_payload_0_3069 : _zz_dataOut_payload_0_3058);
  assign _zz_dataOut_payload_0_5001 = (_zz_dataOut_payload_0_3059 < _zz_dataOut_payload_0_3068);
  assign _zz_dataOut_payload_0_5002 = (_zz_dataOut_payload_0_5001 ? _zz_dataOut_payload_0_3059 : _zz_dataOut_payload_0_3068);
  assign _zz_dataOut_payload_0_5003 = (_zz_dataOut_payload_0_5001 ? _zz_dataOut_payload_0_3068 : _zz_dataOut_payload_0_3059);
  assign _zz_dataOut_payload_0_5004 = (_zz_dataOut_payload_0_3060 < _zz_dataOut_payload_0_3067);
  assign _zz_dataOut_payload_0_5005 = (_zz_dataOut_payload_0_5004 ? _zz_dataOut_payload_0_3060 : _zz_dataOut_payload_0_3067);
  assign _zz_dataOut_payload_0_5006 = (_zz_dataOut_payload_0_5004 ? _zz_dataOut_payload_0_3067 : _zz_dataOut_payload_0_3060);
  assign _zz_dataOut_payload_0_5007 = (_zz_dataOut_payload_0_3061 < _zz_dataOut_payload_0_3066);
  assign _zz_dataOut_payload_0_5008 = (_zz_dataOut_payload_0_5007 ? _zz_dataOut_payload_0_3061 : _zz_dataOut_payload_0_3066);
  assign _zz_dataOut_payload_0_5009 = (_zz_dataOut_payload_0_5007 ? _zz_dataOut_payload_0_3066 : _zz_dataOut_payload_0_3061);
  assign _zz_dataOut_payload_0_5010 = (_zz_dataOut_payload_0_3062 < _zz_dataOut_payload_0_3065);
  assign _zz_dataOut_payload_0_5011 = (_zz_dataOut_payload_0_5010 ? _zz_dataOut_payload_0_3062 : _zz_dataOut_payload_0_3065);
  assign _zz_dataOut_payload_0_5012 = (_zz_dataOut_payload_0_5010 ? _zz_dataOut_payload_0_3065 : _zz_dataOut_payload_0_3062);
  assign _zz_dataOut_payload_0_5013 = (_zz_dataOut_payload_0_3063 < _zz_dataOut_payload_0_3064);
  assign _zz_dataOut_payload_0_5014 = (_zz_dataOut_payload_0_5013 ? _zz_dataOut_payload_0_3063 : _zz_dataOut_payload_0_3064);
  assign _zz_dataOut_payload_0_5015 = (_zz_dataOut_payload_0_5013 ? _zz_dataOut_payload_0_3064 : _zz_dataOut_payload_0_3063);
  assign _zz_dataOut_payload_0_5016 = (_zz_dataOut_payload_0_4993 < _zz_dataOut_payload_0_5005);
  assign _zz_dataOut_payload_0_5017 = (_zz_dataOut_payload_0_5016 ? _zz_dataOut_payload_0_4993 : _zz_dataOut_payload_0_5005);
  assign _zz_dataOut_payload_0_5018 = (_zz_dataOut_payload_0_5016 ? _zz_dataOut_payload_0_5005 : _zz_dataOut_payload_0_4993);
  assign _zz_dataOut_payload_0_5019 = (_zz_dataOut_payload_0_4996 < _zz_dataOut_payload_0_5008);
  assign _zz_dataOut_payload_0_5020 = (_zz_dataOut_payload_0_5019 ? _zz_dataOut_payload_0_4996 : _zz_dataOut_payload_0_5008);
  assign _zz_dataOut_payload_0_5021 = (_zz_dataOut_payload_0_5019 ? _zz_dataOut_payload_0_5008 : _zz_dataOut_payload_0_4996);
  assign _zz_dataOut_payload_0_5022 = (_zz_dataOut_payload_0_4999 < _zz_dataOut_payload_0_5011);
  assign _zz_dataOut_payload_0_5023 = (_zz_dataOut_payload_0_5022 ? _zz_dataOut_payload_0_4999 : _zz_dataOut_payload_0_5011);
  assign _zz_dataOut_payload_0_5024 = (_zz_dataOut_payload_0_5022 ? _zz_dataOut_payload_0_5011 : _zz_dataOut_payload_0_4999);
  assign _zz_dataOut_payload_0_5025 = (_zz_dataOut_payload_0_5002 < _zz_dataOut_payload_0_5014);
  assign _zz_dataOut_payload_0_5026 = (_zz_dataOut_payload_0_5025 ? _zz_dataOut_payload_0_5002 : _zz_dataOut_payload_0_5014);
  assign _zz_dataOut_payload_0_5027 = (_zz_dataOut_payload_0_5025 ? _zz_dataOut_payload_0_5014 : _zz_dataOut_payload_0_5002);
  assign _zz_dataOut_payload_0_5028 = (_zz_dataOut_payload_0_5017 < _zz_dataOut_payload_0_5023);
  assign _zz_dataOut_payload_0_5029 = (_zz_dataOut_payload_0_5028 ? _zz_dataOut_payload_0_5017 : _zz_dataOut_payload_0_5023);
  assign _zz_dataOut_payload_0_5030 = (_zz_dataOut_payload_0_5028 ? _zz_dataOut_payload_0_5023 : _zz_dataOut_payload_0_5017);
  assign _zz_dataOut_payload_0_5031 = (_zz_dataOut_payload_0_5020 < _zz_dataOut_payload_0_5026);
  assign _zz_dataOut_payload_0_5032 = (_zz_dataOut_payload_0_5031 ? _zz_dataOut_payload_0_5020 : _zz_dataOut_payload_0_5026);
  assign _zz_dataOut_payload_0_5033 = (_zz_dataOut_payload_0_5031 ? _zz_dataOut_payload_0_5026 : _zz_dataOut_payload_0_5020);
  assign _zz_dataOut_payload_0_5034 = (_zz_dataOut_payload_0_5029 < _zz_dataOut_payload_0_5032);
  assign _zz_dataOut_payload_0_5035 = (_zz_dataOut_payload_0_5030 < _zz_dataOut_payload_0_5033);
  assign _zz_dataOut_payload_0_5040 = (_zz_dataOut_payload_0_5018 < _zz_dataOut_payload_0_5024);
  assign _zz_dataOut_payload_0_5041 = (_zz_dataOut_payload_0_5040 ? _zz_dataOut_payload_0_5018 : _zz_dataOut_payload_0_5024);
  assign _zz_dataOut_payload_0_5042 = (_zz_dataOut_payload_0_5040 ? _zz_dataOut_payload_0_5024 : _zz_dataOut_payload_0_5018);
  assign _zz_dataOut_payload_0_5043 = (_zz_dataOut_payload_0_5021 < _zz_dataOut_payload_0_5027);
  assign _zz_dataOut_payload_0_5044 = (_zz_dataOut_payload_0_5043 ? _zz_dataOut_payload_0_5021 : _zz_dataOut_payload_0_5027);
  assign _zz_dataOut_payload_0_5045 = (_zz_dataOut_payload_0_5043 ? _zz_dataOut_payload_0_5027 : _zz_dataOut_payload_0_5021);
  assign _zz_dataOut_payload_0_5046 = (_zz_dataOut_payload_0_5041 < _zz_dataOut_payload_0_5044);
  assign _zz_dataOut_payload_0_5047 = (_zz_dataOut_payload_0_5042 < _zz_dataOut_payload_0_5045);
  assign _zz_dataOut_payload_0_5060 = (_zz_dataOut_payload_0_5015 < _zz_dataOut_payload_0_5003);
  assign _zz_dataOut_payload_0_5061 = (_zz_dataOut_payload_0_5060 ? _zz_dataOut_payload_0_5015 : _zz_dataOut_payload_0_5003);
  assign _zz_dataOut_payload_0_5062 = (_zz_dataOut_payload_0_5060 ? _zz_dataOut_payload_0_5003 : _zz_dataOut_payload_0_5015);
  assign _zz_dataOut_payload_0_5063 = (_zz_dataOut_payload_0_5012 < _zz_dataOut_payload_0_5000);
  assign _zz_dataOut_payload_0_5064 = (_zz_dataOut_payload_0_5063 ? _zz_dataOut_payload_0_5012 : _zz_dataOut_payload_0_5000);
  assign _zz_dataOut_payload_0_5065 = (_zz_dataOut_payload_0_5063 ? _zz_dataOut_payload_0_5000 : _zz_dataOut_payload_0_5012);
  assign _zz_dataOut_payload_0_5066 = (_zz_dataOut_payload_0_5009 < _zz_dataOut_payload_0_4997);
  assign _zz_dataOut_payload_0_5067 = (_zz_dataOut_payload_0_5066 ? _zz_dataOut_payload_0_5009 : _zz_dataOut_payload_0_4997);
  assign _zz_dataOut_payload_0_5068 = (_zz_dataOut_payload_0_5066 ? _zz_dataOut_payload_0_4997 : _zz_dataOut_payload_0_5009);
  assign _zz_dataOut_payload_0_5069 = (_zz_dataOut_payload_0_5006 < _zz_dataOut_payload_0_4994);
  assign _zz_dataOut_payload_0_5070 = (_zz_dataOut_payload_0_5069 ? _zz_dataOut_payload_0_5006 : _zz_dataOut_payload_0_4994);
  assign _zz_dataOut_payload_0_5071 = (_zz_dataOut_payload_0_5069 ? _zz_dataOut_payload_0_4994 : _zz_dataOut_payload_0_5006);
  assign _zz_dataOut_payload_0_5072 = (_zz_dataOut_payload_0_5061 < _zz_dataOut_payload_0_5067);
  assign _zz_dataOut_payload_0_5073 = (_zz_dataOut_payload_0_5072 ? _zz_dataOut_payload_0_5061 : _zz_dataOut_payload_0_5067);
  assign _zz_dataOut_payload_0_5074 = (_zz_dataOut_payload_0_5072 ? _zz_dataOut_payload_0_5067 : _zz_dataOut_payload_0_5061);
  assign _zz_dataOut_payload_0_5075 = (_zz_dataOut_payload_0_5064 < _zz_dataOut_payload_0_5070);
  assign _zz_dataOut_payload_0_5076 = (_zz_dataOut_payload_0_5075 ? _zz_dataOut_payload_0_5064 : _zz_dataOut_payload_0_5070);
  assign _zz_dataOut_payload_0_5077 = (_zz_dataOut_payload_0_5075 ? _zz_dataOut_payload_0_5070 : _zz_dataOut_payload_0_5064);
  assign _zz_dataOut_payload_0_5078 = (_zz_dataOut_payload_0_5073 < _zz_dataOut_payload_0_5076);
  assign _zz_dataOut_payload_0_5079 = (_zz_dataOut_payload_0_5074 < _zz_dataOut_payload_0_5077);
  assign _zz_dataOut_payload_0_5084 = (_zz_dataOut_payload_0_5062 < _zz_dataOut_payload_0_5068);
  assign _zz_dataOut_payload_0_5085 = (_zz_dataOut_payload_0_5084 ? _zz_dataOut_payload_0_5062 : _zz_dataOut_payload_0_5068);
  assign _zz_dataOut_payload_0_5086 = (_zz_dataOut_payload_0_5084 ? _zz_dataOut_payload_0_5068 : _zz_dataOut_payload_0_5062);
  assign _zz_dataOut_payload_0_5087 = (_zz_dataOut_payload_0_5065 < _zz_dataOut_payload_0_5071);
  assign _zz_dataOut_payload_0_5088 = (_zz_dataOut_payload_0_5087 ? _zz_dataOut_payload_0_5065 : _zz_dataOut_payload_0_5071);
  assign _zz_dataOut_payload_0_5089 = (_zz_dataOut_payload_0_5087 ? _zz_dataOut_payload_0_5071 : _zz_dataOut_payload_0_5065);
  assign _zz_dataOut_payload_0_5090 = (_zz_dataOut_payload_0_5085 < _zz_dataOut_payload_0_5088);
  assign _zz_dataOut_payload_0_5091 = (_zz_dataOut_payload_0_5086 < _zz_dataOut_payload_0_5089);
  assign _zz_dataOut_payload_0_5376 = (_zz_dataOut_payload_0_5120 < _zz_dataOut_payload_0_5151);
  assign _zz_dataOut_payload_0_5377 = (_zz_dataOut_payload_0_5376 ? _zz_dataOut_payload_0_5120 : _zz_dataOut_payload_0_5151);
  assign _zz_dataOut_payload_0_5378 = (_zz_dataOut_payload_0_5376 ? _zz_dataOut_payload_0_5151 : _zz_dataOut_payload_0_5120);
  assign _zz_dataOut_payload_0_5379 = (_zz_dataOut_payload_0_5121 < _zz_dataOut_payload_0_5150);
  assign _zz_dataOut_payload_0_5380 = (_zz_dataOut_payload_0_5379 ? _zz_dataOut_payload_0_5121 : _zz_dataOut_payload_0_5150);
  assign _zz_dataOut_payload_0_5381 = (_zz_dataOut_payload_0_5379 ? _zz_dataOut_payload_0_5150 : _zz_dataOut_payload_0_5121);
  assign _zz_dataOut_payload_0_5382 = (_zz_dataOut_payload_0_5122 < _zz_dataOut_payload_0_5149);
  assign _zz_dataOut_payload_0_5383 = (_zz_dataOut_payload_0_5382 ? _zz_dataOut_payload_0_5122 : _zz_dataOut_payload_0_5149);
  assign _zz_dataOut_payload_0_5384 = (_zz_dataOut_payload_0_5382 ? _zz_dataOut_payload_0_5149 : _zz_dataOut_payload_0_5122);
  assign _zz_dataOut_payload_0_5385 = (_zz_dataOut_payload_0_5123 < _zz_dataOut_payload_0_5148);
  assign _zz_dataOut_payload_0_5386 = (_zz_dataOut_payload_0_5385 ? _zz_dataOut_payload_0_5123 : _zz_dataOut_payload_0_5148);
  assign _zz_dataOut_payload_0_5387 = (_zz_dataOut_payload_0_5385 ? _zz_dataOut_payload_0_5148 : _zz_dataOut_payload_0_5123);
  assign _zz_dataOut_payload_0_5388 = (_zz_dataOut_payload_0_5124 < _zz_dataOut_payload_0_5147);
  assign _zz_dataOut_payload_0_5389 = (_zz_dataOut_payload_0_5388 ? _zz_dataOut_payload_0_5124 : _zz_dataOut_payload_0_5147);
  assign _zz_dataOut_payload_0_5390 = (_zz_dataOut_payload_0_5388 ? _zz_dataOut_payload_0_5147 : _zz_dataOut_payload_0_5124);
  assign _zz_dataOut_payload_0_5391 = (_zz_dataOut_payload_0_5125 < _zz_dataOut_payload_0_5146);
  assign _zz_dataOut_payload_0_5392 = (_zz_dataOut_payload_0_5391 ? _zz_dataOut_payload_0_5125 : _zz_dataOut_payload_0_5146);
  assign _zz_dataOut_payload_0_5393 = (_zz_dataOut_payload_0_5391 ? _zz_dataOut_payload_0_5146 : _zz_dataOut_payload_0_5125);
  assign _zz_dataOut_payload_0_5394 = (_zz_dataOut_payload_0_5126 < _zz_dataOut_payload_0_5145);
  assign _zz_dataOut_payload_0_5395 = (_zz_dataOut_payload_0_5394 ? _zz_dataOut_payload_0_5126 : _zz_dataOut_payload_0_5145);
  assign _zz_dataOut_payload_0_5396 = (_zz_dataOut_payload_0_5394 ? _zz_dataOut_payload_0_5145 : _zz_dataOut_payload_0_5126);
  assign _zz_dataOut_payload_0_5397 = (_zz_dataOut_payload_0_5127 < _zz_dataOut_payload_0_5144);
  assign _zz_dataOut_payload_0_5398 = (_zz_dataOut_payload_0_5397 ? _zz_dataOut_payload_0_5127 : _zz_dataOut_payload_0_5144);
  assign _zz_dataOut_payload_0_5399 = (_zz_dataOut_payload_0_5397 ? _zz_dataOut_payload_0_5144 : _zz_dataOut_payload_0_5127);
  assign _zz_dataOut_payload_0_5400 = (_zz_dataOut_payload_0_5128 < _zz_dataOut_payload_0_5143);
  assign _zz_dataOut_payload_0_5401 = (_zz_dataOut_payload_0_5400 ? _zz_dataOut_payload_0_5128 : _zz_dataOut_payload_0_5143);
  assign _zz_dataOut_payload_0_5402 = (_zz_dataOut_payload_0_5400 ? _zz_dataOut_payload_0_5143 : _zz_dataOut_payload_0_5128);
  assign _zz_dataOut_payload_0_5403 = (_zz_dataOut_payload_0_5129 < _zz_dataOut_payload_0_5142);
  assign _zz_dataOut_payload_0_5404 = (_zz_dataOut_payload_0_5403 ? _zz_dataOut_payload_0_5129 : _zz_dataOut_payload_0_5142);
  assign _zz_dataOut_payload_0_5405 = (_zz_dataOut_payload_0_5403 ? _zz_dataOut_payload_0_5142 : _zz_dataOut_payload_0_5129);
  assign _zz_dataOut_payload_0_5406 = (_zz_dataOut_payload_0_5130 < _zz_dataOut_payload_0_5141);
  assign _zz_dataOut_payload_0_5407 = (_zz_dataOut_payload_0_5406 ? _zz_dataOut_payload_0_5130 : _zz_dataOut_payload_0_5141);
  assign _zz_dataOut_payload_0_5408 = (_zz_dataOut_payload_0_5406 ? _zz_dataOut_payload_0_5141 : _zz_dataOut_payload_0_5130);
  assign _zz_dataOut_payload_0_5409 = (_zz_dataOut_payload_0_5131 < _zz_dataOut_payload_0_5140);
  assign _zz_dataOut_payload_0_5410 = (_zz_dataOut_payload_0_5409 ? _zz_dataOut_payload_0_5131 : _zz_dataOut_payload_0_5140);
  assign _zz_dataOut_payload_0_5411 = (_zz_dataOut_payload_0_5409 ? _zz_dataOut_payload_0_5140 : _zz_dataOut_payload_0_5131);
  assign _zz_dataOut_payload_0_5412 = (_zz_dataOut_payload_0_5132 < _zz_dataOut_payload_0_5139);
  assign _zz_dataOut_payload_0_5413 = (_zz_dataOut_payload_0_5412 ? _zz_dataOut_payload_0_5132 : _zz_dataOut_payload_0_5139);
  assign _zz_dataOut_payload_0_5414 = (_zz_dataOut_payload_0_5412 ? _zz_dataOut_payload_0_5139 : _zz_dataOut_payload_0_5132);
  assign _zz_dataOut_payload_0_5415 = (_zz_dataOut_payload_0_5133 < _zz_dataOut_payload_0_5138);
  assign _zz_dataOut_payload_0_5416 = (_zz_dataOut_payload_0_5415 ? _zz_dataOut_payload_0_5133 : _zz_dataOut_payload_0_5138);
  assign _zz_dataOut_payload_0_5417 = (_zz_dataOut_payload_0_5415 ? _zz_dataOut_payload_0_5138 : _zz_dataOut_payload_0_5133);
  assign _zz_dataOut_payload_0_5418 = (_zz_dataOut_payload_0_5134 < _zz_dataOut_payload_0_5137);
  assign _zz_dataOut_payload_0_5419 = (_zz_dataOut_payload_0_5418 ? _zz_dataOut_payload_0_5134 : _zz_dataOut_payload_0_5137);
  assign _zz_dataOut_payload_0_5420 = (_zz_dataOut_payload_0_5418 ? _zz_dataOut_payload_0_5137 : _zz_dataOut_payload_0_5134);
  assign _zz_dataOut_payload_0_5421 = (_zz_dataOut_payload_0_5135 < _zz_dataOut_payload_0_5136);
  assign _zz_dataOut_payload_0_5422 = (_zz_dataOut_payload_0_5421 ? _zz_dataOut_payload_0_5135 : _zz_dataOut_payload_0_5136);
  assign _zz_dataOut_payload_0_5423 = (_zz_dataOut_payload_0_5421 ? _zz_dataOut_payload_0_5136 : _zz_dataOut_payload_0_5135);
  assign _zz_dataOut_payload_0_5424 = (_zz_dataOut_payload_0_5377 < _zz_dataOut_payload_0_5401);
  assign _zz_dataOut_payload_0_5425 = (_zz_dataOut_payload_0_5424 ? _zz_dataOut_payload_0_5377 : _zz_dataOut_payload_0_5401);
  assign _zz_dataOut_payload_0_5426 = (_zz_dataOut_payload_0_5424 ? _zz_dataOut_payload_0_5401 : _zz_dataOut_payload_0_5377);
  assign _zz_dataOut_payload_0_5427 = (_zz_dataOut_payload_0_5380 < _zz_dataOut_payload_0_5404);
  assign _zz_dataOut_payload_0_5428 = (_zz_dataOut_payload_0_5427 ? _zz_dataOut_payload_0_5380 : _zz_dataOut_payload_0_5404);
  assign _zz_dataOut_payload_0_5429 = (_zz_dataOut_payload_0_5427 ? _zz_dataOut_payload_0_5404 : _zz_dataOut_payload_0_5380);
  assign _zz_dataOut_payload_0_5430 = (_zz_dataOut_payload_0_5383 < _zz_dataOut_payload_0_5407);
  assign _zz_dataOut_payload_0_5431 = (_zz_dataOut_payload_0_5430 ? _zz_dataOut_payload_0_5383 : _zz_dataOut_payload_0_5407);
  assign _zz_dataOut_payload_0_5432 = (_zz_dataOut_payload_0_5430 ? _zz_dataOut_payload_0_5407 : _zz_dataOut_payload_0_5383);
  assign _zz_dataOut_payload_0_5433 = (_zz_dataOut_payload_0_5386 < _zz_dataOut_payload_0_5410);
  assign _zz_dataOut_payload_0_5434 = (_zz_dataOut_payload_0_5433 ? _zz_dataOut_payload_0_5386 : _zz_dataOut_payload_0_5410);
  assign _zz_dataOut_payload_0_5435 = (_zz_dataOut_payload_0_5433 ? _zz_dataOut_payload_0_5410 : _zz_dataOut_payload_0_5386);
  assign _zz_dataOut_payload_0_5436 = (_zz_dataOut_payload_0_5389 < _zz_dataOut_payload_0_5413);
  assign _zz_dataOut_payload_0_5437 = (_zz_dataOut_payload_0_5436 ? _zz_dataOut_payload_0_5389 : _zz_dataOut_payload_0_5413);
  assign _zz_dataOut_payload_0_5438 = (_zz_dataOut_payload_0_5436 ? _zz_dataOut_payload_0_5413 : _zz_dataOut_payload_0_5389);
  assign _zz_dataOut_payload_0_5439 = (_zz_dataOut_payload_0_5392 < _zz_dataOut_payload_0_5416);
  assign _zz_dataOut_payload_0_5440 = (_zz_dataOut_payload_0_5439 ? _zz_dataOut_payload_0_5392 : _zz_dataOut_payload_0_5416);
  assign _zz_dataOut_payload_0_5441 = (_zz_dataOut_payload_0_5439 ? _zz_dataOut_payload_0_5416 : _zz_dataOut_payload_0_5392);
  assign _zz_dataOut_payload_0_5442 = (_zz_dataOut_payload_0_5395 < _zz_dataOut_payload_0_5419);
  assign _zz_dataOut_payload_0_5443 = (_zz_dataOut_payload_0_5442 ? _zz_dataOut_payload_0_5395 : _zz_dataOut_payload_0_5419);
  assign _zz_dataOut_payload_0_5444 = (_zz_dataOut_payload_0_5442 ? _zz_dataOut_payload_0_5419 : _zz_dataOut_payload_0_5395);
  assign _zz_dataOut_payload_0_5445 = (_zz_dataOut_payload_0_5398 < _zz_dataOut_payload_0_5422);
  assign _zz_dataOut_payload_0_5446 = (_zz_dataOut_payload_0_5445 ? _zz_dataOut_payload_0_5398 : _zz_dataOut_payload_0_5422);
  assign _zz_dataOut_payload_0_5447 = (_zz_dataOut_payload_0_5445 ? _zz_dataOut_payload_0_5422 : _zz_dataOut_payload_0_5398);
  assign _zz_dataOut_payload_0_5448 = (_zz_dataOut_payload_0_5425 < _zz_dataOut_payload_0_5437);
  assign _zz_dataOut_payload_0_5449 = (_zz_dataOut_payload_0_5448 ? _zz_dataOut_payload_0_5425 : _zz_dataOut_payload_0_5437);
  assign _zz_dataOut_payload_0_5450 = (_zz_dataOut_payload_0_5448 ? _zz_dataOut_payload_0_5437 : _zz_dataOut_payload_0_5425);
  assign _zz_dataOut_payload_0_5451 = (_zz_dataOut_payload_0_5428 < _zz_dataOut_payload_0_5440);
  assign _zz_dataOut_payload_0_5452 = (_zz_dataOut_payload_0_5451 ? _zz_dataOut_payload_0_5428 : _zz_dataOut_payload_0_5440);
  assign _zz_dataOut_payload_0_5453 = (_zz_dataOut_payload_0_5451 ? _zz_dataOut_payload_0_5440 : _zz_dataOut_payload_0_5428);
  assign _zz_dataOut_payload_0_5454 = (_zz_dataOut_payload_0_5431 < _zz_dataOut_payload_0_5443);
  assign _zz_dataOut_payload_0_5455 = (_zz_dataOut_payload_0_5454 ? _zz_dataOut_payload_0_5431 : _zz_dataOut_payload_0_5443);
  assign _zz_dataOut_payload_0_5456 = (_zz_dataOut_payload_0_5454 ? _zz_dataOut_payload_0_5443 : _zz_dataOut_payload_0_5431);
  assign _zz_dataOut_payload_0_5457 = (_zz_dataOut_payload_0_5434 < _zz_dataOut_payload_0_5446);
  assign _zz_dataOut_payload_0_5458 = (_zz_dataOut_payload_0_5457 ? _zz_dataOut_payload_0_5434 : _zz_dataOut_payload_0_5446);
  assign _zz_dataOut_payload_0_5459 = (_zz_dataOut_payload_0_5457 ? _zz_dataOut_payload_0_5446 : _zz_dataOut_payload_0_5434);
  assign _zz_dataOut_payload_0_5460 = (_zz_dataOut_payload_0_5449 < _zz_dataOut_payload_0_5455);
  assign _zz_dataOut_payload_0_5461 = (_zz_dataOut_payload_0_5460 ? _zz_dataOut_payload_0_5449 : _zz_dataOut_payload_0_5455);
  assign _zz_dataOut_payload_0_5462 = (_zz_dataOut_payload_0_5460 ? _zz_dataOut_payload_0_5455 : _zz_dataOut_payload_0_5449);
  assign _zz_dataOut_payload_0_5463 = (_zz_dataOut_payload_0_5452 < _zz_dataOut_payload_0_5458);
  assign _zz_dataOut_payload_0_5464 = (_zz_dataOut_payload_0_5463 ? _zz_dataOut_payload_0_5452 : _zz_dataOut_payload_0_5458);
  assign _zz_dataOut_payload_0_5465 = (_zz_dataOut_payload_0_5463 ? _zz_dataOut_payload_0_5458 : _zz_dataOut_payload_0_5452);
  assign _zz_dataOut_payload_0_5466 = (_zz_dataOut_payload_0_5461 < _zz_dataOut_payload_0_5464);
  assign _zz_dataOut_payload_0_5467 = (_zz_dataOut_payload_0_5462 < _zz_dataOut_payload_0_5465);
  assign _zz_dataOut_payload_0_5472 = (_zz_dataOut_payload_0_5450 < _zz_dataOut_payload_0_5456);
  assign _zz_dataOut_payload_0_5473 = (_zz_dataOut_payload_0_5472 ? _zz_dataOut_payload_0_5450 : _zz_dataOut_payload_0_5456);
  assign _zz_dataOut_payload_0_5474 = (_zz_dataOut_payload_0_5472 ? _zz_dataOut_payload_0_5456 : _zz_dataOut_payload_0_5450);
  assign _zz_dataOut_payload_0_5475 = (_zz_dataOut_payload_0_5453 < _zz_dataOut_payload_0_5459);
  assign _zz_dataOut_payload_0_5476 = (_zz_dataOut_payload_0_5475 ? _zz_dataOut_payload_0_5453 : _zz_dataOut_payload_0_5459);
  assign _zz_dataOut_payload_0_5477 = (_zz_dataOut_payload_0_5475 ? _zz_dataOut_payload_0_5459 : _zz_dataOut_payload_0_5453);
  assign _zz_dataOut_payload_0_5478 = (_zz_dataOut_payload_0_5473 < _zz_dataOut_payload_0_5476);
  assign _zz_dataOut_payload_0_5479 = (_zz_dataOut_payload_0_5474 < _zz_dataOut_payload_0_5477);
  assign _zz_dataOut_payload_0_5492 = (_zz_dataOut_payload_0_5426 < _zz_dataOut_payload_0_5438);
  assign _zz_dataOut_payload_0_5493 = (_zz_dataOut_payload_0_5492 ? _zz_dataOut_payload_0_5426 : _zz_dataOut_payload_0_5438);
  assign _zz_dataOut_payload_0_5494 = (_zz_dataOut_payload_0_5492 ? _zz_dataOut_payload_0_5438 : _zz_dataOut_payload_0_5426);
  assign _zz_dataOut_payload_0_5495 = (_zz_dataOut_payload_0_5429 < _zz_dataOut_payload_0_5441);
  assign _zz_dataOut_payload_0_5496 = (_zz_dataOut_payload_0_5495 ? _zz_dataOut_payload_0_5429 : _zz_dataOut_payload_0_5441);
  assign _zz_dataOut_payload_0_5497 = (_zz_dataOut_payload_0_5495 ? _zz_dataOut_payload_0_5441 : _zz_dataOut_payload_0_5429);
  assign _zz_dataOut_payload_0_5498 = (_zz_dataOut_payload_0_5432 < _zz_dataOut_payload_0_5444);
  assign _zz_dataOut_payload_0_5499 = (_zz_dataOut_payload_0_5498 ? _zz_dataOut_payload_0_5432 : _zz_dataOut_payload_0_5444);
  assign _zz_dataOut_payload_0_5500 = (_zz_dataOut_payload_0_5498 ? _zz_dataOut_payload_0_5444 : _zz_dataOut_payload_0_5432);
  assign _zz_dataOut_payload_0_5501 = (_zz_dataOut_payload_0_5435 < _zz_dataOut_payload_0_5447);
  assign _zz_dataOut_payload_0_5502 = (_zz_dataOut_payload_0_5501 ? _zz_dataOut_payload_0_5435 : _zz_dataOut_payload_0_5447);
  assign _zz_dataOut_payload_0_5503 = (_zz_dataOut_payload_0_5501 ? _zz_dataOut_payload_0_5447 : _zz_dataOut_payload_0_5435);
  assign _zz_dataOut_payload_0_5504 = (_zz_dataOut_payload_0_5493 < _zz_dataOut_payload_0_5499);
  assign _zz_dataOut_payload_0_5505 = (_zz_dataOut_payload_0_5504 ? _zz_dataOut_payload_0_5493 : _zz_dataOut_payload_0_5499);
  assign _zz_dataOut_payload_0_5506 = (_zz_dataOut_payload_0_5504 ? _zz_dataOut_payload_0_5499 : _zz_dataOut_payload_0_5493);
  assign _zz_dataOut_payload_0_5507 = (_zz_dataOut_payload_0_5496 < _zz_dataOut_payload_0_5502);
  assign _zz_dataOut_payload_0_5508 = (_zz_dataOut_payload_0_5507 ? _zz_dataOut_payload_0_5496 : _zz_dataOut_payload_0_5502);
  assign _zz_dataOut_payload_0_5509 = (_zz_dataOut_payload_0_5507 ? _zz_dataOut_payload_0_5502 : _zz_dataOut_payload_0_5496);
  assign _zz_dataOut_payload_0_5510 = (_zz_dataOut_payload_0_5505 < _zz_dataOut_payload_0_5508);
  assign _zz_dataOut_payload_0_5511 = (_zz_dataOut_payload_0_5506 < _zz_dataOut_payload_0_5509);
  assign _zz_dataOut_payload_0_5516 = (_zz_dataOut_payload_0_5494 < _zz_dataOut_payload_0_5500);
  assign _zz_dataOut_payload_0_5517 = (_zz_dataOut_payload_0_5516 ? _zz_dataOut_payload_0_5494 : _zz_dataOut_payload_0_5500);
  assign _zz_dataOut_payload_0_5518 = (_zz_dataOut_payload_0_5516 ? _zz_dataOut_payload_0_5500 : _zz_dataOut_payload_0_5494);
  assign _zz_dataOut_payload_0_5519 = (_zz_dataOut_payload_0_5497 < _zz_dataOut_payload_0_5503);
  assign _zz_dataOut_payload_0_5520 = (_zz_dataOut_payload_0_5519 ? _zz_dataOut_payload_0_5497 : _zz_dataOut_payload_0_5503);
  assign _zz_dataOut_payload_0_5521 = (_zz_dataOut_payload_0_5519 ? _zz_dataOut_payload_0_5503 : _zz_dataOut_payload_0_5497);
  assign _zz_dataOut_payload_0_5522 = (_zz_dataOut_payload_0_5517 < _zz_dataOut_payload_0_5520);
  assign _zz_dataOut_payload_0_5523 = (_zz_dataOut_payload_0_5518 < _zz_dataOut_payload_0_5521);
  assign _zz_dataOut_payload_0_5552 = (_zz_dataOut_payload_0_5423 < _zz_dataOut_payload_0_5399);
  assign _zz_dataOut_payload_0_5553 = (_zz_dataOut_payload_0_5552 ? _zz_dataOut_payload_0_5423 : _zz_dataOut_payload_0_5399);
  assign _zz_dataOut_payload_0_5554 = (_zz_dataOut_payload_0_5552 ? _zz_dataOut_payload_0_5399 : _zz_dataOut_payload_0_5423);
  assign _zz_dataOut_payload_0_5555 = (_zz_dataOut_payload_0_5420 < _zz_dataOut_payload_0_5396);
  assign _zz_dataOut_payload_0_5556 = (_zz_dataOut_payload_0_5555 ? _zz_dataOut_payload_0_5420 : _zz_dataOut_payload_0_5396);
  assign _zz_dataOut_payload_0_5557 = (_zz_dataOut_payload_0_5555 ? _zz_dataOut_payload_0_5396 : _zz_dataOut_payload_0_5420);
  assign _zz_dataOut_payload_0_5558 = (_zz_dataOut_payload_0_5417 < _zz_dataOut_payload_0_5393);
  assign _zz_dataOut_payload_0_5559 = (_zz_dataOut_payload_0_5558 ? _zz_dataOut_payload_0_5417 : _zz_dataOut_payload_0_5393);
  assign _zz_dataOut_payload_0_5560 = (_zz_dataOut_payload_0_5558 ? _zz_dataOut_payload_0_5393 : _zz_dataOut_payload_0_5417);
  assign _zz_dataOut_payload_0_5561 = (_zz_dataOut_payload_0_5414 < _zz_dataOut_payload_0_5390);
  assign _zz_dataOut_payload_0_5562 = (_zz_dataOut_payload_0_5561 ? _zz_dataOut_payload_0_5414 : _zz_dataOut_payload_0_5390);
  assign _zz_dataOut_payload_0_5563 = (_zz_dataOut_payload_0_5561 ? _zz_dataOut_payload_0_5390 : _zz_dataOut_payload_0_5414);
  assign _zz_dataOut_payload_0_5564 = (_zz_dataOut_payload_0_5411 < _zz_dataOut_payload_0_5387);
  assign _zz_dataOut_payload_0_5565 = (_zz_dataOut_payload_0_5564 ? _zz_dataOut_payload_0_5411 : _zz_dataOut_payload_0_5387);
  assign _zz_dataOut_payload_0_5566 = (_zz_dataOut_payload_0_5564 ? _zz_dataOut_payload_0_5387 : _zz_dataOut_payload_0_5411);
  assign _zz_dataOut_payload_0_5567 = (_zz_dataOut_payload_0_5408 < _zz_dataOut_payload_0_5384);
  assign _zz_dataOut_payload_0_5568 = (_zz_dataOut_payload_0_5567 ? _zz_dataOut_payload_0_5408 : _zz_dataOut_payload_0_5384);
  assign _zz_dataOut_payload_0_5569 = (_zz_dataOut_payload_0_5567 ? _zz_dataOut_payload_0_5384 : _zz_dataOut_payload_0_5408);
  assign _zz_dataOut_payload_0_5570 = (_zz_dataOut_payload_0_5405 < _zz_dataOut_payload_0_5381);
  assign _zz_dataOut_payload_0_5571 = (_zz_dataOut_payload_0_5570 ? _zz_dataOut_payload_0_5405 : _zz_dataOut_payload_0_5381);
  assign _zz_dataOut_payload_0_5572 = (_zz_dataOut_payload_0_5570 ? _zz_dataOut_payload_0_5381 : _zz_dataOut_payload_0_5405);
  assign _zz_dataOut_payload_0_5573 = (_zz_dataOut_payload_0_5402 < _zz_dataOut_payload_0_5378);
  assign _zz_dataOut_payload_0_5574 = (_zz_dataOut_payload_0_5573 ? _zz_dataOut_payload_0_5402 : _zz_dataOut_payload_0_5378);
  assign _zz_dataOut_payload_0_5575 = (_zz_dataOut_payload_0_5573 ? _zz_dataOut_payload_0_5378 : _zz_dataOut_payload_0_5402);
  assign _zz_dataOut_payload_0_5576 = (_zz_dataOut_payload_0_5553 < _zz_dataOut_payload_0_5565);
  assign _zz_dataOut_payload_0_5577 = (_zz_dataOut_payload_0_5576 ? _zz_dataOut_payload_0_5553 : _zz_dataOut_payload_0_5565);
  assign _zz_dataOut_payload_0_5578 = (_zz_dataOut_payload_0_5576 ? _zz_dataOut_payload_0_5565 : _zz_dataOut_payload_0_5553);
  assign _zz_dataOut_payload_0_5579 = (_zz_dataOut_payload_0_5556 < _zz_dataOut_payload_0_5568);
  assign _zz_dataOut_payload_0_5580 = (_zz_dataOut_payload_0_5579 ? _zz_dataOut_payload_0_5556 : _zz_dataOut_payload_0_5568);
  assign _zz_dataOut_payload_0_5581 = (_zz_dataOut_payload_0_5579 ? _zz_dataOut_payload_0_5568 : _zz_dataOut_payload_0_5556);
  assign _zz_dataOut_payload_0_5582 = (_zz_dataOut_payload_0_5559 < _zz_dataOut_payload_0_5571);
  assign _zz_dataOut_payload_0_5583 = (_zz_dataOut_payload_0_5582 ? _zz_dataOut_payload_0_5559 : _zz_dataOut_payload_0_5571);
  assign _zz_dataOut_payload_0_5584 = (_zz_dataOut_payload_0_5582 ? _zz_dataOut_payload_0_5571 : _zz_dataOut_payload_0_5559);
  assign _zz_dataOut_payload_0_5585 = (_zz_dataOut_payload_0_5562 < _zz_dataOut_payload_0_5574);
  assign _zz_dataOut_payload_0_5586 = (_zz_dataOut_payload_0_5585 ? _zz_dataOut_payload_0_5562 : _zz_dataOut_payload_0_5574);
  assign _zz_dataOut_payload_0_5587 = (_zz_dataOut_payload_0_5585 ? _zz_dataOut_payload_0_5574 : _zz_dataOut_payload_0_5562);
  assign _zz_dataOut_payload_0_5588 = (_zz_dataOut_payload_0_5577 < _zz_dataOut_payload_0_5583);
  assign _zz_dataOut_payload_0_5589 = (_zz_dataOut_payload_0_5588 ? _zz_dataOut_payload_0_5577 : _zz_dataOut_payload_0_5583);
  assign _zz_dataOut_payload_0_5590 = (_zz_dataOut_payload_0_5588 ? _zz_dataOut_payload_0_5583 : _zz_dataOut_payload_0_5577);
  assign _zz_dataOut_payload_0_5591 = (_zz_dataOut_payload_0_5580 < _zz_dataOut_payload_0_5586);
  assign _zz_dataOut_payload_0_5592 = (_zz_dataOut_payload_0_5591 ? _zz_dataOut_payload_0_5580 : _zz_dataOut_payload_0_5586);
  assign _zz_dataOut_payload_0_5593 = (_zz_dataOut_payload_0_5591 ? _zz_dataOut_payload_0_5586 : _zz_dataOut_payload_0_5580);
  assign _zz_dataOut_payload_0_5594 = (_zz_dataOut_payload_0_5589 < _zz_dataOut_payload_0_5592);
  assign _zz_dataOut_payload_0_5595 = (_zz_dataOut_payload_0_5590 < _zz_dataOut_payload_0_5593);
  assign _zz_dataOut_payload_0_5600 = (_zz_dataOut_payload_0_5578 < _zz_dataOut_payload_0_5584);
  assign _zz_dataOut_payload_0_5601 = (_zz_dataOut_payload_0_5600 ? _zz_dataOut_payload_0_5578 : _zz_dataOut_payload_0_5584);
  assign _zz_dataOut_payload_0_5602 = (_zz_dataOut_payload_0_5600 ? _zz_dataOut_payload_0_5584 : _zz_dataOut_payload_0_5578);
  assign _zz_dataOut_payload_0_5603 = (_zz_dataOut_payload_0_5581 < _zz_dataOut_payload_0_5587);
  assign _zz_dataOut_payload_0_5604 = (_zz_dataOut_payload_0_5603 ? _zz_dataOut_payload_0_5581 : _zz_dataOut_payload_0_5587);
  assign _zz_dataOut_payload_0_5605 = (_zz_dataOut_payload_0_5603 ? _zz_dataOut_payload_0_5587 : _zz_dataOut_payload_0_5581);
  assign _zz_dataOut_payload_0_5606 = (_zz_dataOut_payload_0_5601 < _zz_dataOut_payload_0_5604);
  assign _zz_dataOut_payload_0_5607 = (_zz_dataOut_payload_0_5602 < _zz_dataOut_payload_0_5605);
  assign _zz_dataOut_payload_0_5620 = (_zz_dataOut_payload_0_5554 < _zz_dataOut_payload_0_5566);
  assign _zz_dataOut_payload_0_5621 = (_zz_dataOut_payload_0_5620 ? _zz_dataOut_payload_0_5554 : _zz_dataOut_payload_0_5566);
  assign _zz_dataOut_payload_0_5622 = (_zz_dataOut_payload_0_5620 ? _zz_dataOut_payload_0_5566 : _zz_dataOut_payload_0_5554);
  assign _zz_dataOut_payload_0_5623 = (_zz_dataOut_payload_0_5557 < _zz_dataOut_payload_0_5569);
  assign _zz_dataOut_payload_0_5624 = (_zz_dataOut_payload_0_5623 ? _zz_dataOut_payload_0_5557 : _zz_dataOut_payload_0_5569);
  assign _zz_dataOut_payload_0_5625 = (_zz_dataOut_payload_0_5623 ? _zz_dataOut_payload_0_5569 : _zz_dataOut_payload_0_5557);
  assign _zz_dataOut_payload_0_5626 = (_zz_dataOut_payload_0_5560 < _zz_dataOut_payload_0_5572);
  assign _zz_dataOut_payload_0_5627 = (_zz_dataOut_payload_0_5626 ? _zz_dataOut_payload_0_5560 : _zz_dataOut_payload_0_5572);
  assign _zz_dataOut_payload_0_5628 = (_zz_dataOut_payload_0_5626 ? _zz_dataOut_payload_0_5572 : _zz_dataOut_payload_0_5560);
  assign _zz_dataOut_payload_0_5629 = (_zz_dataOut_payload_0_5563 < _zz_dataOut_payload_0_5575);
  assign _zz_dataOut_payload_0_5630 = (_zz_dataOut_payload_0_5629 ? _zz_dataOut_payload_0_5563 : _zz_dataOut_payload_0_5575);
  assign _zz_dataOut_payload_0_5631 = (_zz_dataOut_payload_0_5629 ? _zz_dataOut_payload_0_5575 : _zz_dataOut_payload_0_5563);
  assign _zz_dataOut_payload_0_5632 = (_zz_dataOut_payload_0_5621 < _zz_dataOut_payload_0_5627);
  assign _zz_dataOut_payload_0_5633 = (_zz_dataOut_payload_0_5632 ? _zz_dataOut_payload_0_5621 : _zz_dataOut_payload_0_5627);
  assign _zz_dataOut_payload_0_5634 = (_zz_dataOut_payload_0_5632 ? _zz_dataOut_payload_0_5627 : _zz_dataOut_payload_0_5621);
  assign _zz_dataOut_payload_0_5635 = (_zz_dataOut_payload_0_5624 < _zz_dataOut_payload_0_5630);
  assign _zz_dataOut_payload_0_5636 = (_zz_dataOut_payload_0_5635 ? _zz_dataOut_payload_0_5624 : _zz_dataOut_payload_0_5630);
  assign _zz_dataOut_payload_0_5637 = (_zz_dataOut_payload_0_5635 ? _zz_dataOut_payload_0_5630 : _zz_dataOut_payload_0_5624);
  assign _zz_dataOut_payload_0_5638 = (_zz_dataOut_payload_0_5633 < _zz_dataOut_payload_0_5636);
  assign _zz_dataOut_payload_0_5639 = (_zz_dataOut_payload_0_5634 < _zz_dataOut_payload_0_5637);
  assign _zz_dataOut_payload_0_5644 = (_zz_dataOut_payload_0_5622 < _zz_dataOut_payload_0_5628);
  assign _zz_dataOut_payload_0_5645 = (_zz_dataOut_payload_0_5644 ? _zz_dataOut_payload_0_5622 : _zz_dataOut_payload_0_5628);
  assign _zz_dataOut_payload_0_5646 = (_zz_dataOut_payload_0_5644 ? _zz_dataOut_payload_0_5628 : _zz_dataOut_payload_0_5622);
  assign _zz_dataOut_payload_0_5647 = (_zz_dataOut_payload_0_5625 < _zz_dataOut_payload_0_5631);
  assign _zz_dataOut_payload_0_5648 = (_zz_dataOut_payload_0_5647 ? _zz_dataOut_payload_0_5625 : _zz_dataOut_payload_0_5631);
  assign _zz_dataOut_payload_0_5649 = (_zz_dataOut_payload_0_5647 ? _zz_dataOut_payload_0_5631 : _zz_dataOut_payload_0_5625);
  assign _zz_dataOut_payload_0_5650 = (_zz_dataOut_payload_0_5645 < _zz_dataOut_payload_0_5648);
  assign _zz_dataOut_payload_0_5651 = (_zz_dataOut_payload_0_5646 < _zz_dataOut_payload_0_5649);
  assign _zz_dataOut_payload_0_5712 = (_zz_dataOut_payload_0_5152 < _zz_dataOut_payload_0_5183);
  assign _zz_dataOut_payload_0_5713 = (_zz_dataOut_payload_0_5712 ? _zz_dataOut_payload_0_5152 : _zz_dataOut_payload_0_5183);
  assign _zz_dataOut_payload_0_5714 = (_zz_dataOut_payload_0_5712 ? _zz_dataOut_payload_0_5183 : _zz_dataOut_payload_0_5152);
  assign _zz_dataOut_payload_0_5715 = (_zz_dataOut_payload_0_5153 < _zz_dataOut_payload_0_5182);
  assign _zz_dataOut_payload_0_5716 = (_zz_dataOut_payload_0_5715 ? _zz_dataOut_payload_0_5153 : _zz_dataOut_payload_0_5182);
  assign _zz_dataOut_payload_0_5717 = (_zz_dataOut_payload_0_5715 ? _zz_dataOut_payload_0_5182 : _zz_dataOut_payload_0_5153);
  assign _zz_dataOut_payload_0_5718 = (_zz_dataOut_payload_0_5154 < _zz_dataOut_payload_0_5181);
  assign _zz_dataOut_payload_0_5719 = (_zz_dataOut_payload_0_5718 ? _zz_dataOut_payload_0_5154 : _zz_dataOut_payload_0_5181);
  assign _zz_dataOut_payload_0_5720 = (_zz_dataOut_payload_0_5718 ? _zz_dataOut_payload_0_5181 : _zz_dataOut_payload_0_5154);
  assign _zz_dataOut_payload_0_5721 = (_zz_dataOut_payload_0_5155 < _zz_dataOut_payload_0_5180);
  assign _zz_dataOut_payload_0_5722 = (_zz_dataOut_payload_0_5721 ? _zz_dataOut_payload_0_5155 : _zz_dataOut_payload_0_5180);
  assign _zz_dataOut_payload_0_5723 = (_zz_dataOut_payload_0_5721 ? _zz_dataOut_payload_0_5180 : _zz_dataOut_payload_0_5155);
  assign _zz_dataOut_payload_0_5724 = (_zz_dataOut_payload_0_5156 < _zz_dataOut_payload_0_5179);
  assign _zz_dataOut_payload_0_5725 = (_zz_dataOut_payload_0_5724 ? _zz_dataOut_payload_0_5156 : _zz_dataOut_payload_0_5179);
  assign _zz_dataOut_payload_0_5726 = (_zz_dataOut_payload_0_5724 ? _zz_dataOut_payload_0_5179 : _zz_dataOut_payload_0_5156);
  assign _zz_dataOut_payload_0_5727 = (_zz_dataOut_payload_0_5157 < _zz_dataOut_payload_0_5178);
  assign _zz_dataOut_payload_0_5728 = (_zz_dataOut_payload_0_5727 ? _zz_dataOut_payload_0_5157 : _zz_dataOut_payload_0_5178);
  assign _zz_dataOut_payload_0_5729 = (_zz_dataOut_payload_0_5727 ? _zz_dataOut_payload_0_5178 : _zz_dataOut_payload_0_5157);
  assign _zz_dataOut_payload_0_5730 = (_zz_dataOut_payload_0_5158 < _zz_dataOut_payload_0_5177);
  assign _zz_dataOut_payload_0_5731 = (_zz_dataOut_payload_0_5730 ? _zz_dataOut_payload_0_5158 : _zz_dataOut_payload_0_5177);
  assign _zz_dataOut_payload_0_5732 = (_zz_dataOut_payload_0_5730 ? _zz_dataOut_payload_0_5177 : _zz_dataOut_payload_0_5158);
  assign _zz_dataOut_payload_0_5733 = (_zz_dataOut_payload_0_5159 < _zz_dataOut_payload_0_5176);
  assign _zz_dataOut_payload_0_5734 = (_zz_dataOut_payload_0_5733 ? _zz_dataOut_payload_0_5159 : _zz_dataOut_payload_0_5176);
  assign _zz_dataOut_payload_0_5735 = (_zz_dataOut_payload_0_5733 ? _zz_dataOut_payload_0_5176 : _zz_dataOut_payload_0_5159);
  assign _zz_dataOut_payload_0_5736 = (_zz_dataOut_payload_0_5160 < _zz_dataOut_payload_0_5175);
  assign _zz_dataOut_payload_0_5737 = (_zz_dataOut_payload_0_5736 ? _zz_dataOut_payload_0_5160 : _zz_dataOut_payload_0_5175);
  assign _zz_dataOut_payload_0_5738 = (_zz_dataOut_payload_0_5736 ? _zz_dataOut_payload_0_5175 : _zz_dataOut_payload_0_5160);
  assign _zz_dataOut_payload_0_5739 = (_zz_dataOut_payload_0_5161 < _zz_dataOut_payload_0_5174);
  assign _zz_dataOut_payload_0_5740 = (_zz_dataOut_payload_0_5739 ? _zz_dataOut_payload_0_5161 : _zz_dataOut_payload_0_5174);
  assign _zz_dataOut_payload_0_5741 = (_zz_dataOut_payload_0_5739 ? _zz_dataOut_payload_0_5174 : _zz_dataOut_payload_0_5161);
  assign _zz_dataOut_payload_0_5742 = (_zz_dataOut_payload_0_5162 < _zz_dataOut_payload_0_5173);
  assign _zz_dataOut_payload_0_5743 = (_zz_dataOut_payload_0_5742 ? _zz_dataOut_payload_0_5162 : _zz_dataOut_payload_0_5173);
  assign _zz_dataOut_payload_0_5744 = (_zz_dataOut_payload_0_5742 ? _zz_dataOut_payload_0_5173 : _zz_dataOut_payload_0_5162);
  assign _zz_dataOut_payload_0_5745 = (_zz_dataOut_payload_0_5163 < _zz_dataOut_payload_0_5172);
  assign _zz_dataOut_payload_0_5746 = (_zz_dataOut_payload_0_5745 ? _zz_dataOut_payload_0_5163 : _zz_dataOut_payload_0_5172);
  assign _zz_dataOut_payload_0_5747 = (_zz_dataOut_payload_0_5745 ? _zz_dataOut_payload_0_5172 : _zz_dataOut_payload_0_5163);
  assign _zz_dataOut_payload_0_5748 = (_zz_dataOut_payload_0_5164 < _zz_dataOut_payload_0_5171);
  assign _zz_dataOut_payload_0_5749 = (_zz_dataOut_payload_0_5748 ? _zz_dataOut_payload_0_5164 : _zz_dataOut_payload_0_5171);
  assign _zz_dataOut_payload_0_5750 = (_zz_dataOut_payload_0_5748 ? _zz_dataOut_payload_0_5171 : _zz_dataOut_payload_0_5164);
  assign _zz_dataOut_payload_0_5751 = (_zz_dataOut_payload_0_5165 < _zz_dataOut_payload_0_5170);
  assign _zz_dataOut_payload_0_5752 = (_zz_dataOut_payload_0_5751 ? _zz_dataOut_payload_0_5165 : _zz_dataOut_payload_0_5170);
  assign _zz_dataOut_payload_0_5753 = (_zz_dataOut_payload_0_5751 ? _zz_dataOut_payload_0_5170 : _zz_dataOut_payload_0_5165);
  assign _zz_dataOut_payload_0_5754 = (_zz_dataOut_payload_0_5166 < _zz_dataOut_payload_0_5169);
  assign _zz_dataOut_payload_0_5755 = (_zz_dataOut_payload_0_5754 ? _zz_dataOut_payload_0_5166 : _zz_dataOut_payload_0_5169);
  assign _zz_dataOut_payload_0_5756 = (_zz_dataOut_payload_0_5754 ? _zz_dataOut_payload_0_5169 : _zz_dataOut_payload_0_5166);
  assign _zz_dataOut_payload_0_5757 = (_zz_dataOut_payload_0_5167 < _zz_dataOut_payload_0_5168);
  assign _zz_dataOut_payload_0_5758 = (_zz_dataOut_payload_0_5757 ? _zz_dataOut_payload_0_5167 : _zz_dataOut_payload_0_5168);
  assign _zz_dataOut_payload_0_5759 = (_zz_dataOut_payload_0_5757 ? _zz_dataOut_payload_0_5168 : _zz_dataOut_payload_0_5167);
  assign _zz_dataOut_payload_0_5760 = (_zz_dataOut_payload_0_5713 < _zz_dataOut_payload_0_5737);
  assign _zz_dataOut_payload_0_5761 = (_zz_dataOut_payload_0_5760 ? _zz_dataOut_payload_0_5713 : _zz_dataOut_payload_0_5737);
  assign _zz_dataOut_payload_0_5762 = (_zz_dataOut_payload_0_5760 ? _zz_dataOut_payload_0_5737 : _zz_dataOut_payload_0_5713);
  assign _zz_dataOut_payload_0_5763 = (_zz_dataOut_payload_0_5716 < _zz_dataOut_payload_0_5740);
  assign _zz_dataOut_payload_0_5764 = (_zz_dataOut_payload_0_5763 ? _zz_dataOut_payload_0_5716 : _zz_dataOut_payload_0_5740);
  assign _zz_dataOut_payload_0_5765 = (_zz_dataOut_payload_0_5763 ? _zz_dataOut_payload_0_5740 : _zz_dataOut_payload_0_5716);
  assign _zz_dataOut_payload_0_5766 = (_zz_dataOut_payload_0_5719 < _zz_dataOut_payload_0_5743);
  assign _zz_dataOut_payload_0_5767 = (_zz_dataOut_payload_0_5766 ? _zz_dataOut_payload_0_5719 : _zz_dataOut_payload_0_5743);
  assign _zz_dataOut_payload_0_5768 = (_zz_dataOut_payload_0_5766 ? _zz_dataOut_payload_0_5743 : _zz_dataOut_payload_0_5719);
  assign _zz_dataOut_payload_0_5769 = (_zz_dataOut_payload_0_5722 < _zz_dataOut_payload_0_5746);
  assign _zz_dataOut_payload_0_5770 = (_zz_dataOut_payload_0_5769 ? _zz_dataOut_payload_0_5722 : _zz_dataOut_payload_0_5746);
  assign _zz_dataOut_payload_0_5771 = (_zz_dataOut_payload_0_5769 ? _zz_dataOut_payload_0_5746 : _zz_dataOut_payload_0_5722);
  assign _zz_dataOut_payload_0_5772 = (_zz_dataOut_payload_0_5725 < _zz_dataOut_payload_0_5749);
  assign _zz_dataOut_payload_0_5773 = (_zz_dataOut_payload_0_5772 ? _zz_dataOut_payload_0_5725 : _zz_dataOut_payload_0_5749);
  assign _zz_dataOut_payload_0_5774 = (_zz_dataOut_payload_0_5772 ? _zz_dataOut_payload_0_5749 : _zz_dataOut_payload_0_5725);
  assign _zz_dataOut_payload_0_5775 = (_zz_dataOut_payload_0_5728 < _zz_dataOut_payload_0_5752);
  assign _zz_dataOut_payload_0_5776 = (_zz_dataOut_payload_0_5775 ? _zz_dataOut_payload_0_5728 : _zz_dataOut_payload_0_5752);
  assign _zz_dataOut_payload_0_5777 = (_zz_dataOut_payload_0_5775 ? _zz_dataOut_payload_0_5752 : _zz_dataOut_payload_0_5728);
  assign _zz_dataOut_payload_0_5778 = (_zz_dataOut_payload_0_5731 < _zz_dataOut_payload_0_5755);
  assign _zz_dataOut_payload_0_5779 = (_zz_dataOut_payload_0_5778 ? _zz_dataOut_payload_0_5731 : _zz_dataOut_payload_0_5755);
  assign _zz_dataOut_payload_0_5780 = (_zz_dataOut_payload_0_5778 ? _zz_dataOut_payload_0_5755 : _zz_dataOut_payload_0_5731);
  assign _zz_dataOut_payload_0_5781 = (_zz_dataOut_payload_0_5734 < _zz_dataOut_payload_0_5758);
  assign _zz_dataOut_payload_0_5782 = (_zz_dataOut_payload_0_5781 ? _zz_dataOut_payload_0_5734 : _zz_dataOut_payload_0_5758);
  assign _zz_dataOut_payload_0_5783 = (_zz_dataOut_payload_0_5781 ? _zz_dataOut_payload_0_5758 : _zz_dataOut_payload_0_5734);
  assign _zz_dataOut_payload_0_5784 = (_zz_dataOut_payload_0_5761 < _zz_dataOut_payload_0_5773);
  assign _zz_dataOut_payload_0_5785 = (_zz_dataOut_payload_0_5784 ? _zz_dataOut_payload_0_5761 : _zz_dataOut_payload_0_5773);
  assign _zz_dataOut_payload_0_5786 = (_zz_dataOut_payload_0_5784 ? _zz_dataOut_payload_0_5773 : _zz_dataOut_payload_0_5761);
  assign _zz_dataOut_payload_0_5787 = (_zz_dataOut_payload_0_5764 < _zz_dataOut_payload_0_5776);
  assign _zz_dataOut_payload_0_5788 = (_zz_dataOut_payload_0_5787 ? _zz_dataOut_payload_0_5764 : _zz_dataOut_payload_0_5776);
  assign _zz_dataOut_payload_0_5789 = (_zz_dataOut_payload_0_5787 ? _zz_dataOut_payload_0_5776 : _zz_dataOut_payload_0_5764);
  assign _zz_dataOut_payload_0_5790 = (_zz_dataOut_payload_0_5767 < _zz_dataOut_payload_0_5779);
  assign _zz_dataOut_payload_0_5791 = (_zz_dataOut_payload_0_5790 ? _zz_dataOut_payload_0_5767 : _zz_dataOut_payload_0_5779);
  assign _zz_dataOut_payload_0_5792 = (_zz_dataOut_payload_0_5790 ? _zz_dataOut_payload_0_5779 : _zz_dataOut_payload_0_5767);
  assign _zz_dataOut_payload_0_5793 = (_zz_dataOut_payload_0_5770 < _zz_dataOut_payload_0_5782);
  assign _zz_dataOut_payload_0_5794 = (_zz_dataOut_payload_0_5793 ? _zz_dataOut_payload_0_5770 : _zz_dataOut_payload_0_5782);
  assign _zz_dataOut_payload_0_5795 = (_zz_dataOut_payload_0_5793 ? _zz_dataOut_payload_0_5782 : _zz_dataOut_payload_0_5770);
  assign _zz_dataOut_payload_0_5796 = (_zz_dataOut_payload_0_5785 < _zz_dataOut_payload_0_5791);
  assign _zz_dataOut_payload_0_5797 = (_zz_dataOut_payload_0_5796 ? _zz_dataOut_payload_0_5785 : _zz_dataOut_payload_0_5791);
  assign _zz_dataOut_payload_0_5798 = (_zz_dataOut_payload_0_5796 ? _zz_dataOut_payload_0_5791 : _zz_dataOut_payload_0_5785);
  assign _zz_dataOut_payload_0_5799 = (_zz_dataOut_payload_0_5788 < _zz_dataOut_payload_0_5794);
  assign _zz_dataOut_payload_0_5800 = (_zz_dataOut_payload_0_5799 ? _zz_dataOut_payload_0_5788 : _zz_dataOut_payload_0_5794);
  assign _zz_dataOut_payload_0_5801 = (_zz_dataOut_payload_0_5799 ? _zz_dataOut_payload_0_5794 : _zz_dataOut_payload_0_5788);
  assign _zz_dataOut_payload_0_5802 = (_zz_dataOut_payload_0_5797 < _zz_dataOut_payload_0_5800);
  assign _zz_dataOut_payload_0_5803 = (_zz_dataOut_payload_0_5798 < _zz_dataOut_payload_0_5801);
  assign _zz_dataOut_payload_0_5808 = (_zz_dataOut_payload_0_5786 < _zz_dataOut_payload_0_5792);
  assign _zz_dataOut_payload_0_5809 = (_zz_dataOut_payload_0_5808 ? _zz_dataOut_payload_0_5786 : _zz_dataOut_payload_0_5792);
  assign _zz_dataOut_payload_0_5810 = (_zz_dataOut_payload_0_5808 ? _zz_dataOut_payload_0_5792 : _zz_dataOut_payload_0_5786);
  assign _zz_dataOut_payload_0_5811 = (_zz_dataOut_payload_0_5789 < _zz_dataOut_payload_0_5795);
  assign _zz_dataOut_payload_0_5812 = (_zz_dataOut_payload_0_5811 ? _zz_dataOut_payload_0_5789 : _zz_dataOut_payload_0_5795);
  assign _zz_dataOut_payload_0_5813 = (_zz_dataOut_payload_0_5811 ? _zz_dataOut_payload_0_5795 : _zz_dataOut_payload_0_5789);
  assign _zz_dataOut_payload_0_5814 = (_zz_dataOut_payload_0_5809 < _zz_dataOut_payload_0_5812);
  assign _zz_dataOut_payload_0_5815 = (_zz_dataOut_payload_0_5810 < _zz_dataOut_payload_0_5813);
  assign _zz_dataOut_payload_0_5828 = (_zz_dataOut_payload_0_5762 < _zz_dataOut_payload_0_5774);
  assign _zz_dataOut_payload_0_5829 = (_zz_dataOut_payload_0_5828 ? _zz_dataOut_payload_0_5762 : _zz_dataOut_payload_0_5774);
  assign _zz_dataOut_payload_0_5830 = (_zz_dataOut_payload_0_5828 ? _zz_dataOut_payload_0_5774 : _zz_dataOut_payload_0_5762);
  assign _zz_dataOut_payload_0_5831 = (_zz_dataOut_payload_0_5765 < _zz_dataOut_payload_0_5777);
  assign _zz_dataOut_payload_0_5832 = (_zz_dataOut_payload_0_5831 ? _zz_dataOut_payload_0_5765 : _zz_dataOut_payload_0_5777);
  assign _zz_dataOut_payload_0_5833 = (_zz_dataOut_payload_0_5831 ? _zz_dataOut_payload_0_5777 : _zz_dataOut_payload_0_5765);
  assign _zz_dataOut_payload_0_5834 = (_zz_dataOut_payload_0_5768 < _zz_dataOut_payload_0_5780);
  assign _zz_dataOut_payload_0_5835 = (_zz_dataOut_payload_0_5834 ? _zz_dataOut_payload_0_5768 : _zz_dataOut_payload_0_5780);
  assign _zz_dataOut_payload_0_5836 = (_zz_dataOut_payload_0_5834 ? _zz_dataOut_payload_0_5780 : _zz_dataOut_payload_0_5768);
  assign _zz_dataOut_payload_0_5837 = (_zz_dataOut_payload_0_5771 < _zz_dataOut_payload_0_5783);
  assign _zz_dataOut_payload_0_5838 = (_zz_dataOut_payload_0_5837 ? _zz_dataOut_payload_0_5771 : _zz_dataOut_payload_0_5783);
  assign _zz_dataOut_payload_0_5839 = (_zz_dataOut_payload_0_5837 ? _zz_dataOut_payload_0_5783 : _zz_dataOut_payload_0_5771);
  assign _zz_dataOut_payload_0_5840 = (_zz_dataOut_payload_0_5829 < _zz_dataOut_payload_0_5835);
  assign _zz_dataOut_payload_0_5841 = (_zz_dataOut_payload_0_5840 ? _zz_dataOut_payload_0_5829 : _zz_dataOut_payload_0_5835);
  assign _zz_dataOut_payload_0_5842 = (_zz_dataOut_payload_0_5840 ? _zz_dataOut_payload_0_5835 : _zz_dataOut_payload_0_5829);
  assign _zz_dataOut_payload_0_5843 = (_zz_dataOut_payload_0_5832 < _zz_dataOut_payload_0_5838);
  assign _zz_dataOut_payload_0_5844 = (_zz_dataOut_payload_0_5843 ? _zz_dataOut_payload_0_5832 : _zz_dataOut_payload_0_5838);
  assign _zz_dataOut_payload_0_5845 = (_zz_dataOut_payload_0_5843 ? _zz_dataOut_payload_0_5838 : _zz_dataOut_payload_0_5832);
  assign _zz_dataOut_payload_0_5846 = (_zz_dataOut_payload_0_5841 < _zz_dataOut_payload_0_5844);
  assign _zz_dataOut_payload_0_5847 = (_zz_dataOut_payload_0_5842 < _zz_dataOut_payload_0_5845);
  assign _zz_dataOut_payload_0_5852 = (_zz_dataOut_payload_0_5830 < _zz_dataOut_payload_0_5836);
  assign _zz_dataOut_payload_0_5853 = (_zz_dataOut_payload_0_5852 ? _zz_dataOut_payload_0_5830 : _zz_dataOut_payload_0_5836);
  assign _zz_dataOut_payload_0_5854 = (_zz_dataOut_payload_0_5852 ? _zz_dataOut_payload_0_5836 : _zz_dataOut_payload_0_5830);
  assign _zz_dataOut_payload_0_5855 = (_zz_dataOut_payload_0_5833 < _zz_dataOut_payload_0_5839);
  assign _zz_dataOut_payload_0_5856 = (_zz_dataOut_payload_0_5855 ? _zz_dataOut_payload_0_5833 : _zz_dataOut_payload_0_5839);
  assign _zz_dataOut_payload_0_5857 = (_zz_dataOut_payload_0_5855 ? _zz_dataOut_payload_0_5839 : _zz_dataOut_payload_0_5833);
  assign _zz_dataOut_payload_0_5858 = (_zz_dataOut_payload_0_5853 < _zz_dataOut_payload_0_5856);
  assign _zz_dataOut_payload_0_5859 = (_zz_dataOut_payload_0_5854 < _zz_dataOut_payload_0_5857);
  assign _zz_dataOut_payload_0_5888 = (_zz_dataOut_payload_0_5759 < _zz_dataOut_payload_0_5735);
  assign _zz_dataOut_payload_0_5889 = (_zz_dataOut_payload_0_5888 ? _zz_dataOut_payload_0_5759 : _zz_dataOut_payload_0_5735);
  assign _zz_dataOut_payload_0_5890 = (_zz_dataOut_payload_0_5888 ? _zz_dataOut_payload_0_5735 : _zz_dataOut_payload_0_5759);
  assign _zz_dataOut_payload_0_5891 = (_zz_dataOut_payload_0_5756 < _zz_dataOut_payload_0_5732);
  assign _zz_dataOut_payload_0_5892 = (_zz_dataOut_payload_0_5891 ? _zz_dataOut_payload_0_5756 : _zz_dataOut_payload_0_5732);
  assign _zz_dataOut_payload_0_5893 = (_zz_dataOut_payload_0_5891 ? _zz_dataOut_payload_0_5732 : _zz_dataOut_payload_0_5756);
  assign _zz_dataOut_payload_0_5894 = (_zz_dataOut_payload_0_5753 < _zz_dataOut_payload_0_5729);
  assign _zz_dataOut_payload_0_5895 = (_zz_dataOut_payload_0_5894 ? _zz_dataOut_payload_0_5753 : _zz_dataOut_payload_0_5729);
  assign _zz_dataOut_payload_0_5896 = (_zz_dataOut_payload_0_5894 ? _zz_dataOut_payload_0_5729 : _zz_dataOut_payload_0_5753);
  assign _zz_dataOut_payload_0_5897 = (_zz_dataOut_payload_0_5750 < _zz_dataOut_payload_0_5726);
  assign _zz_dataOut_payload_0_5898 = (_zz_dataOut_payload_0_5897 ? _zz_dataOut_payload_0_5750 : _zz_dataOut_payload_0_5726);
  assign _zz_dataOut_payload_0_5899 = (_zz_dataOut_payload_0_5897 ? _zz_dataOut_payload_0_5726 : _zz_dataOut_payload_0_5750);
  assign _zz_dataOut_payload_0_5900 = (_zz_dataOut_payload_0_5747 < _zz_dataOut_payload_0_5723);
  assign _zz_dataOut_payload_0_5901 = (_zz_dataOut_payload_0_5900 ? _zz_dataOut_payload_0_5747 : _zz_dataOut_payload_0_5723);
  assign _zz_dataOut_payload_0_5902 = (_zz_dataOut_payload_0_5900 ? _zz_dataOut_payload_0_5723 : _zz_dataOut_payload_0_5747);
  assign _zz_dataOut_payload_0_5903 = (_zz_dataOut_payload_0_5744 < _zz_dataOut_payload_0_5720);
  assign _zz_dataOut_payload_0_5904 = (_zz_dataOut_payload_0_5903 ? _zz_dataOut_payload_0_5744 : _zz_dataOut_payload_0_5720);
  assign _zz_dataOut_payload_0_5905 = (_zz_dataOut_payload_0_5903 ? _zz_dataOut_payload_0_5720 : _zz_dataOut_payload_0_5744);
  assign _zz_dataOut_payload_0_5906 = (_zz_dataOut_payload_0_5741 < _zz_dataOut_payload_0_5717);
  assign _zz_dataOut_payload_0_5907 = (_zz_dataOut_payload_0_5906 ? _zz_dataOut_payload_0_5741 : _zz_dataOut_payload_0_5717);
  assign _zz_dataOut_payload_0_5908 = (_zz_dataOut_payload_0_5906 ? _zz_dataOut_payload_0_5717 : _zz_dataOut_payload_0_5741);
  assign _zz_dataOut_payload_0_5909 = (_zz_dataOut_payload_0_5738 < _zz_dataOut_payload_0_5714);
  assign _zz_dataOut_payload_0_5910 = (_zz_dataOut_payload_0_5909 ? _zz_dataOut_payload_0_5738 : _zz_dataOut_payload_0_5714);
  assign _zz_dataOut_payload_0_5911 = (_zz_dataOut_payload_0_5909 ? _zz_dataOut_payload_0_5714 : _zz_dataOut_payload_0_5738);
  assign _zz_dataOut_payload_0_5912 = (_zz_dataOut_payload_0_5889 < _zz_dataOut_payload_0_5901);
  assign _zz_dataOut_payload_0_5913 = (_zz_dataOut_payload_0_5912 ? _zz_dataOut_payload_0_5889 : _zz_dataOut_payload_0_5901);
  assign _zz_dataOut_payload_0_5914 = (_zz_dataOut_payload_0_5912 ? _zz_dataOut_payload_0_5901 : _zz_dataOut_payload_0_5889);
  assign _zz_dataOut_payload_0_5915 = (_zz_dataOut_payload_0_5892 < _zz_dataOut_payload_0_5904);
  assign _zz_dataOut_payload_0_5916 = (_zz_dataOut_payload_0_5915 ? _zz_dataOut_payload_0_5892 : _zz_dataOut_payload_0_5904);
  assign _zz_dataOut_payload_0_5917 = (_zz_dataOut_payload_0_5915 ? _zz_dataOut_payload_0_5904 : _zz_dataOut_payload_0_5892);
  assign _zz_dataOut_payload_0_5918 = (_zz_dataOut_payload_0_5895 < _zz_dataOut_payload_0_5907);
  assign _zz_dataOut_payload_0_5919 = (_zz_dataOut_payload_0_5918 ? _zz_dataOut_payload_0_5895 : _zz_dataOut_payload_0_5907);
  assign _zz_dataOut_payload_0_5920 = (_zz_dataOut_payload_0_5918 ? _zz_dataOut_payload_0_5907 : _zz_dataOut_payload_0_5895);
  assign _zz_dataOut_payload_0_5921 = (_zz_dataOut_payload_0_5898 < _zz_dataOut_payload_0_5910);
  assign _zz_dataOut_payload_0_5922 = (_zz_dataOut_payload_0_5921 ? _zz_dataOut_payload_0_5898 : _zz_dataOut_payload_0_5910);
  assign _zz_dataOut_payload_0_5923 = (_zz_dataOut_payload_0_5921 ? _zz_dataOut_payload_0_5910 : _zz_dataOut_payload_0_5898);
  assign _zz_dataOut_payload_0_5924 = (_zz_dataOut_payload_0_5913 < _zz_dataOut_payload_0_5919);
  assign _zz_dataOut_payload_0_5925 = (_zz_dataOut_payload_0_5924 ? _zz_dataOut_payload_0_5913 : _zz_dataOut_payload_0_5919);
  assign _zz_dataOut_payload_0_5926 = (_zz_dataOut_payload_0_5924 ? _zz_dataOut_payload_0_5919 : _zz_dataOut_payload_0_5913);
  assign _zz_dataOut_payload_0_5927 = (_zz_dataOut_payload_0_5916 < _zz_dataOut_payload_0_5922);
  assign _zz_dataOut_payload_0_5928 = (_zz_dataOut_payload_0_5927 ? _zz_dataOut_payload_0_5916 : _zz_dataOut_payload_0_5922);
  assign _zz_dataOut_payload_0_5929 = (_zz_dataOut_payload_0_5927 ? _zz_dataOut_payload_0_5922 : _zz_dataOut_payload_0_5916);
  assign _zz_dataOut_payload_0_5930 = (_zz_dataOut_payload_0_5925 < _zz_dataOut_payload_0_5928);
  assign _zz_dataOut_payload_0_5931 = (_zz_dataOut_payload_0_5926 < _zz_dataOut_payload_0_5929);
  assign _zz_dataOut_payload_0_5936 = (_zz_dataOut_payload_0_5914 < _zz_dataOut_payload_0_5920);
  assign _zz_dataOut_payload_0_5937 = (_zz_dataOut_payload_0_5936 ? _zz_dataOut_payload_0_5914 : _zz_dataOut_payload_0_5920);
  assign _zz_dataOut_payload_0_5938 = (_zz_dataOut_payload_0_5936 ? _zz_dataOut_payload_0_5920 : _zz_dataOut_payload_0_5914);
  assign _zz_dataOut_payload_0_5939 = (_zz_dataOut_payload_0_5917 < _zz_dataOut_payload_0_5923);
  assign _zz_dataOut_payload_0_5940 = (_zz_dataOut_payload_0_5939 ? _zz_dataOut_payload_0_5917 : _zz_dataOut_payload_0_5923);
  assign _zz_dataOut_payload_0_5941 = (_zz_dataOut_payload_0_5939 ? _zz_dataOut_payload_0_5923 : _zz_dataOut_payload_0_5917);
  assign _zz_dataOut_payload_0_5942 = (_zz_dataOut_payload_0_5937 < _zz_dataOut_payload_0_5940);
  assign _zz_dataOut_payload_0_5943 = (_zz_dataOut_payload_0_5938 < _zz_dataOut_payload_0_5941);
  assign _zz_dataOut_payload_0_5956 = (_zz_dataOut_payload_0_5890 < _zz_dataOut_payload_0_5902);
  assign _zz_dataOut_payload_0_5957 = (_zz_dataOut_payload_0_5956 ? _zz_dataOut_payload_0_5890 : _zz_dataOut_payload_0_5902);
  assign _zz_dataOut_payload_0_5958 = (_zz_dataOut_payload_0_5956 ? _zz_dataOut_payload_0_5902 : _zz_dataOut_payload_0_5890);
  assign _zz_dataOut_payload_0_5959 = (_zz_dataOut_payload_0_5893 < _zz_dataOut_payload_0_5905);
  assign _zz_dataOut_payload_0_5960 = (_zz_dataOut_payload_0_5959 ? _zz_dataOut_payload_0_5893 : _zz_dataOut_payload_0_5905);
  assign _zz_dataOut_payload_0_5961 = (_zz_dataOut_payload_0_5959 ? _zz_dataOut_payload_0_5905 : _zz_dataOut_payload_0_5893);
  assign _zz_dataOut_payload_0_5962 = (_zz_dataOut_payload_0_5896 < _zz_dataOut_payload_0_5908);
  assign _zz_dataOut_payload_0_5963 = (_zz_dataOut_payload_0_5962 ? _zz_dataOut_payload_0_5896 : _zz_dataOut_payload_0_5908);
  assign _zz_dataOut_payload_0_5964 = (_zz_dataOut_payload_0_5962 ? _zz_dataOut_payload_0_5908 : _zz_dataOut_payload_0_5896);
  assign _zz_dataOut_payload_0_5965 = (_zz_dataOut_payload_0_5899 < _zz_dataOut_payload_0_5911);
  assign _zz_dataOut_payload_0_5966 = (_zz_dataOut_payload_0_5965 ? _zz_dataOut_payload_0_5899 : _zz_dataOut_payload_0_5911);
  assign _zz_dataOut_payload_0_5967 = (_zz_dataOut_payload_0_5965 ? _zz_dataOut_payload_0_5911 : _zz_dataOut_payload_0_5899);
  assign _zz_dataOut_payload_0_5968 = (_zz_dataOut_payload_0_5957 < _zz_dataOut_payload_0_5963);
  assign _zz_dataOut_payload_0_5969 = (_zz_dataOut_payload_0_5968 ? _zz_dataOut_payload_0_5957 : _zz_dataOut_payload_0_5963);
  assign _zz_dataOut_payload_0_5970 = (_zz_dataOut_payload_0_5968 ? _zz_dataOut_payload_0_5963 : _zz_dataOut_payload_0_5957);
  assign _zz_dataOut_payload_0_5971 = (_zz_dataOut_payload_0_5960 < _zz_dataOut_payload_0_5966);
  assign _zz_dataOut_payload_0_5972 = (_zz_dataOut_payload_0_5971 ? _zz_dataOut_payload_0_5960 : _zz_dataOut_payload_0_5966);
  assign _zz_dataOut_payload_0_5973 = (_zz_dataOut_payload_0_5971 ? _zz_dataOut_payload_0_5966 : _zz_dataOut_payload_0_5960);
  assign _zz_dataOut_payload_0_5974 = (_zz_dataOut_payload_0_5969 < _zz_dataOut_payload_0_5972);
  assign _zz_dataOut_payload_0_5975 = (_zz_dataOut_payload_0_5970 < _zz_dataOut_payload_0_5973);
  assign _zz_dataOut_payload_0_5980 = (_zz_dataOut_payload_0_5958 < _zz_dataOut_payload_0_5964);
  assign _zz_dataOut_payload_0_5981 = (_zz_dataOut_payload_0_5980 ? _zz_dataOut_payload_0_5958 : _zz_dataOut_payload_0_5964);
  assign _zz_dataOut_payload_0_5982 = (_zz_dataOut_payload_0_5980 ? _zz_dataOut_payload_0_5964 : _zz_dataOut_payload_0_5958);
  assign _zz_dataOut_payload_0_5983 = (_zz_dataOut_payload_0_5961 < _zz_dataOut_payload_0_5967);
  assign _zz_dataOut_payload_0_5984 = (_zz_dataOut_payload_0_5983 ? _zz_dataOut_payload_0_5961 : _zz_dataOut_payload_0_5967);
  assign _zz_dataOut_payload_0_5985 = (_zz_dataOut_payload_0_5983 ? _zz_dataOut_payload_0_5967 : _zz_dataOut_payload_0_5961);
  assign _zz_dataOut_payload_0_5986 = (_zz_dataOut_payload_0_5981 < _zz_dataOut_payload_0_5984);
  assign _zz_dataOut_payload_0_5987 = (_zz_dataOut_payload_0_5982 < _zz_dataOut_payload_0_5985);
  assign _zz_dataOut_payload_0_6048 = (_zz_dataOut_payload_0_5184 < _zz_dataOut_payload_0_5215);
  assign _zz_dataOut_payload_0_6049 = (_zz_dataOut_payload_0_6048 ? _zz_dataOut_payload_0_5184 : _zz_dataOut_payload_0_5215);
  assign _zz_dataOut_payload_0_6050 = (_zz_dataOut_payload_0_6048 ? _zz_dataOut_payload_0_5215 : _zz_dataOut_payload_0_5184);
  assign _zz_dataOut_payload_0_6051 = (_zz_dataOut_payload_0_5185 < _zz_dataOut_payload_0_5214);
  assign _zz_dataOut_payload_0_6052 = (_zz_dataOut_payload_0_6051 ? _zz_dataOut_payload_0_5185 : _zz_dataOut_payload_0_5214);
  assign _zz_dataOut_payload_0_6053 = (_zz_dataOut_payload_0_6051 ? _zz_dataOut_payload_0_5214 : _zz_dataOut_payload_0_5185);
  assign _zz_dataOut_payload_0_6054 = (_zz_dataOut_payload_0_5186 < _zz_dataOut_payload_0_5213);
  assign _zz_dataOut_payload_0_6055 = (_zz_dataOut_payload_0_6054 ? _zz_dataOut_payload_0_5186 : _zz_dataOut_payload_0_5213);
  assign _zz_dataOut_payload_0_6056 = (_zz_dataOut_payload_0_6054 ? _zz_dataOut_payload_0_5213 : _zz_dataOut_payload_0_5186);
  assign _zz_dataOut_payload_0_6057 = (_zz_dataOut_payload_0_5187 < _zz_dataOut_payload_0_5212);
  assign _zz_dataOut_payload_0_6058 = (_zz_dataOut_payload_0_6057 ? _zz_dataOut_payload_0_5187 : _zz_dataOut_payload_0_5212);
  assign _zz_dataOut_payload_0_6059 = (_zz_dataOut_payload_0_6057 ? _zz_dataOut_payload_0_5212 : _zz_dataOut_payload_0_5187);
  assign _zz_dataOut_payload_0_6060 = (_zz_dataOut_payload_0_5188 < _zz_dataOut_payload_0_5211);
  assign _zz_dataOut_payload_0_6061 = (_zz_dataOut_payload_0_6060 ? _zz_dataOut_payload_0_5188 : _zz_dataOut_payload_0_5211);
  assign _zz_dataOut_payload_0_6062 = (_zz_dataOut_payload_0_6060 ? _zz_dataOut_payload_0_5211 : _zz_dataOut_payload_0_5188);
  assign _zz_dataOut_payload_0_6063 = (_zz_dataOut_payload_0_5189 < _zz_dataOut_payload_0_5210);
  assign _zz_dataOut_payload_0_6064 = (_zz_dataOut_payload_0_6063 ? _zz_dataOut_payload_0_5189 : _zz_dataOut_payload_0_5210);
  assign _zz_dataOut_payload_0_6065 = (_zz_dataOut_payload_0_6063 ? _zz_dataOut_payload_0_5210 : _zz_dataOut_payload_0_5189);
  assign _zz_dataOut_payload_0_6066 = (_zz_dataOut_payload_0_5190 < _zz_dataOut_payload_0_5209);
  assign _zz_dataOut_payload_0_6067 = (_zz_dataOut_payload_0_6066 ? _zz_dataOut_payload_0_5190 : _zz_dataOut_payload_0_5209);
  assign _zz_dataOut_payload_0_6068 = (_zz_dataOut_payload_0_6066 ? _zz_dataOut_payload_0_5209 : _zz_dataOut_payload_0_5190);
  assign _zz_dataOut_payload_0_6069 = (_zz_dataOut_payload_0_5191 < _zz_dataOut_payload_0_5208);
  assign _zz_dataOut_payload_0_6070 = (_zz_dataOut_payload_0_6069 ? _zz_dataOut_payload_0_5191 : _zz_dataOut_payload_0_5208);
  assign _zz_dataOut_payload_0_6071 = (_zz_dataOut_payload_0_6069 ? _zz_dataOut_payload_0_5208 : _zz_dataOut_payload_0_5191);
  assign _zz_dataOut_payload_0_6072 = (_zz_dataOut_payload_0_5192 < _zz_dataOut_payload_0_5207);
  assign _zz_dataOut_payload_0_6073 = (_zz_dataOut_payload_0_6072 ? _zz_dataOut_payload_0_5192 : _zz_dataOut_payload_0_5207);
  assign _zz_dataOut_payload_0_6074 = (_zz_dataOut_payload_0_6072 ? _zz_dataOut_payload_0_5207 : _zz_dataOut_payload_0_5192);
  assign _zz_dataOut_payload_0_6075 = (_zz_dataOut_payload_0_5193 < _zz_dataOut_payload_0_5206);
  assign _zz_dataOut_payload_0_6076 = (_zz_dataOut_payload_0_6075 ? _zz_dataOut_payload_0_5193 : _zz_dataOut_payload_0_5206);
  assign _zz_dataOut_payload_0_6077 = (_zz_dataOut_payload_0_6075 ? _zz_dataOut_payload_0_5206 : _zz_dataOut_payload_0_5193);
  assign _zz_dataOut_payload_0_6078 = (_zz_dataOut_payload_0_5194 < _zz_dataOut_payload_0_5205);
  assign _zz_dataOut_payload_0_6079 = (_zz_dataOut_payload_0_6078 ? _zz_dataOut_payload_0_5194 : _zz_dataOut_payload_0_5205);
  assign _zz_dataOut_payload_0_6080 = (_zz_dataOut_payload_0_6078 ? _zz_dataOut_payload_0_5205 : _zz_dataOut_payload_0_5194);
  assign _zz_dataOut_payload_0_6081 = (_zz_dataOut_payload_0_5195 < _zz_dataOut_payload_0_5204);
  assign _zz_dataOut_payload_0_6082 = (_zz_dataOut_payload_0_6081 ? _zz_dataOut_payload_0_5195 : _zz_dataOut_payload_0_5204);
  assign _zz_dataOut_payload_0_6083 = (_zz_dataOut_payload_0_6081 ? _zz_dataOut_payload_0_5204 : _zz_dataOut_payload_0_5195);
  assign _zz_dataOut_payload_0_6084 = (_zz_dataOut_payload_0_5196 < _zz_dataOut_payload_0_5203);
  assign _zz_dataOut_payload_0_6085 = (_zz_dataOut_payload_0_6084 ? _zz_dataOut_payload_0_5196 : _zz_dataOut_payload_0_5203);
  assign _zz_dataOut_payload_0_6086 = (_zz_dataOut_payload_0_6084 ? _zz_dataOut_payload_0_5203 : _zz_dataOut_payload_0_5196);
  assign _zz_dataOut_payload_0_6087 = (_zz_dataOut_payload_0_5197 < _zz_dataOut_payload_0_5202);
  assign _zz_dataOut_payload_0_6088 = (_zz_dataOut_payload_0_6087 ? _zz_dataOut_payload_0_5197 : _zz_dataOut_payload_0_5202);
  assign _zz_dataOut_payload_0_6089 = (_zz_dataOut_payload_0_6087 ? _zz_dataOut_payload_0_5202 : _zz_dataOut_payload_0_5197);
  assign _zz_dataOut_payload_0_6090 = (_zz_dataOut_payload_0_5198 < _zz_dataOut_payload_0_5201);
  assign _zz_dataOut_payload_0_6091 = (_zz_dataOut_payload_0_6090 ? _zz_dataOut_payload_0_5198 : _zz_dataOut_payload_0_5201);
  assign _zz_dataOut_payload_0_6092 = (_zz_dataOut_payload_0_6090 ? _zz_dataOut_payload_0_5201 : _zz_dataOut_payload_0_5198);
  assign _zz_dataOut_payload_0_6093 = (_zz_dataOut_payload_0_5199 < _zz_dataOut_payload_0_5200);
  assign _zz_dataOut_payload_0_6094 = (_zz_dataOut_payload_0_6093 ? _zz_dataOut_payload_0_5199 : _zz_dataOut_payload_0_5200);
  assign _zz_dataOut_payload_0_6095 = (_zz_dataOut_payload_0_6093 ? _zz_dataOut_payload_0_5200 : _zz_dataOut_payload_0_5199);
  assign _zz_dataOut_payload_0_6096 = (_zz_dataOut_payload_0_6049 < _zz_dataOut_payload_0_6073);
  assign _zz_dataOut_payload_0_6097 = (_zz_dataOut_payload_0_6096 ? _zz_dataOut_payload_0_6049 : _zz_dataOut_payload_0_6073);
  assign _zz_dataOut_payload_0_6098 = (_zz_dataOut_payload_0_6096 ? _zz_dataOut_payload_0_6073 : _zz_dataOut_payload_0_6049);
  assign _zz_dataOut_payload_0_6099 = (_zz_dataOut_payload_0_6052 < _zz_dataOut_payload_0_6076);
  assign _zz_dataOut_payload_0_6100 = (_zz_dataOut_payload_0_6099 ? _zz_dataOut_payload_0_6052 : _zz_dataOut_payload_0_6076);
  assign _zz_dataOut_payload_0_6101 = (_zz_dataOut_payload_0_6099 ? _zz_dataOut_payload_0_6076 : _zz_dataOut_payload_0_6052);
  assign _zz_dataOut_payload_0_6102 = (_zz_dataOut_payload_0_6055 < _zz_dataOut_payload_0_6079);
  assign _zz_dataOut_payload_0_6103 = (_zz_dataOut_payload_0_6102 ? _zz_dataOut_payload_0_6055 : _zz_dataOut_payload_0_6079);
  assign _zz_dataOut_payload_0_6104 = (_zz_dataOut_payload_0_6102 ? _zz_dataOut_payload_0_6079 : _zz_dataOut_payload_0_6055);
  assign _zz_dataOut_payload_0_6105 = (_zz_dataOut_payload_0_6058 < _zz_dataOut_payload_0_6082);
  assign _zz_dataOut_payload_0_6106 = (_zz_dataOut_payload_0_6105 ? _zz_dataOut_payload_0_6058 : _zz_dataOut_payload_0_6082);
  assign _zz_dataOut_payload_0_6107 = (_zz_dataOut_payload_0_6105 ? _zz_dataOut_payload_0_6082 : _zz_dataOut_payload_0_6058);
  assign _zz_dataOut_payload_0_6108 = (_zz_dataOut_payload_0_6061 < _zz_dataOut_payload_0_6085);
  assign _zz_dataOut_payload_0_6109 = (_zz_dataOut_payload_0_6108 ? _zz_dataOut_payload_0_6061 : _zz_dataOut_payload_0_6085);
  assign _zz_dataOut_payload_0_6110 = (_zz_dataOut_payload_0_6108 ? _zz_dataOut_payload_0_6085 : _zz_dataOut_payload_0_6061);
  assign _zz_dataOut_payload_0_6111 = (_zz_dataOut_payload_0_6064 < _zz_dataOut_payload_0_6088);
  assign _zz_dataOut_payload_0_6112 = (_zz_dataOut_payload_0_6111 ? _zz_dataOut_payload_0_6064 : _zz_dataOut_payload_0_6088);
  assign _zz_dataOut_payload_0_6113 = (_zz_dataOut_payload_0_6111 ? _zz_dataOut_payload_0_6088 : _zz_dataOut_payload_0_6064);
  assign _zz_dataOut_payload_0_6114 = (_zz_dataOut_payload_0_6067 < _zz_dataOut_payload_0_6091);
  assign _zz_dataOut_payload_0_6115 = (_zz_dataOut_payload_0_6114 ? _zz_dataOut_payload_0_6067 : _zz_dataOut_payload_0_6091);
  assign _zz_dataOut_payload_0_6116 = (_zz_dataOut_payload_0_6114 ? _zz_dataOut_payload_0_6091 : _zz_dataOut_payload_0_6067);
  assign _zz_dataOut_payload_0_6117 = (_zz_dataOut_payload_0_6070 < _zz_dataOut_payload_0_6094);
  assign _zz_dataOut_payload_0_6118 = (_zz_dataOut_payload_0_6117 ? _zz_dataOut_payload_0_6070 : _zz_dataOut_payload_0_6094);
  assign _zz_dataOut_payload_0_6119 = (_zz_dataOut_payload_0_6117 ? _zz_dataOut_payload_0_6094 : _zz_dataOut_payload_0_6070);
  assign _zz_dataOut_payload_0_6120 = (_zz_dataOut_payload_0_6097 < _zz_dataOut_payload_0_6109);
  assign _zz_dataOut_payload_0_6121 = (_zz_dataOut_payload_0_6120 ? _zz_dataOut_payload_0_6097 : _zz_dataOut_payload_0_6109);
  assign _zz_dataOut_payload_0_6122 = (_zz_dataOut_payload_0_6120 ? _zz_dataOut_payload_0_6109 : _zz_dataOut_payload_0_6097);
  assign _zz_dataOut_payload_0_6123 = (_zz_dataOut_payload_0_6100 < _zz_dataOut_payload_0_6112);
  assign _zz_dataOut_payload_0_6124 = (_zz_dataOut_payload_0_6123 ? _zz_dataOut_payload_0_6100 : _zz_dataOut_payload_0_6112);
  assign _zz_dataOut_payload_0_6125 = (_zz_dataOut_payload_0_6123 ? _zz_dataOut_payload_0_6112 : _zz_dataOut_payload_0_6100);
  assign _zz_dataOut_payload_0_6126 = (_zz_dataOut_payload_0_6103 < _zz_dataOut_payload_0_6115);
  assign _zz_dataOut_payload_0_6127 = (_zz_dataOut_payload_0_6126 ? _zz_dataOut_payload_0_6103 : _zz_dataOut_payload_0_6115);
  assign _zz_dataOut_payload_0_6128 = (_zz_dataOut_payload_0_6126 ? _zz_dataOut_payload_0_6115 : _zz_dataOut_payload_0_6103);
  assign _zz_dataOut_payload_0_6129 = (_zz_dataOut_payload_0_6106 < _zz_dataOut_payload_0_6118);
  assign _zz_dataOut_payload_0_6130 = (_zz_dataOut_payload_0_6129 ? _zz_dataOut_payload_0_6106 : _zz_dataOut_payload_0_6118);
  assign _zz_dataOut_payload_0_6131 = (_zz_dataOut_payload_0_6129 ? _zz_dataOut_payload_0_6118 : _zz_dataOut_payload_0_6106);
  assign _zz_dataOut_payload_0_6132 = (_zz_dataOut_payload_0_6121 < _zz_dataOut_payload_0_6127);
  assign _zz_dataOut_payload_0_6133 = (_zz_dataOut_payload_0_6132 ? _zz_dataOut_payload_0_6121 : _zz_dataOut_payload_0_6127);
  assign _zz_dataOut_payload_0_6134 = (_zz_dataOut_payload_0_6132 ? _zz_dataOut_payload_0_6127 : _zz_dataOut_payload_0_6121);
  assign _zz_dataOut_payload_0_6135 = (_zz_dataOut_payload_0_6124 < _zz_dataOut_payload_0_6130);
  assign _zz_dataOut_payload_0_6136 = (_zz_dataOut_payload_0_6135 ? _zz_dataOut_payload_0_6124 : _zz_dataOut_payload_0_6130);
  assign _zz_dataOut_payload_0_6137 = (_zz_dataOut_payload_0_6135 ? _zz_dataOut_payload_0_6130 : _zz_dataOut_payload_0_6124);
  assign _zz_dataOut_payload_0_6138 = (_zz_dataOut_payload_0_6133 < _zz_dataOut_payload_0_6136);
  assign _zz_dataOut_payload_0_6139 = (_zz_dataOut_payload_0_6134 < _zz_dataOut_payload_0_6137);
  assign _zz_dataOut_payload_0_6144 = (_zz_dataOut_payload_0_6122 < _zz_dataOut_payload_0_6128);
  assign _zz_dataOut_payload_0_6145 = (_zz_dataOut_payload_0_6144 ? _zz_dataOut_payload_0_6122 : _zz_dataOut_payload_0_6128);
  assign _zz_dataOut_payload_0_6146 = (_zz_dataOut_payload_0_6144 ? _zz_dataOut_payload_0_6128 : _zz_dataOut_payload_0_6122);
  assign _zz_dataOut_payload_0_6147 = (_zz_dataOut_payload_0_6125 < _zz_dataOut_payload_0_6131);
  assign _zz_dataOut_payload_0_6148 = (_zz_dataOut_payload_0_6147 ? _zz_dataOut_payload_0_6125 : _zz_dataOut_payload_0_6131);
  assign _zz_dataOut_payload_0_6149 = (_zz_dataOut_payload_0_6147 ? _zz_dataOut_payload_0_6131 : _zz_dataOut_payload_0_6125);
  assign _zz_dataOut_payload_0_6150 = (_zz_dataOut_payload_0_6145 < _zz_dataOut_payload_0_6148);
  assign _zz_dataOut_payload_0_6151 = (_zz_dataOut_payload_0_6146 < _zz_dataOut_payload_0_6149);
  assign _zz_dataOut_payload_0_6164 = (_zz_dataOut_payload_0_6098 < _zz_dataOut_payload_0_6110);
  assign _zz_dataOut_payload_0_6165 = (_zz_dataOut_payload_0_6164 ? _zz_dataOut_payload_0_6098 : _zz_dataOut_payload_0_6110);
  assign _zz_dataOut_payload_0_6166 = (_zz_dataOut_payload_0_6164 ? _zz_dataOut_payload_0_6110 : _zz_dataOut_payload_0_6098);
  assign _zz_dataOut_payload_0_6167 = (_zz_dataOut_payload_0_6101 < _zz_dataOut_payload_0_6113);
  assign _zz_dataOut_payload_0_6168 = (_zz_dataOut_payload_0_6167 ? _zz_dataOut_payload_0_6101 : _zz_dataOut_payload_0_6113);
  assign _zz_dataOut_payload_0_6169 = (_zz_dataOut_payload_0_6167 ? _zz_dataOut_payload_0_6113 : _zz_dataOut_payload_0_6101);
  assign _zz_dataOut_payload_0_6170 = (_zz_dataOut_payload_0_6104 < _zz_dataOut_payload_0_6116);
  assign _zz_dataOut_payload_0_6171 = (_zz_dataOut_payload_0_6170 ? _zz_dataOut_payload_0_6104 : _zz_dataOut_payload_0_6116);
  assign _zz_dataOut_payload_0_6172 = (_zz_dataOut_payload_0_6170 ? _zz_dataOut_payload_0_6116 : _zz_dataOut_payload_0_6104);
  assign _zz_dataOut_payload_0_6173 = (_zz_dataOut_payload_0_6107 < _zz_dataOut_payload_0_6119);
  assign _zz_dataOut_payload_0_6174 = (_zz_dataOut_payload_0_6173 ? _zz_dataOut_payload_0_6107 : _zz_dataOut_payload_0_6119);
  assign _zz_dataOut_payload_0_6175 = (_zz_dataOut_payload_0_6173 ? _zz_dataOut_payload_0_6119 : _zz_dataOut_payload_0_6107);
  assign _zz_dataOut_payload_0_6176 = (_zz_dataOut_payload_0_6165 < _zz_dataOut_payload_0_6171);
  assign _zz_dataOut_payload_0_6177 = (_zz_dataOut_payload_0_6176 ? _zz_dataOut_payload_0_6165 : _zz_dataOut_payload_0_6171);
  assign _zz_dataOut_payload_0_6178 = (_zz_dataOut_payload_0_6176 ? _zz_dataOut_payload_0_6171 : _zz_dataOut_payload_0_6165);
  assign _zz_dataOut_payload_0_6179 = (_zz_dataOut_payload_0_6168 < _zz_dataOut_payload_0_6174);
  assign _zz_dataOut_payload_0_6180 = (_zz_dataOut_payload_0_6179 ? _zz_dataOut_payload_0_6168 : _zz_dataOut_payload_0_6174);
  assign _zz_dataOut_payload_0_6181 = (_zz_dataOut_payload_0_6179 ? _zz_dataOut_payload_0_6174 : _zz_dataOut_payload_0_6168);
  assign _zz_dataOut_payload_0_6182 = (_zz_dataOut_payload_0_6177 < _zz_dataOut_payload_0_6180);
  assign _zz_dataOut_payload_0_6183 = (_zz_dataOut_payload_0_6178 < _zz_dataOut_payload_0_6181);
  assign _zz_dataOut_payload_0_6188 = (_zz_dataOut_payload_0_6166 < _zz_dataOut_payload_0_6172);
  assign _zz_dataOut_payload_0_6189 = (_zz_dataOut_payload_0_6188 ? _zz_dataOut_payload_0_6166 : _zz_dataOut_payload_0_6172);
  assign _zz_dataOut_payload_0_6190 = (_zz_dataOut_payload_0_6188 ? _zz_dataOut_payload_0_6172 : _zz_dataOut_payload_0_6166);
  assign _zz_dataOut_payload_0_6191 = (_zz_dataOut_payload_0_6169 < _zz_dataOut_payload_0_6175);
  assign _zz_dataOut_payload_0_6192 = (_zz_dataOut_payload_0_6191 ? _zz_dataOut_payload_0_6169 : _zz_dataOut_payload_0_6175);
  assign _zz_dataOut_payload_0_6193 = (_zz_dataOut_payload_0_6191 ? _zz_dataOut_payload_0_6175 : _zz_dataOut_payload_0_6169);
  assign _zz_dataOut_payload_0_6194 = (_zz_dataOut_payload_0_6189 < _zz_dataOut_payload_0_6192);
  assign _zz_dataOut_payload_0_6195 = (_zz_dataOut_payload_0_6190 < _zz_dataOut_payload_0_6193);
  assign _zz_dataOut_payload_0_6224 = (_zz_dataOut_payload_0_6095 < _zz_dataOut_payload_0_6071);
  assign _zz_dataOut_payload_0_6225 = (_zz_dataOut_payload_0_6224 ? _zz_dataOut_payload_0_6095 : _zz_dataOut_payload_0_6071);
  assign _zz_dataOut_payload_0_6226 = (_zz_dataOut_payload_0_6224 ? _zz_dataOut_payload_0_6071 : _zz_dataOut_payload_0_6095);
  assign _zz_dataOut_payload_0_6227 = (_zz_dataOut_payload_0_6092 < _zz_dataOut_payload_0_6068);
  assign _zz_dataOut_payload_0_6228 = (_zz_dataOut_payload_0_6227 ? _zz_dataOut_payload_0_6092 : _zz_dataOut_payload_0_6068);
  assign _zz_dataOut_payload_0_6229 = (_zz_dataOut_payload_0_6227 ? _zz_dataOut_payload_0_6068 : _zz_dataOut_payload_0_6092);
  assign _zz_dataOut_payload_0_6230 = (_zz_dataOut_payload_0_6089 < _zz_dataOut_payload_0_6065);
  assign _zz_dataOut_payload_0_6231 = (_zz_dataOut_payload_0_6230 ? _zz_dataOut_payload_0_6089 : _zz_dataOut_payload_0_6065);
  assign _zz_dataOut_payload_0_6232 = (_zz_dataOut_payload_0_6230 ? _zz_dataOut_payload_0_6065 : _zz_dataOut_payload_0_6089);
  assign _zz_dataOut_payload_0_6233 = (_zz_dataOut_payload_0_6086 < _zz_dataOut_payload_0_6062);
  assign _zz_dataOut_payload_0_6234 = (_zz_dataOut_payload_0_6233 ? _zz_dataOut_payload_0_6086 : _zz_dataOut_payload_0_6062);
  assign _zz_dataOut_payload_0_6235 = (_zz_dataOut_payload_0_6233 ? _zz_dataOut_payload_0_6062 : _zz_dataOut_payload_0_6086);
  assign _zz_dataOut_payload_0_6236 = (_zz_dataOut_payload_0_6083 < _zz_dataOut_payload_0_6059);
  assign _zz_dataOut_payload_0_6237 = (_zz_dataOut_payload_0_6236 ? _zz_dataOut_payload_0_6083 : _zz_dataOut_payload_0_6059);
  assign _zz_dataOut_payload_0_6238 = (_zz_dataOut_payload_0_6236 ? _zz_dataOut_payload_0_6059 : _zz_dataOut_payload_0_6083);
  assign _zz_dataOut_payload_0_6239 = (_zz_dataOut_payload_0_6080 < _zz_dataOut_payload_0_6056);
  assign _zz_dataOut_payload_0_6240 = (_zz_dataOut_payload_0_6239 ? _zz_dataOut_payload_0_6080 : _zz_dataOut_payload_0_6056);
  assign _zz_dataOut_payload_0_6241 = (_zz_dataOut_payload_0_6239 ? _zz_dataOut_payload_0_6056 : _zz_dataOut_payload_0_6080);
  assign _zz_dataOut_payload_0_6242 = (_zz_dataOut_payload_0_6077 < _zz_dataOut_payload_0_6053);
  assign _zz_dataOut_payload_0_6243 = (_zz_dataOut_payload_0_6242 ? _zz_dataOut_payload_0_6077 : _zz_dataOut_payload_0_6053);
  assign _zz_dataOut_payload_0_6244 = (_zz_dataOut_payload_0_6242 ? _zz_dataOut_payload_0_6053 : _zz_dataOut_payload_0_6077);
  assign _zz_dataOut_payload_0_6245 = (_zz_dataOut_payload_0_6074 < _zz_dataOut_payload_0_6050);
  assign _zz_dataOut_payload_0_6246 = (_zz_dataOut_payload_0_6245 ? _zz_dataOut_payload_0_6074 : _zz_dataOut_payload_0_6050);
  assign _zz_dataOut_payload_0_6247 = (_zz_dataOut_payload_0_6245 ? _zz_dataOut_payload_0_6050 : _zz_dataOut_payload_0_6074);
  assign _zz_dataOut_payload_0_6248 = (_zz_dataOut_payload_0_6225 < _zz_dataOut_payload_0_6237);
  assign _zz_dataOut_payload_0_6249 = (_zz_dataOut_payload_0_6248 ? _zz_dataOut_payload_0_6225 : _zz_dataOut_payload_0_6237);
  assign _zz_dataOut_payload_0_6250 = (_zz_dataOut_payload_0_6248 ? _zz_dataOut_payload_0_6237 : _zz_dataOut_payload_0_6225);
  assign _zz_dataOut_payload_0_6251 = (_zz_dataOut_payload_0_6228 < _zz_dataOut_payload_0_6240);
  assign _zz_dataOut_payload_0_6252 = (_zz_dataOut_payload_0_6251 ? _zz_dataOut_payload_0_6228 : _zz_dataOut_payload_0_6240);
  assign _zz_dataOut_payload_0_6253 = (_zz_dataOut_payload_0_6251 ? _zz_dataOut_payload_0_6240 : _zz_dataOut_payload_0_6228);
  assign _zz_dataOut_payload_0_6254 = (_zz_dataOut_payload_0_6231 < _zz_dataOut_payload_0_6243);
  assign _zz_dataOut_payload_0_6255 = (_zz_dataOut_payload_0_6254 ? _zz_dataOut_payload_0_6231 : _zz_dataOut_payload_0_6243);
  assign _zz_dataOut_payload_0_6256 = (_zz_dataOut_payload_0_6254 ? _zz_dataOut_payload_0_6243 : _zz_dataOut_payload_0_6231);
  assign _zz_dataOut_payload_0_6257 = (_zz_dataOut_payload_0_6234 < _zz_dataOut_payload_0_6246);
  assign _zz_dataOut_payload_0_6258 = (_zz_dataOut_payload_0_6257 ? _zz_dataOut_payload_0_6234 : _zz_dataOut_payload_0_6246);
  assign _zz_dataOut_payload_0_6259 = (_zz_dataOut_payload_0_6257 ? _zz_dataOut_payload_0_6246 : _zz_dataOut_payload_0_6234);
  assign _zz_dataOut_payload_0_6260 = (_zz_dataOut_payload_0_6249 < _zz_dataOut_payload_0_6255);
  assign _zz_dataOut_payload_0_6261 = (_zz_dataOut_payload_0_6260 ? _zz_dataOut_payload_0_6249 : _zz_dataOut_payload_0_6255);
  assign _zz_dataOut_payload_0_6262 = (_zz_dataOut_payload_0_6260 ? _zz_dataOut_payload_0_6255 : _zz_dataOut_payload_0_6249);
  assign _zz_dataOut_payload_0_6263 = (_zz_dataOut_payload_0_6252 < _zz_dataOut_payload_0_6258);
  assign _zz_dataOut_payload_0_6264 = (_zz_dataOut_payload_0_6263 ? _zz_dataOut_payload_0_6252 : _zz_dataOut_payload_0_6258);
  assign _zz_dataOut_payload_0_6265 = (_zz_dataOut_payload_0_6263 ? _zz_dataOut_payload_0_6258 : _zz_dataOut_payload_0_6252);
  assign _zz_dataOut_payload_0_6266 = (_zz_dataOut_payload_0_6261 < _zz_dataOut_payload_0_6264);
  assign _zz_dataOut_payload_0_6267 = (_zz_dataOut_payload_0_6262 < _zz_dataOut_payload_0_6265);
  assign _zz_dataOut_payload_0_6272 = (_zz_dataOut_payload_0_6250 < _zz_dataOut_payload_0_6256);
  assign _zz_dataOut_payload_0_6273 = (_zz_dataOut_payload_0_6272 ? _zz_dataOut_payload_0_6250 : _zz_dataOut_payload_0_6256);
  assign _zz_dataOut_payload_0_6274 = (_zz_dataOut_payload_0_6272 ? _zz_dataOut_payload_0_6256 : _zz_dataOut_payload_0_6250);
  assign _zz_dataOut_payload_0_6275 = (_zz_dataOut_payload_0_6253 < _zz_dataOut_payload_0_6259);
  assign _zz_dataOut_payload_0_6276 = (_zz_dataOut_payload_0_6275 ? _zz_dataOut_payload_0_6253 : _zz_dataOut_payload_0_6259);
  assign _zz_dataOut_payload_0_6277 = (_zz_dataOut_payload_0_6275 ? _zz_dataOut_payload_0_6259 : _zz_dataOut_payload_0_6253);
  assign _zz_dataOut_payload_0_6278 = (_zz_dataOut_payload_0_6273 < _zz_dataOut_payload_0_6276);
  assign _zz_dataOut_payload_0_6279 = (_zz_dataOut_payload_0_6274 < _zz_dataOut_payload_0_6277);
  assign _zz_dataOut_payload_0_6292 = (_zz_dataOut_payload_0_6226 < _zz_dataOut_payload_0_6238);
  assign _zz_dataOut_payload_0_6293 = (_zz_dataOut_payload_0_6292 ? _zz_dataOut_payload_0_6226 : _zz_dataOut_payload_0_6238);
  assign _zz_dataOut_payload_0_6294 = (_zz_dataOut_payload_0_6292 ? _zz_dataOut_payload_0_6238 : _zz_dataOut_payload_0_6226);
  assign _zz_dataOut_payload_0_6295 = (_zz_dataOut_payload_0_6229 < _zz_dataOut_payload_0_6241);
  assign _zz_dataOut_payload_0_6296 = (_zz_dataOut_payload_0_6295 ? _zz_dataOut_payload_0_6229 : _zz_dataOut_payload_0_6241);
  assign _zz_dataOut_payload_0_6297 = (_zz_dataOut_payload_0_6295 ? _zz_dataOut_payload_0_6241 : _zz_dataOut_payload_0_6229);
  assign _zz_dataOut_payload_0_6298 = (_zz_dataOut_payload_0_6232 < _zz_dataOut_payload_0_6244);
  assign _zz_dataOut_payload_0_6299 = (_zz_dataOut_payload_0_6298 ? _zz_dataOut_payload_0_6232 : _zz_dataOut_payload_0_6244);
  assign _zz_dataOut_payload_0_6300 = (_zz_dataOut_payload_0_6298 ? _zz_dataOut_payload_0_6244 : _zz_dataOut_payload_0_6232);
  assign _zz_dataOut_payload_0_6301 = (_zz_dataOut_payload_0_6235 < _zz_dataOut_payload_0_6247);
  assign _zz_dataOut_payload_0_6302 = (_zz_dataOut_payload_0_6301 ? _zz_dataOut_payload_0_6235 : _zz_dataOut_payload_0_6247);
  assign _zz_dataOut_payload_0_6303 = (_zz_dataOut_payload_0_6301 ? _zz_dataOut_payload_0_6247 : _zz_dataOut_payload_0_6235);
  assign _zz_dataOut_payload_0_6304 = (_zz_dataOut_payload_0_6293 < _zz_dataOut_payload_0_6299);
  assign _zz_dataOut_payload_0_6305 = (_zz_dataOut_payload_0_6304 ? _zz_dataOut_payload_0_6293 : _zz_dataOut_payload_0_6299);
  assign _zz_dataOut_payload_0_6306 = (_zz_dataOut_payload_0_6304 ? _zz_dataOut_payload_0_6299 : _zz_dataOut_payload_0_6293);
  assign _zz_dataOut_payload_0_6307 = (_zz_dataOut_payload_0_6296 < _zz_dataOut_payload_0_6302);
  assign _zz_dataOut_payload_0_6308 = (_zz_dataOut_payload_0_6307 ? _zz_dataOut_payload_0_6296 : _zz_dataOut_payload_0_6302);
  assign _zz_dataOut_payload_0_6309 = (_zz_dataOut_payload_0_6307 ? _zz_dataOut_payload_0_6302 : _zz_dataOut_payload_0_6296);
  assign _zz_dataOut_payload_0_6310 = (_zz_dataOut_payload_0_6305 < _zz_dataOut_payload_0_6308);
  assign _zz_dataOut_payload_0_6311 = (_zz_dataOut_payload_0_6306 < _zz_dataOut_payload_0_6309);
  assign _zz_dataOut_payload_0_6316 = (_zz_dataOut_payload_0_6294 < _zz_dataOut_payload_0_6300);
  assign _zz_dataOut_payload_0_6317 = (_zz_dataOut_payload_0_6316 ? _zz_dataOut_payload_0_6294 : _zz_dataOut_payload_0_6300);
  assign _zz_dataOut_payload_0_6318 = (_zz_dataOut_payload_0_6316 ? _zz_dataOut_payload_0_6300 : _zz_dataOut_payload_0_6294);
  assign _zz_dataOut_payload_0_6319 = (_zz_dataOut_payload_0_6297 < _zz_dataOut_payload_0_6303);
  assign _zz_dataOut_payload_0_6320 = (_zz_dataOut_payload_0_6319 ? _zz_dataOut_payload_0_6297 : _zz_dataOut_payload_0_6303);
  assign _zz_dataOut_payload_0_6321 = (_zz_dataOut_payload_0_6319 ? _zz_dataOut_payload_0_6303 : _zz_dataOut_payload_0_6297);
  assign _zz_dataOut_payload_0_6322 = (_zz_dataOut_payload_0_6317 < _zz_dataOut_payload_0_6320);
  assign _zz_dataOut_payload_0_6323 = (_zz_dataOut_payload_0_6318 < _zz_dataOut_payload_0_6321);
  assign _zz_dataOut_payload_0_6384 = (_zz_dataOut_payload_0_5216 < _zz_dataOut_payload_0_5247);
  assign _zz_dataOut_payload_0_6385 = (_zz_dataOut_payload_0_6384 ? _zz_dataOut_payload_0_5216 : _zz_dataOut_payload_0_5247);
  assign _zz_dataOut_payload_0_6386 = (_zz_dataOut_payload_0_6384 ? _zz_dataOut_payload_0_5247 : _zz_dataOut_payload_0_5216);
  assign _zz_dataOut_payload_0_6387 = (_zz_dataOut_payload_0_5217 < _zz_dataOut_payload_0_5246);
  assign _zz_dataOut_payload_0_6388 = (_zz_dataOut_payload_0_6387 ? _zz_dataOut_payload_0_5217 : _zz_dataOut_payload_0_5246);
  assign _zz_dataOut_payload_0_6389 = (_zz_dataOut_payload_0_6387 ? _zz_dataOut_payload_0_5246 : _zz_dataOut_payload_0_5217);
  assign _zz_dataOut_payload_0_6390 = (_zz_dataOut_payload_0_5218 < _zz_dataOut_payload_0_5245);
  assign _zz_dataOut_payload_0_6391 = (_zz_dataOut_payload_0_6390 ? _zz_dataOut_payload_0_5218 : _zz_dataOut_payload_0_5245);
  assign _zz_dataOut_payload_0_6392 = (_zz_dataOut_payload_0_6390 ? _zz_dataOut_payload_0_5245 : _zz_dataOut_payload_0_5218);
  assign _zz_dataOut_payload_0_6393 = (_zz_dataOut_payload_0_5219 < _zz_dataOut_payload_0_5244);
  assign _zz_dataOut_payload_0_6394 = (_zz_dataOut_payload_0_6393 ? _zz_dataOut_payload_0_5219 : _zz_dataOut_payload_0_5244);
  assign _zz_dataOut_payload_0_6395 = (_zz_dataOut_payload_0_6393 ? _zz_dataOut_payload_0_5244 : _zz_dataOut_payload_0_5219);
  assign _zz_dataOut_payload_0_6396 = (_zz_dataOut_payload_0_5220 < _zz_dataOut_payload_0_5243);
  assign _zz_dataOut_payload_0_6397 = (_zz_dataOut_payload_0_6396 ? _zz_dataOut_payload_0_5220 : _zz_dataOut_payload_0_5243);
  assign _zz_dataOut_payload_0_6398 = (_zz_dataOut_payload_0_6396 ? _zz_dataOut_payload_0_5243 : _zz_dataOut_payload_0_5220);
  assign _zz_dataOut_payload_0_6399 = (_zz_dataOut_payload_0_5221 < _zz_dataOut_payload_0_5242);
  assign _zz_dataOut_payload_0_6400 = (_zz_dataOut_payload_0_6399 ? _zz_dataOut_payload_0_5221 : _zz_dataOut_payload_0_5242);
  assign _zz_dataOut_payload_0_6401 = (_zz_dataOut_payload_0_6399 ? _zz_dataOut_payload_0_5242 : _zz_dataOut_payload_0_5221);
  assign _zz_dataOut_payload_0_6402 = (_zz_dataOut_payload_0_5222 < _zz_dataOut_payload_0_5241);
  assign _zz_dataOut_payload_0_6403 = (_zz_dataOut_payload_0_6402 ? _zz_dataOut_payload_0_5222 : _zz_dataOut_payload_0_5241);
  assign _zz_dataOut_payload_0_6404 = (_zz_dataOut_payload_0_6402 ? _zz_dataOut_payload_0_5241 : _zz_dataOut_payload_0_5222);
  assign _zz_dataOut_payload_0_6405 = (_zz_dataOut_payload_0_5223 < _zz_dataOut_payload_0_5240);
  assign _zz_dataOut_payload_0_6406 = (_zz_dataOut_payload_0_6405 ? _zz_dataOut_payload_0_5223 : _zz_dataOut_payload_0_5240);
  assign _zz_dataOut_payload_0_6407 = (_zz_dataOut_payload_0_6405 ? _zz_dataOut_payload_0_5240 : _zz_dataOut_payload_0_5223);
  assign _zz_dataOut_payload_0_6408 = (_zz_dataOut_payload_0_5224 < _zz_dataOut_payload_0_5239);
  assign _zz_dataOut_payload_0_6409 = (_zz_dataOut_payload_0_6408 ? _zz_dataOut_payload_0_5224 : _zz_dataOut_payload_0_5239);
  assign _zz_dataOut_payload_0_6410 = (_zz_dataOut_payload_0_6408 ? _zz_dataOut_payload_0_5239 : _zz_dataOut_payload_0_5224);
  assign _zz_dataOut_payload_0_6411 = (_zz_dataOut_payload_0_5225 < _zz_dataOut_payload_0_5238);
  assign _zz_dataOut_payload_0_6412 = (_zz_dataOut_payload_0_6411 ? _zz_dataOut_payload_0_5225 : _zz_dataOut_payload_0_5238);
  assign _zz_dataOut_payload_0_6413 = (_zz_dataOut_payload_0_6411 ? _zz_dataOut_payload_0_5238 : _zz_dataOut_payload_0_5225);
  assign _zz_dataOut_payload_0_6414 = (_zz_dataOut_payload_0_5226 < _zz_dataOut_payload_0_5237);
  assign _zz_dataOut_payload_0_6415 = (_zz_dataOut_payload_0_6414 ? _zz_dataOut_payload_0_5226 : _zz_dataOut_payload_0_5237);
  assign _zz_dataOut_payload_0_6416 = (_zz_dataOut_payload_0_6414 ? _zz_dataOut_payload_0_5237 : _zz_dataOut_payload_0_5226);
  assign _zz_dataOut_payload_0_6417 = (_zz_dataOut_payload_0_5227 < _zz_dataOut_payload_0_5236);
  assign _zz_dataOut_payload_0_6418 = (_zz_dataOut_payload_0_6417 ? _zz_dataOut_payload_0_5227 : _zz_dataOut_payload_0_5236);
  assign _zz_dataOut_payload_0_6419 = (_zz_dataOut_payload_0_6417 ? _zz_dataOut_payload_0_5236 : _zz_dataOut_payload_0_5227);
  assign _zz_dataOut_payload_0_6420 = (_zz_dataOut_payload_0_5228 < _zz_dataOut_payload_0_5235);
  assign _zz_dataOut_payload_0_6421 = (_zz_dataOut_payload_0_6420 ? _zz_dataOut_payload_0_5228 : _zz_dataOut_payload_0_5235);
  assign _zz_dataOut_payload_0_6422 = (_zz_dataOut_payload_0_6420 ? _zz_dataOut_payload_0_5235 : _zz_dataOut_payload_0_5228);
  assign _zz_dataOut_payload_0_6423 = (_zz_dataOut_payload_0_5229 < _zz_dataOut_payload_0_5234);
  assign _zz_dataOut_payload_0_6424 = (_zz_dataOut_payload_0_6423 ? _zz_dataOut_payload_0_5229 : _zz_dataOut_payload_0_5234);
  assign _zz_dataOut_payload_0_6425 = (_zz_dataOut_payload_0_6423 ? _zz_dataOut_payload_0_5234 : _zz_dataOut_payload_0_5229);
  assign _zz_dataOut_payload_0_6426 = (_zz_dataOut_payload_0_5230 < _zz_dataOut_payload_0_5233);
  assign _zz_dataOut_payload_0_6427 = (_zz_dataOut_payload_0_6426 ? _zz_dataOut_payload_0_5230 : _zz_dataOut_payload_0_5233);
  assign _zz_dataOut_payload_0_6428 = (_zz_dataOut_payload_0_6426 ? _zz_dataOut_payload_0_5233 : _zz_dataOut_payload_0_5230);
  assign _zz_dataOut_payload_0_6429 = (_zz_dataOut_payload_0_5231 < _zz_dataOut_payload_0_5232);
  assign _zz_dataOut_payload_0_6430 = (_zz_dataOut_payload_0_6429 ? _zz_dataOut_payload_0_5231 : _zz_dataOut_payload_0_5232);
  assign _zz_dataOut_payload_0_6431 = (_zz_dataOut_payload_0_6429 ? _zz_dataOut_payload_0_5232 : _zz_dataOut_payload_0_5231);
  assign _zz_dataOut_payload_0_6432 = (_zz_dataOut_payload_0_6385 < _zz_dataOut_payload_0_6409);
  assign _zz_dataOut_payload_0_6433 = (_zz_dataOut_payload_0_6432 ? _zz_dataOut_payload_0_6385 : _zz_dataOut_payload_0_6409);
  assign _zz_dataOut_payload_0_6434 = (_zz_dataOut_payload_0_6432 ? _zz_dataOut_payload_0_6409 : _zz_dataOut_payload_0_6385);
  assign _zz_dataOut_payload_0_6435 = (_zz_dataOut_payload_0_6388 < _zz_dataOut_payload_0_6412);
  assign _zz_dataOut_payload_0_6436 = (_zz_dataOut_payload_0_6435 ? _zz_dataOut_payload_0_6388 : _zz_dataOut_payload_0_6412);
  assign _zz_dataOut_payload_0_6437 = (_zz_dataOut_payload_0_6435 ? _zz_dataOut_payload_0_6412 : _zz_dataOut_payload_0_6388);
  assign _zz_dataOut_payload_0_6438 = (_zz_dataOut_payload_0_6391 < _zz_dataOut_payload_0_6415);
  assign _zz_dataOut_payload_0_6439 = (_zz_dataOut_payload_0_6438 ? _zz_dataOut_payload_0_6391 : _zz_dataOut_payload_0_6415);
  assign _zz_dataOut_payload_0_6440 = (_zz_dataOut_payload_0_6438 ? _zz_dataOut_payload_0_6415 : _zz_dataOut_payload_0_6391);
  assign _zz_dataOut_payload_0_6441 = (_zz_dataOut_payload_0_6394 < _zz_dataOut_payload_0_6418);
  assign _zz_dataOut_payload_0_6442 = (_zz_dataOut_payload_0_6441 ? _zz_dataOut_payload_0_6394 : _zz_dataOut_payload_0_6418);
  assign _zz_dataOut_payload_0_6443 = (_zz_dataOut_payload_0_6441 ? _zz_dataOut_payload_0_6418 : _zz_dataOut_payload_0_6394);
  assign _zz_dataOut_payload_0_6444 = (_zz_dataOut_payload_0_6397 < _zz_dataOut_payload_0_6421);
  assign _zz_dataOut_payload_0_6445 = (_zz_dataOut_payload_0_6444 ? _zz_dataOut_payload_0_6397 : _zz_dataOut_payload_0_6421);
  assign _zz_dataOut_payload_0_6446 = (_zz_dataOut_payload_0_6444 ? _zz_dataOut_payload_0_6421 : _zz_dataOut_payload_0_6397);
  assign _zz_dataOut_payload_0_6447 = (_zz_dataOut_payload_0_6400 < _zz_dataOut_payload_0_6424);
  assign _zz_dataOut_payload_0_6448 = (_zz_dataOut_payload_0_6447 ? _zz_dataOut_payload_0_6400 : _zz_dataOut_payload_0_6424);
  assign _zz_dataOut_payload_0_6449 = (_zz_dataOut_payload_0_6447 ? _zz_dataOut_payload_0_6424 : _zz_dataOut_payload_0_6400);
  assign _zz_dataOut_payload_0_6450 = (_zz_dataOut_payload_0_6403 < _zz_dataOut_payload_0_6427);
  assign _zz_dataOut_payload_0_6451 = (_zz_dataOut_payload_0_6450 ? _zz_dataOut_payload_0_6403 : _zz_dataOut_payload_0_6427);
  assign _zz_dataOut_payload_0_6452 = (_zz_dataOut_payload_0_6450 ? _zz_dataOut_payload_0_6427 : _zz_dataOut_payload_0_6403);
  assign _zz_dataOut_payload_0_6453 = (_zz_dataOut_payload_0_6406 < _zz_dataOut_payload_0_6430);
  assign _zz_dataOut_payload_0_6454 = (_zz_dataOut_payload_0_6453 ? _zz_dataOut_payload_0_6406 : _zz_dataOut_payload_0_6430);
  assign _zz_dataOut_payload_0_6455 = (_zz_dataOut_payload_0_6453 ? _zz_dataOut_payload_0_6430 : _zz_dataOut_payload_0_6406);
  assign _zz_dataOut_payload_0_6456 = (_zz_dataOut_payload_0_6433 < _zz_dataOut_payload_0_6445);
  assign _zz_dataOut_payload_0_6457 = (_zz_dataOut_payload_0_6456 ? _zz_dataOut_payload_0_6433 : _zz_dataOut_payload_0_6445);
  assign _zz_dataOut_payload_0_6458 = (_zz_dataOut_payload_0_6456 ? _zz_dataOut_payload_0_6445 : _zz_dataOut_payload_0_6433);
  assign _zz_dataOut_payload_0_6459 = (_zz_dataOut_payload_0_6436 < _zz_dataOut_payload_0_6448);
  assign _zz_dataOut_payload_0_6460 = (_zz_dataOut_payload_0_6459 ? _zz_dataOut_payload_0_6436 : _zz_dataOut_payload_0_6448);
  assign _zz_dataOut_payload_0_6461 = (_zz_dataOut_payload_0_6459 ? _zz_dataOut_payload_0_6448 : _zz_dataOut_payload_0_6436);
  assign _zz_dataOut_payload_0_6462 = (_zz_dataOut_payload_0_6439 < _zz_dataOut_payload_0_6451);
  assign _zz_dataOut_payload_0_6463 = (_zz_dataOut_payload_0_6462 ? _zz_dataOut_payload_0_6439 : _zz_dataOut_payload_0_6451);
  assign _zz_dataOut_payload_0_6464 = (_zz_dataOut_payload_0_6462 ? _zz_dataOut_payload_0_6451 : _zz_dataOut_payload_0_6439);
  assign _zz_dataOut_payload_0_6465 = (_zz_dataOut_payload_0_6442 < _zz_dataOut_payload_0_6454);
  assign _zz_dataOut_payload_0_6466 = (_zz_dataOut_payload_0_6465 ? _zz_dataOut_payload_0_6442 : _zz_dataOut_payload_0_6454);
  assign _zz_dataOut_payload_0_6467 = (_zz_dataOut_payload_0_6465 ? _zz_dataOut_payload_0_6454 : _zz_dataOut_payload_0_6442);
  assign _zz_dataOut_payload_0_6468 = (_zz_dataOut_payload_0_6457 < _zz_dataOut_payload_0_6463);
  assign _zz_dataOut_payload_0_6469 = (_zz_dataOut_payload_0_6468 ? _zz_dataOut_payload_0_6457 : _zz_dataOut_payload_0_6463);
  assign _zz_dataOut_payload_0_6470 = (_zz_dataOut_payload_0_6468 ? _zz_dataOut_payload_0_6463 : _zz_dataOut_payload_0_6457);
  assign _zz_dataOut_payload_0_6471 = (_zz_dataOut_payload_0_6460 < _zz_dataOut_payload_0_6466);
  assign _zz_dataOut_payload_0_6472 = (_zz_dataOut_payload_0_6471 ? _zz_dataOut_payload_0_6460 : _zz_dataOut_payload_0_6466);
  assign _zz_dataOut_payload_0_6473 = (_zz_dataOut_payload_0_6471 ? _zz_dataOut_payload_0_6466 : _zz_dataOut_payload_0_6460);
  assign _zz_dataOut_payload_0_6474 = (_zz_dataOut_payload_0_6469 < _zz_dataOut_payload_0_6472);
  assign _zz_dataOut_payload_0_6475 = (_zz_dataOut_payload_0_6470 < _zz_dataOut_payload_0_6473);
  assign _zz_dataOut_payload_0_6480 = (_zz_dataOut_payload_0_6458 < _zz_dataOut_payload_0_6464);
  assign _zz_dataOut_payload_0_6481 = (_zz_dataOut_payload_0_6480 ? _zz_dataOut_payload_0_6458 : _zz_dataOut_payload_0_6464);
  assign _zz_dataOut_payload_0_6482 = (_zz_dataOut_payload_0_6480 ? _zz_dataOut_payload_0_6464 : _zz_dataOut_payload_0_6458);
  assign _zz_dataOut_payload_0_6483 = (_zz_dataOut_payload_0_6461 < _zz_dataOut_payload_0_6467);
  assign _zz_dataOut_payload_0_6484 = (_zz_dataOut_payload_0_6483 ? _zz_dataOut_payload_0_6461 : _zz_dataOut_payload_0_6467);
  assign _zz_dataOut_payload_0_6485 = (_zz_dataOut_payload_0_6483 ? _zz_dataOut_payload_0_6467 : _zz_dataOut_payload_0_6461);
  assign _zz_dataOut_payload_0_6486 = (_zz_dataOut_payload_0_6481 < _zz_dataOut_payload_0_6484);
  assign _zz_dataOut_payload_0_6487 = (_zz_dataOut_payload_0_6482 < _zz_dataOut_payload_0_6485);
  assign _zz_dataOut_payload_0_6500 = (_zz_dataOut_payload_0_6434 < _zz_dataOut_payload_0_6446);
  assign _zz_dataOut_payload_0_6501 = (_zz_dataOut_payload_0_6500 ? _zz_dataOut_payload_0_6434 : _zz_dataOut_payload_0_6446);
  assign _zz_dataOut_payload_0_6502 = (_zz_dataOut_payload_0_6500 ? _zz_dataOut_payload_0_6446 : _zz_dataOut_payload_0_6434);
  assign _zz_dataOut_payload_0_6503 = (_zz_dataOut_payload_0_6437 < _zz_dataOut_payload_0_6449);
  assign _zz_dataOut_payload_0_6504 = (_zz_dataOut_payload_0_6503 ? _zz_dataOut_payload_0_6437 : _zz_dataOut_payload_0_6449);
  assign _zz_dataOut_payload_0_6505 = (_zz_dataOut_payload_0_6503 ? _zz_dataOut_payload_0_6449 : _zz_dataOut_payload_0_6437);
  assign _zz_dataOut_payload_0_6506 = (_zz_dataOut_payload_0_6440 < _zz_dataOut_payload_0_6452);
  assign _zz_dataOut_payload_0_6507 = (_zz_dataOut_payload_0_6506 ? _zz_dataOut_payload_0_6440 : _zz_dataOut_payload_0_6452);
  assign _zz_dataOut_payload_0_6508 = (_zz_dataOut_payload_0_6506 ? _zz_dataOut_payload_0_6452 : _zz_dataOut_payload_0_6440);
  assign _zz_dataOut_payload_0_6509 = (_zz_dataOut_payload_0_6443 < _zz_dataOut_payload_0_6455);
  assign _zz_dataOut_payload_0_6510 = (_zz_dataOut_payload_0_6509 ? _zz_dataOut_payload_0_6443 : _zz_dataOut_payload_0_6455);
  assign _zz_dataOut_payload_0_6511 = (_zz_dataOut_payload_0_6509 ? _zz_dataOut_payload_0_6455 : _zz_dataOut_payload_0_6443);
  assign _zz_dataOut_payload_0_6512 = (_zz_dataOut_payload_0_6501 < _zz_dataOut_payload_0_6507);
  assign _zz_dataOut_payload_0_6513 = (_zz_dataOut_payload_0_6512 ? _zz_dataOut_payload_0_6501 : _zz_dataOut_payload_0_6507);
  assign _zz_dataOut_payload_0_6514 = (_zz_dataOut_payload_0_6512 ? _zz_dataOut_payload_0_6507 : _zz_dataOut_payload_0_6501);
  assign _zz_dataOut_payload_0_6515 = (_zz_dataOut_payload_0_6504 < _zz_dataOut_payload_0_6510);
  assign _zz_dataOut_payload_0_6516 = (_zz_dataOut_payload_0_6515 ? _zz_dataOut_payload_0_6504 : _zz_dataOut_payload_0_6510);
  assign _zz_dataOut_payload_0_6517 = (_zz_dataOut_payload_0_6515 ? _zz_dataOut_payload_0_6510 : _zz_dataOut_payload_0_6504);
  assign _zz_dataOut_payload_0_6518 = (_zz_dataOut_payload_0_6513 < _zz_dataOut_payload_0_6516);
  assign _zz_dataOut_payload_0_6519 = (_zz_dataOut_payload_0_6514 < _zz_dataOut_payload_0_6517);
  assign _zz_dataOut_payload_0_6524 = (_zz_dataOut_payload_0_6502 < _zz_dataOut_payload_0_6508);
  assign _zz_dataOut_payload_0_6525 = (_zz_dataOut_payload_0_6524 ? _zz_dataOut_payload_0_6502 : _zz_dataOut_payload_0_6508);
  assign _zz_dataOut_payload_0_6526 = (_zz_dataOut_payload_0_6524 ? _zz_dataOut_payload_0_6508 : _zz_dataOut_payload_0_6502);
  assign _zz_dataOut_payload_0_6527 = (_zz_dataOut_payload_0_6505 < _zz_dataOut_payload_0_6511);
  assign _zz_dataOut_payload_0_6528 = (_zz_dataOut_payload_0_6527 ? _zz_dataOut_payload_0_6505 : _zz_dataOut_payload_0_6511);
  assign _zz_dataOut_payload_0_6529 = (_zz_dataOut_payload_0_6527 ? _zz_dataOut_payload_0_6511 : _zz_dataOut_payload_0_6505);
  assign _zz_dataOut_payload_0_6530 = (_zz_dataOut_payload_0_6525 < _zz_dataOut_payload_0_6528);
  assign _zz_dataOut_payload_0_6531 = (_zz_dataOut_payload_0_6526 < _zz_dataOut_payload_0_6529);
  assign _zz_dataOut_payload_0_6560 = (_zz_dataOut_payload_0_6431 < _zz_dataOut_payload_0_6407);
  assign _zz_dataOut_payload_0_6561 = (_zz_dataOut_payload_0_6560 ? _zz_dataOut_payload_0_6431 : _zz_dataOut_payload_0_6407);
  assign _zz_dataOut_payload_0_6562 = (_zz_dataOut_payload_0_6560 ? _zz_dataOut_payload_0_6407 : _zz_dataOut_payload_0_6431);
  assign _zz_dataOut_payload_0_6563 = (_zz_dataOut_payload_0_6428 < _zz_dataOut_payload_0_6404);
  assign _zz_dataOut_payload_0_6564 = (_zz_dataOut_payload_0_6563 ? _zz_dataOut_payload_0_6428 : _zz_dataOut_payload_0_6404);
  assign _zz_dataOut_payload_0_6565 = (_zz_dataOut_payload_0_6563 ? _zz_dataOut_payload_0_6404 : _zz_dataOut_payload_0_6428);
  assign _zz_dataOut_payload_0_6566 = (_zz_dataOut_payload_0_6425 < _zz_dataOut_payload_0_6401);
  assign _zz_dataOut_payload_0_6567 = (_zz_dataOut_payload_0_6566 ? _zz_dataOut_payload_0_6425 : _zz_dataOut_payload_0_6401);
  assign _zz_dataOut_payload_0_6568 = (_zz_dataOut_payload_0_6566 ? _zz_dataOut_payload_0_6401 : _zz_dataOut_payload_0_6425);
  assign _zz_dataOut_payload_0_6569 = (_zz_dataOut_payload_0_6422 < _zz_dataOut_payload_0_6398);
  assign _zz_dataOut_payload_0_6570 = (_zz_dataOut_payload_0_6569 ? _zz_dataOut_payload_0_6422 : _zz_dataOut_payload_0_6398);
  assign _zz_dataOut_payload_0_6571 = (_zz_dataOut_payload_0_6569 ? _zz_dataOut_payload_0_6398 : _zz_dataOut_payload_0_6422);
  assign _zz_dataOut_payload_0_6572 = (_zz_dataOut_payload_0_6419 < _zz_dataOut_payload_0_6395);
  assign _zz_dataOut_payload_0_6573 = (_zz_dataOut_payload_0_6572 ? _zz_dataOut_payload_0_6419 : _zz_dataOut_payload_0_6395);
  assign _zz_dataOut_payload_0_6574 = (_zz_dataOut_payload_0_6572 ? _zz_dataOut_payload_0_6395 : _zz_dataOut_payload_0_6419);
  assign _zz_dataOut_payload_0_6575 = (_zz_dataOut_payload_0_6416 < _zz_dataOut_payload_0_6392);
  assign _zz_dataOut_payload_0_6576 = (_zz_dataOut_payload_0_6575 ? _zz_dataOut_payload_0_6416 : _zz_dataOut_payload_0_6392);
  assign _zz_dataOut_payload_0_6577 = (_zz_dataOut_payload_0_6575 ? _zz_dataOut_payload_0_6392 : _zz_dataOut_payload_0_6416);
  assign _zz_dataOut_payload_0_6578 = (_zz_dataOut_payload_0_6413 < _zz_dataOut_payload_0_6389);
  assign _zz_dataOut_payload_0_6579 = (_zz_dataOut_payload_0_6578 ? _zz_dataOut_payload_0_6413 : _zz_dataOut_payload_0_6389);
  assign _zz_dataOut_payload_0_6580 = (_zz_dataOut_payload_0_6578 ? _zz_dataOut_payload_0_6389 : _zz_dataOut_payload_0_6413);
  assign _zz_dataOut_payload_0_6581 = (_zz_dataOut_payload_0_6410 < _zz_dataOut_payload_0_6386);
  assign _zz_dataOut_payload_0_6582 = (_zz_dataOut_payload_0_6581 ? _zz_dataOut_payload_0_6410 : _zz_dataOut_payload_0_6386);
  assign _zz_dataOut_payload_0_6583 = (_zz_dataOut_payload_0_6581 ? _zz_dataOut_payload_0_6386 : _zz_dataOut_payload_0_6410);
  assign _zz_dataOut_payload_0_6584 = (_zz_dataOut_payload_0_6561 < _zz_dataOut_payload_0_6573);
  assign _zz_dataOut_payload_0_6585 = (_zz_dataOut_payload_0_6584 ? _zz_dataOut_payload_0_6561 : _zz_dataOut_payload_0_6573);
  assign _zz_dataOut_payload_0_6586 = (_zz_dataOut_payload_0_6584 ? _zz_dataOut_payload_0_6573 : _zz_dataOut_payload_0_6561);
  assign _zz_dataOut_payload_0_6587 = (_zz_dataOut_payload_0_6564 < _zz_dataOut_payload_0_6576);
  assign _zz_dataOut_payload_0_6588 = (_zz_dataOut_payload_0_6587 ? _zz_dataOut_payload_0_6564 : _zz_dataOut_payload_0_6576);
  assign _zz_dataOut_payload_0_6589 = (_zz_dataOut_payload_0_6587 ? _zz_dataOut_payload_0_6576 : _zz_dataOut_payload_0_6564);
  assign _zz_dataOut_payload_0_6590 = (_zz_dataOut_payload_0_6567 < _zz_dataOut_payload_0_6579);
  assign _zz_dataOut_payload_0_6591 = (_zz_dataOut_payload_0_6590 ? _zz_dataOut_payload_0_6567 : _zz_dataOut_payload_0_6579);
  assign _zz_dataOut_payload_0_6592 = (_zz_dataOut_payload_0_6590 ? _zz_dataOut_payload_0_6579 : _zz_dataOut_payload_0_6567);
  assign _zz_dataOut_payload_0_6593 = (_zz_dataOut_payload_0_6570 < _zz_dataOut_payload_0_6582);
  assign _zz_dataOut_payload_0_6594 = (_zz_dataOut_payload_0_6593 ? _zz_dataOut_payload_0_6570 : _zz_dataOut_payload_0_6582);
  assign _zz_dataOut_payload_0_6595 = (_zz_dataOut_payload_0_6593 ? _zz_dataOut_payload_0_6582 : _zz_dataOut_payload_0_6570);
  assign _zz_dataOut_payload_0_6596 = (_zz_dataOut_payload_0_6585 < _zz_dataOut_payload_0_6591);
  assign _zz_dataOut_payload_0_6597 = (_zz_dataOut_payload_0_6596 ? _zz_dataOut_payload_0_6585 : _zz_dataOut_payload_0_6591);
  assign _zz_dataOut_payload_0_6598 = (_zz_dataOut_payload_0_6596 ? _zz_dataOut_payload_0_6591 : _zz_dataOut_payload_0_6585);
  assign _zz_dataOut_payload_0_6599 = (_zz_dataOut_payload_0_6588 < _zz_dataOut_payload_0_6594);
  assign _zz_dataOut_payload_0_6600 = (_zz_dataOut_payload_0_6599 ? _zz_dataOut_payload_0_6588 : _zz_dataOut_payload_0_6594);
  assign _zz_dataOut_payload_0_6601 = (_zz_dataOut_payload_0_6599 ? _zz_dataOut_payload_0_6594 : _zz_dataOut_payload_0_6588);
  assign _zz_dataOut_payload_0_6602 = (_zz_dataOut_payload_0_6597 < _zz_dataOut_payload_0_6600);
  assign _zz_dataOut_payload_0_6603 = (_zz_dataOut_payload_0_6598 < _zz_dataOut_payload_0_6601);
  assign _zz_dataOut_payload_0_6608 = (_zz_dataOut_payload_0_6586 < _zz_dataOut_payload_0_6592);
  assign _zz_dataOut_payload_0_6609 = (_zz_dataOut_payload_0_6608 ? _zz_dataOut_payload_0_6586 : _zz_dataOut_payload_0_6592);
  assign _zz_dataOut_payload_0_6610 = (_zz_dataOut_payload_0_6608 ? _zz_dataOut_payload_0_6592 : _zz_dataOut_payload_0_6586);
  assign _zz_dataOut_payload_0_6611 = (_zz_dataOut_payload_0_6589 < _zz_dataOut_payload_0_6595);
  assign _zz_dataOut_payload_0_6612 = (_zz_dataOut_payload_0_6611 ? _zz_dataOut_payload_0_6589 : _zz_dataOut_payload_0_6595);
  assign _zz_dataOut_payload_0_6613 = (_zz_dataOut_payload_0_6611 ? _zz_dataOut_payload_0_6595 : _zz_dataOut_payload_0_6589);
  assign _zz_dataOut_payload_0_6614 = (_zz_dataOut_payload_0_6609 < _zz_dataOut_payload_0_6612);
  assign _zz_dataOut_payload_0_6615 = (_zz_dataOut_payload_0_6610 < _zz_dataOut_payload_0_6613);
  assign _zz_dataOut_payload_0_6628 = (_zz_dataOut_payload_0_6562 < _zz_dataOut_payload_0_6574);
  assign _zz_dataOut_payload_0_6629 = (_zz_dataOut_payload_0_6628 ? _zz_dataOut_payload_0_6562 : _zz_dataOut_payload_0_6574);
  assign _zz_dataOut_payload_0_6630 = (_zz_dataOut_payload_0_6628 ? _zz_dataOut_payload_0_6574 : _zz_dataOut_payload_0_6562);
  assign _zz_dataOut_payload_0_6631 = (_zz_dataOut_payload_0_6565 < _zz_dataOut_payload_0_6577);
  assign _zz_dataOut_payload_0_6632 = (_zz_dataOut_payload_0_6631 ? _zz_dataOut_payload_0_6565 : _zz_dataOut_payload_0_6577);
  assign _zz_dataOut_payload_0_6633 = (_zz_dataOut_payload_0_6631 ? _zz_dataOut_payload_0_6577 : _zz_dataOut_payload_0_6565);
  assign _zz_dataOut_payload_0_6634 = (_zz_dataOut_payload_0_6568 < _zz_dataOut_payload_0_6580);
  assign _zz_dataOut_payload_0_6635 = (_zz_dataOut_payload_0_6634 ? _zz_dataOut_payload_0_6568 : _zz_dataOut_payload_0_6580);
  assign _zz_dataOut_payload_0_6636 = (_zz_dataOut_payload_0_6634 ? _zz_dataOut_payload_0_6580 : _zz_dataOut_payload_0_6568);
  assign _zz_dataOut_payload_0_6637 = (_zz_dataOut_payload_0_6571 < _zz_dataOut_payload_0_6583);
  assign _zz_dataOut_payload_0_6638 = (_zz_dataOut_payload_0_6637 ? _zz_dataOut_payload_0_6571 : _zz_dataOut_payload_0_6583);
  assign _zz_dataOut_payload_0_6639 = (_zz_dataOut_payload_0_6637 ? _zz_dataOut_payload_0_6583 : _zz_dataOut_payload_0_6571);
  assign _zz_dataOut_payload_0_6640 = (_zz_dataOut_payload_0_6629 < _zz_dataOut_payload_0_6635);
  assign _zz_dataOut_payload_0_6641 = (_zz_dataOut_payload_0_6640 ? _zz_dataOut_payload_0_6629 : _zz_dataOut_payload_0_6635);
  assign _zz_dataOut_payload_0_6642 = (_zz_dataOut_payload_0_6640 ? _zz_dataOut_payload_0_6635 : _zz_dataOut_payload_0_6629);
  assign _zz_dataOut_payload_0_6643 = (_zz_dataOut_payload_0_6632 < _zz_dataOut_payload_0_6638);
  assign _zz_dataOut_payload_0_6644 = (_zz_dataOut_payload_0_6643 ? _zz_dataOut_payload_0_6632 : _zz_dataOut_payload_0_6638);
  assign _zz_dataOut_payload_0_6645 = (_zz_dataOut_payload_0_6643 ? _zz_dataOut_payload_0_6638 : _zz_dataOut_payload_0_6632);
  assign _zz_dataOut_payload_0_6646 = (_zz_dataOut_payload_0_6641 < _zz_dataOut_payload_0_6644);
  assign _zz_dataOut_payload_0_6647 = (_zz_dataOut_payload_0_6642 < _zz_dataOut_payload_0_6645);
  assign _zz_dataOut_payload_0_6652 = (_zz_dataOut_payload_0_6630 < _zz_dataOut_payload_0_6636);
  assign _zz_dataOut_payload_0_6653 = (_zz_dataOut_payload_0_6652 ? _zz_dataOut_payload_0_6630 : _zz_dataOut_payload_0_6636);
  assign _zz_dataOut_payload_0_6654 = (_zz_dataOut_payload_0_6652 ? _zz_dataOut_payload_0_6636 : _zz_dataOut_payload_0_6630);
  assign _zz_dataOut_payload_0_6655 = (_zz_dataOut_payload_0_6633 < _zz_dataOut_payload_0_6639);
  assign _zz_dataOut_payload_0_6656 = (_zz_dataOut_payload_0_6655 ? _zz_dataOut_payload_0_6633 : _zz_dataOut_payload_0_6639);
  assign _zz_dataOut_payload_0_6657 = (_zz_dataOut_payload_0_6655 ? _zz_dataOut_payload_0_6639 : _zz_dataOut_payload_0_6633);
  assign _zz_dataOut_payload_0_6658 = (_zz_dataOut_payload_0_6653 < _zz_dataOut_payload_0_6656);
  assign _zz_dataOut_payload_0_6659 = (_zz_dataOut_payload_0_6654 < _zz_dataOut_payload_0_6657);
  assign _zz_dataOut_payload_0_6720 = (_zz_dataOut_payload_0_5248 < _zz_dataOut_payload_0_5279);
  assign _zz_dataOut_payload_0_6721 = (_zz_dataOut_payload_0_6720 ? _zz_dataOut_payload_0_5248 : _zz_dataOut_payload_0_5279);
  assign _zz_dataOut_payload_0_6722 = (_zz_dataOut_payload_0_6720 ? _zz_dataOut_payload_0_5279 : _zz_dataOut_payload_0_5248);
  assign _zz_dataOut_payload_0_6723 = (_zz_dataOut_payload_0_5249 < _zz_dataOut_payload_0_5278);
  assign _zz_dataOut_payload_0_6724 = (_zz_dataOut_payload_0_6723 ? _zz_dataOut_payload_0_5249 : _zz_dataOut_payload_0_5278);
  assign _zz_dataOut_payload_0_6725 = (_zz_dataOut_payload_0_6723 ? _zz_dataOut_payload_0_5278 : _zz_dataOut_payload_0_5249);
  assign _zz_dataOut_payload_0_6726 = (_zz_dataOut_payload_0_5250 < _zz_dataOut_payload_0_5277);
  assign _zz_dataOut_payload_0_6727 = (_zz_dataOut_payload_0_6726 ? _zz_dataOut_payload_0_5250 : _zz_dataOut_payload_0_5277);
  assign _zz_dataOut_payload_0_6728 = (_zz_dataOut_payload_0_6726 ? _zz_dataOut_payload_0_5277 : _zz_dataOut_payload_0_5250);
  assign _zz_dataOut_payload_0_6729 = (_zz_dataOut_payload_0_5251 < _zz_dataOut_payload_0_5276);
  assign _zz_dataOut_payload_0_6730 = (_zz_dataOut_payload_0_6729 ? _zz_dataOut_payload_0_5251 : _zz_dataOut_payload_0_5276);
  assign _zz_dataOut_payload_0_6731 = (_zz_dataOut_payload_0_6729 ? _zz_dataOut_payload_0_5276 : _zz_dataOut_payload_0_5251);
  assign _zz_dataOut_payload_0_6732 = (_zz_dataOut_payload_0_5252 < _zz_dataOut_payload_0_5275);
  assign _zz_dataOut_payload_0_6733 = (_zz_dataOut_payload_0_6732 ? _zz_dataOut_payload_0_5252 : _zz_dataOut_payload_0_5275);
  assign _zz_dataOut_payload_0_6734 = (_zz_dataOut_payload_0_6732 ? _zz_dataOut_payload_0_5275 : _zz_dataOut_payload_0_5252);
  assign _zz_dataOut_payload_0_6735 = (_zz_dataOut_payload_0_5253 < _zz_dataOut_payload_0_5274);
  assign _zz_dataOut_payload_0_6736 = (_zz_dataOut_payload_0_6735 ? _zz_dataOut_payload_0_5253 : _zz_dataOut_payload_0_5274);
  assign _zz_dataOut_payload_0_6737 = (_zz_dataOut_payload_0_6735 ? _zz_dataOut_payload_0_5274 : _zz_dataOut_payload_0_5253);
  assign _zz_dataOut_payload_0_6738 = (_zz_dataOut_payload_0_5254 < _zz_dataOut_payload_0_5273);
  assign _zz_dataOut_payload_0_6739 = (_zz_dataOut_payload_0_6738 ? _zz_dataOut_payload_0_5254 : _zz_dataOut_payload_0_5273);
  assign _zz_dataOut_payload_0_6740 = (_zz_dataOut_payload_0_6738 ? _zz_dataOut_payload_0_5273 : _zz_dataOut_payload_0_5254);
  assign _zz_dataOut_payload_0_6741 = (_zz_dataOut_payload_0_5255 < _zz_dataOut_payload_0_5272);
  assign _zz_dataOut_payload_0_6742 = (_zz_dataOut_payload_0_6741 ? _zz_dataOut_payload_0_5255 : _zz_dataOut_payload_0_5272);
  assign _zz_dataOut_payload_0_6743 = (_zz_dataOut_payload_0_6741 ? _zz_dataOut_payload_0_5272 : _zz_dataOut_payload_0_5255);
  assign _zz_dataOut_payload_0_6744 = (_zz_dataOut_payload_0_5256 < _zz_dataOut_payload_0_5271);
  assign _zz_dataOut_payload_0_6745 = (_zz_dataOut_payload_0_6744 ? _zz_dataOut_payload_0_5256 : _zz_dataOut_payload_0_5271);
  assign _zz_dataOut_payload_0_6746 = (_zz_dataOut_payload_0_6744 ? _zz_dataOut_payload_0_5271 : _zz_dataOut_payload_0_5256);
  assign _zz_dataOut_payload_0_6747 = (_zz_dataOut_payload_0_5257 < _zz_dataOut_payload_0_5270);
  assign _zz_dataOut_payload_0_6748 = (_zz_dataOut_payload_0_6747 ? _zz_dataOut_payload_0_5257 : _zz_dataOut_payload_0_5270);
  assign _zz_dataOut_payload_0_6749 = (_zz_dataOut_payload_0_6747 ? _zz_dataOut_payload_0_5270 : _zz_dataOut_payload_0_5257);
  assign _zz_dataOut_payload_0_6750 = (_zz_dataOut_payload_0_5258 < _zz_dataOut_payload_0_5269);
  assign _zz_dataOut_payload_0_6751 = (_zz_dataOut_payload_0_6750 ? _zz_dataOut_payload_0_5258 : _zz_dataOut_payload_0_5269);
  assign _zz_dataOut_payload_0_6752 = (_zz_dataOut_payload_0_6750 ? _zz_dataOut_payload_0_5269 : _zz_dataOut_payload_0_5258);
  assign _zz_dataOut_payload_0_6753 = (_zz_dataOut_payload_0_5259 < _zz_dataOut_payload_0_5268);
  assign _zz_dataOut_payload_0_6754 = (_zz_dataOut_payload_0_6753 ? _zz_dataOut_payload_0_5259 : _zz_dataOut_payload_0_5268);
  assign _zz_dataOut_payload_0_6755 = (_zz_dataOut_payload_0_6753 ? _zz_dataOut_payload_0_5268 : _zz_dataOut_payload_0_5259);
  assign _zz_dataOut_payload_0_6756 = (_zz_dataOut_payload_0_5260 < _zz_dataOut_payload_0_5267);
  assign _zz_dataOut_payload_0_6757 = (_zz_dataOut_payload_0_6756 ? _zz_dataOut_payload_0_5260 : _zz_dataOut_payload_0_5267);
  assign _zz_dataOut_payload_0_6758 = (_zz_dataOut_payload_0_6756 ? _zz_dataOut_payload_0_5267 : _zz_dataOut_payload_0_5260);
  assign _zz_dataOut_payload_0_6759 = (_zz_dataOut_payload_0_5261 < _zz_dataOut_payload_0_5266);
  assign _zz_dataOut_payload_0_6760 = (_zz_dataOut_payload_0_6759 ? _zz_dataOut_payload_0_5261 : _zz_dataOut_payload_0_5266);
  assign _zz_dataOut_payload_0_6761 = (_zz_dataOut_payload_0_6759 ? _zz_dataOut_payload_0_5266 : _zz_dataOut_payload_0_5261);
  assign _zz_dataOut_payload_0_6762 = (_zz_dataOut_payload_0_5262 < _zz_dataOut_payload_0_5265);
  assign _zz_dataOut_payload_0_6763 = (_zz_dataOut_payload_0_6762 ? _zz_dataOut_payload_0_5262 : _zz_dataOut_payload_0_5265);
  assign _zz_dataOut_payload_0_6764 = (_zz_dataOut_payload_0_6762 ? _zz_dataOut_payload_0_5265 : _zz_dataOut_payload_0_5262);
  assign _zz_dataOut_payload_0_6765 = (_zz_dataOut_payload_0_5263 < _zz_dataOut_payload_0_5264);
  assign _zz_dataOut_payload_0_6766 = (_zz_dataOut_payload_0_6765 ? _zz_dataOut_payload_0_5263 : _zz_dataOut_payload_0_5264);
  assign _zz_dataOut_payload_0_6767 = (_zz_dataOut_payload_0_6765 ? _zz_dataOut_payload_0_5264 : _zz_dataOut_payload_0_5263);
  assign _zz_dataOut_payload_0_6768 = (_zz_dataOut_payload_0_6721 < _zz_dataOut_payload_0_6745);
  assign _zz_dataOut_payload_0_6769 = (_zz_dataOut_payload_0_6768 ? _zz_dataOut_payload_0_6721 : _zz_dataOut_payload_0_6745);
  assign _zz_dataOut_payload_0_6770 = (_zz_dataOut_payload_0_6768 ? _zz_dataOut_payload_0_6745 : _zz_dataOut_payload_0_6721);
  assign _zz_dataOut_payload_0_6771 = (_zz_dataOut_payload_0_6724 < _zz_dataOut_payload_0_6748);
  assign _zz_dataOut_payload_0_6772 = (_zz_dataOut_payload_0_6771 ? _zz_dataOut_payload_0_6724 : _zz_dataOut_payload_0_6748);
  assign _zz_dataOut_payload_0_6773 = (_zz_dataOut_payload_0_6771 ? _zz_dataOut_payload_0_6748 : _zz_dataOut_payload_0_6724);
  assign _zz_dataOut_payload_0_6774 = (_zz_dataOut_payload_0_6727 < _zz_dataOut_payload_0_6751);
  assign _zz_dataOut_payload_0_6775 = (_zz_dataOut_payload_0_6774 ? _zz_dataOut_payload_0_6727 : _zz_dataOut_payload_0_6751);
  assign _zz_dataOut_payload_0_6776 = (_zz_dataOut_payload_0_6774 ? _zz_dataOut_payload_0_6751 : _zz_dataOut_payload_0_6727);
  assign _zz_dataOut_payload_0_6777 = (_zz_dataOut_payload_0_6730 < _zz_dataOut_payload_0_6754);
  assign _zz_dataOut_payload_0_6778 = (_zz_dataOut_payload_0_6777 ? _zz_dataOut_payload_0_6730 : _zz_dataOut_payload_0_6754);
  assign _zz_dataOut_payload_0_6779 = (_zz_dataOut_payload_0_6777 ? _zz_dataOut_payload_0_6754 : _zz_dataOut_payload_0_6730);
  assign _zz_dataOut_payload_0_6780 = (_zz_dataOut_payload_0_6733 < _zz_dataOut_payload_0_6757);
  assign _zz_dataOut_payload_0_6781 = (_zz_dataOut_payload_0_6780 ? _zz_dataOut_payload_0_6733 : _zz_dataOut_payload_0_6757);
  assign _zz_dataOut_payload_0_6782 = (_zz_dataOut_payload_0_6780 ? _zz_dataOut_payload_0_6757 : _zz_dataOut_payload_0_6733);
  assign _zz_dataOut_payload_0_6783 = (_zz_dataOut_payload_0_6736 < _zz_dataOut_payload_0_6760);
  assign _zz_dataOut_payload_0_6784 = (_zz_dataOut_payload_0_6783 ? _zz_dataOut_payload_0_6736 : _zz_dataOut_payload_0_6760);
  assign _zz_dataOut_payload_0_6785 = (_zz_dataOut_payload_0_6783 ? _zz_dataOut_payload_0_6760 : _zz_dataOut_payload_0_6736);
  assign _zz_dataOut_payload_0_6786 = (_zz_dataOut_payload_0_6739 < _zz_dataOut_payload_0_6763);
  assign _zz_dataOut_payload_0_6787 = (_zz_dataOut_payload_0_6786 ? _zz_dataOut_payload_0_6739 : _zz_dataOut_payload_0_6763);
  assign _zz_dataOut_payload_0_6788 = (_zz_dataOut_payload_0_6786 ? _zz_dataOut_payload_0_6763 : _zz_dataOut_payload_0_6739);
  assign _zz_dataOut_payload_0_6789 = (_zz_dataOut_payload_0_6742 < _zz_dataOut_payload_0_6766);
  assign _zz_dataOut_payload_0_6790 = (_zz_dataOut_payload_0_6789 ? _zz_dataOut_payload_0_6742 : _zz_dataOut_payload_0_6766);
  assign _zz_dataOut_payload_0_6791 = (_zz_dataOut_payload_0_6789 ? _zz_dataOut_payload_0_6766 : _zz_dataOut_payload_0_6742);
  assign _zz_dataOut_payload_0_6792 = (_zz_dataOut_payload_0_6769 < _zz_dataOut_payload_0_6781);
  assign _zz_dataOut_payload_0_6793 = (_zz_dataOut_payload_0_6792 ? _zz_dataOut_payload_0_6769 : _zz_dataOut_payload_0_6781);
  assign _zz_dataOut_payload_0_6794 = (_zz_dataOut_payload_0_6792 ? _zz_dataOut_payload_0_6781 : _zz_dataOut_payload_0_6769);
  assign _zz_dataOut_payload_0_6795 = (_zz_dataOut_payload_0_6772 < _zz_dataOut_payload_0_6784);
  assign _zz_dataOut_payload_0_6796 = (_zz_dataOut_payload_0_6795 ? _zz_dataOut_payload_0_6772 : _zz_dataOut_payload_0_6784);
  assign _zz_dataOut_payload_0_6797 = (_zz_dataOut_payload_0_6795 ? _zz_dataOut_payload_0_6784 : _zz_dataOut_payload_0_6772);
  assign _zz_dataOut_payload_0_6798 = (_zz_dataOut_payload_0_6775 < _zz_dataOut_payload_0_6787);
  assign _zz_dataOut_payload_0_6799 = (_zz_dataOut_payload_0_6798 ? _zz_dataOut_payload_0_6775 : _zz_dataOut_payload_0_6787);
  assign _zz_dataOut_payload_0_6800 = (_zz_dataOut_payload_0_6798 ? _zz_dataOut_payload_0_6787 : _zz_dataOut_payload_0_6775);
  assign _zz_dataOut_payload_0_6801 = (_zz_dataOut_payload_0_6778 < _zz_dataOut_payload_0_6790);
  assign _zz_dataOut_payload_0_6802 = (_zz_dataOut_payload_0_6801 ? _zz_dataOut_payload_0_6778 : _zz_dataOut_payload_0_6790);
  assign _zz_dataOut_payload_0_6803 = (_zz_dataOut_payload_0_6801 ? _zz_dataOut_payload_0_6790 : _zz_dataOut_payload_0_6778);
  assign _zz_dataOut_payload_0_6804 = (_zz_dataOut_payload_0_6793 < _zz_dataOut_payload_0_6799);
  assign _zz_dataOut_payload_0_6805 = (_zz_dataOut_payload_0_6804 ? _zz_dataOut_payload_0_6793 : _zz_dataOut_payload_0_6799);
  assign _zz_dataOut_payload_0_6806 = (_zz_dataOut_payload_0_6804 ? _zz_dataOut_payload_0_6799 : _zz_dataOut_payload_0_6793);
  assign _zz_dataOut_payload_0_6807 = (_zz_dataOut_payload_0_6796 < _zz_dataOut_payload_0_6802);
  assign _zz_dataOut_payload_0_6808 = (_zz_dataOut_payload_0_6807 ? _zz_dataOut_payload_0_6796 : _zz_dataOut_payload_0_6802);
  assign _zz_dataOut_payload_0_6809 = (_zz_dataOut_payload_0_6807 ? _zz_dataOut_payload_0_6802 : _zz_dataOut_payload_0_6796);
  assign _zz_dataOut_payload_0_6810 = (_zz_dataOut_payload_0_6805 < _zz_dataOut_payload_0_6808);
  assign _zz_dataOut_payload_0_6811 = (_zz_dataOut_payload_0_6806 < _zz_dataOut_payload_0_6809);
  assign _zz_dataOut_payload_0_6816 = (_zz_dataOut_payload_0_6794 < _zz_dataOut_payload_0_6800);
  assign _zz_dataOut_payload_0_6817 = (_zz_dataOut_payload_0_6816 ? _zz_dataOut_payload_0_6794 : _zz_dataOut_payload_0_6800);
  assign _zz_dataOut_payload_0_6818 = (_zz_dataOut_payload_0_6816 ? _zz_dataOut_payload_0_6800 : _zz_dataOut_payload_0_6794);
  assign _zz_dataOut_payload_0_6819 = (_zz_dataOut_payload_0_6797 < _zz_dataOut_payload_0_6803);
  assign _zz_dataOut_payload_0_6820 = (_zz_dataOut_payload_0_6819 ? _zz_dataOut_payload_0_6797 : _zz_dataOut_payload_0_6803);
  assign _zz_dataOut_payload_0_6821 = (_zz_dataOut_payload_0_6819 ? _zz_dataOut_payload_0_6803 : _zz_dataOut_payload_0_6797);
  assign _zz_dataOut_payload_0_6822 = (_zz_dataOut_payload_0_6817 < _zz_dataOut_payload_0_6820);
  assign _zz_dataOut_payload_0_6823 = (_zz_dataOut_payload_0_6818 < _zz_dataOut_payload_0_6821);
  assign _zz_dataOut_payload_0_6836 = (_zz_dataOut_payload_0_6770 < _zz_dataOut_payload_0_6782);
  assign _zz_dataOut_payload_0_6837 = (_zz_dataOut_payload_0_6836 ? _zz_dataOut_payload_0_6770 : _zz_dataOut_payload_0_6782);
  assign _zz_dataOut_payload_0_6838 = (_zz_dataOut_payload_0_6836 ? _zz_dataOut_payload_0_6782 : _zz_dataOut_payload_0_6770);
  assign _zz_dataOut_payload_0_6839 = (_zz_dataOut_payload_0_6773 < _zz_dataOut_payload_0_6785);
  assign _zz_dataOut_payload_0_6840 = (_zz_dataOut_payload_0_6839 ? _zz_dataOut_payload_0_6773 : _zz_dataOut_payload_0_6785);
  assign _zz_dataOut_payload_0_6841 = (_zz_dataOut_payload_0_6839 ? _zz_dataOut_payload_0_6785 : _zz_dataOut_payload_0_6773);
  assign _zz_dataOut_payload_0_6842 = (_zz_dataOut_payload_0_6776 < _zz_dataOut_payload_0_6788);
  assign _zz_dataOut_payload_0_6843 = (_zz_dataOut_payload_0_6842 ? _zz_dataOut_payload_0_6776 : _zz_dataOut_payload_0_6788);
  assign _zz_dataOut_payload_0_6844 = (_zz_dataOut_payload_0_6842 ? _zz_dataOut_payload_0_6788 : _zz_dataOut_payload_0_6776);
  assign _zz_dataOut_payload_0_6845 = (_zz_dataOut_payload_0_6779 < _zz_dataOut_payload_0_6791);
  assign _zz_dataOut_payload_0_6846 = (_zz_dataOut_payload_0_6845 ? _zz_dataOut_payload_0_6779 : _zz_dataOut_payload_0_6791);
  assign _zz_dataOut_payload_0_6847 = (_zz_dataOut_payload_0_6845 ? _zz_dataOut_payload_0_6791 : _zz_dataOut_payload_0_6779);
  assign _zz_dataOut_payload_0_6848 = (_zz_dataOut_payload_0_6837 < _zz_dataOut_payload_0_6843);
  assign _zz_dataOut_payload_0_6849 = (_zz_dataOut_payload_0_6848 ? _zz_dataOut_payload_0_6837 : _zz_dataOut_payload_0_6843);
  assign _zz_dataOut_payload_0_6850 = (_zz_dataOut_payload_0_6848 ? _zz_dataOut_payload_0_6843 : _zz_dataOut_payload_0_6837);
  assign _zz_dataOut_payload_0_6851 = (_zz_dataOut_payload_0_6840 < _zz_dataOut_payload_0_6846);
  assign _zz_dataOut_payload_0_6852 = (_zz_dataOut_payload_0_6851 ? _zz_dataOut_payload_0_6840 : _zz_dataOut_payload_0_6846);
  assign _zz_dataOut_payload_0_6853 = (_zz_dataOut_payload_0_6851 ? _zz_dataOut_payload_0_6846 : _zz_dataOut_payload_0_6840);
  assign _zz_dataOut_payload_0_6854 = (_zz_dataOut_payload_0_6849 < _zz_dataOut_payload_0_6852);
  assign _zz_dataOut_payload_0_6855 = (_zz_dataOut_payload_0_6850 < _zz_dataOut_payload_0_6853);
  assign _zz_dataOut_payload_0_6860 = (_zz_dataOut_payload_0_6838 < _zz_dataOut_payload_0_6844);
  assign _zz_dataOut_payload_0_6861 = (_zz_dataOut_payload_0_6860 ? _zz_dataOut_payload_0_6838 : _zz_dataOut_payload_0_6844);
  assign _zz_dataOut_payload_0_6862 = (_zz_dataOut_payload_0_6860 ? _zz_dataOut_payload_0_6844 : _zz_dataOut_payload_0_6838);
  assign _zz_dataOut_payload_0_6863 = (_zz_dataOut_payload_0_6841 < _zz_dataOut_payload_0_6847);
  assign _zz_dataOut_payload_0_6864 = (_zz_dataOut_payload_0_6863 ? _zz_dataOut_payload_0_6841 : _zz_dataOut_payload_0_6847);
  assign _zz_dataOut_payload_0_6865 = (_zz_dataOut_payload_0_6863 ? _zz_dataOut_payload_0_6847 : _zz_dataOut_payload_0_6841);
  assign _zz_dataOut_payload_0_6866 = (_zz_dataOut_payload_0_6861 < _zz_dataOut_payload_0_6864);
  assign _zz_dataOut_payload_0_6867 = (_zz_dataOut_payload_0_6862 < _zz_dataOut_payload_0_6865);
  assign _zz_dataOut_payload_0_6896 = (_zz_dataOut_payload_0_6767 < _zz_dataOut_payload_0_6743);
  assign _zz_dataOut_payload_0_6897 = (_zz_dataOut_payload_0_6896 ? _zz_dataOut_payload_0_6767 : _zz_dataOut_payload_0_6743);
  assign _zz_dataOut_payload_0_6898 = (_zz_dataOut_payload_0_6896 ? _zz_dataOut_payload_0_6743 : _zz_dataOut_payload_0_6767);
  assign _zz_dataOut_payload_0_6899 = (_zz_dataOut_payload_0_6764 < _zz_dataOut_payload_0_6740);
  assign _zz_dataOut_payload_0_6900 = (_zz_dataOut_payload_0_6899 ? _zz_dataOut_payload_0_6764 : _zz_dataOut_payload_0_6740);
  assign _zz_dataOut_payload_0_6901 = (_zz_dataOut_payload_0_6899 ? _zz_dataOut_payload_0_6740 : _zz_dataOut_payload_0_6764);
  assign _zz_dataOut_payload_0_6902 = (_zz_dataOut_payload_0_6761 < _zz_dataOut_payload_0_6737);
  assign _zz_dataOut_payload_0_6903 = (_zz_dataOut_payload_0_6902 ? _zz_dataOut_payload_0_6761 : _zz_dataOut_payload_0_6737);
  assign _zz_dataOut_payload_0_6904 = (_zz_dataOut_payload_0_6902 ? _zz_dataOut_payload_0_6737 : _zz_dataOut_payload_0_6761);
  assign _zz_dataOut_payload_0_6905 = (_zz_dataOut_payload_0_6758 < _zz_dataOut_payload_0_6734);
  assign _zz_dataOut_payload_0_6906 = (_zz_dataOut_payload_0_6905 ? _zz_dataOut_payload_0_6758 : _zz_dataOut_payload_0_6734);
  assign _zz_dataOut_payload_0_6907 = (_zz_dataOut_payload_0_6905 ? _zz_dataOut_payload_0_6734 : _zz_dataOut_payload_0_6758);
  assign _zz_dataOut_payload_0_6908 = (_zz_dataOut_payload_0_6755 < _zz_dataOut_payload_0_6731);
  assign _zz_dataOut_payload_0_6909 = (_zz_dataOut_payload_0_6908 ? _zz_dataOut_payload_0_6755 : _zz_dataOut_payload_0_6731);
  assign _zz_dataOut_payload_0_6910 = (_zz_dataOut_payload_0_6908 ? _zz_dataOut_payload_0_6731 : _zz_dataOut_payload_0_6755);
  assign _zz_dataOut_payload_0_6911 = (_zz_dataOut_payload_0_6752 < _zz_dataOut_payload_0_6728);
  assign _zz_dataOut_payload_0_6912 = (_zz_dataOut_payload_0_6911 ? _zz_dataOut_payload_0_6752 : _zz_dataOut_payload_0_6728);
  assign _zz_dataOut_payload_0_6913 = (_zz_dataOut_payload_0_6911 ? _zz_dataOut_payload_0_6728 : _zz_dataOut_payload_0_6752);
  assign _zz_dataOut_payload_0_6914 = (_zz_dataOut_payload_0_6749 < _zz_dataOut_payload_0_6725);
  assign _zz_dataOut_payload_0_6915 = (_zz_dataOut_payload_0_6914 ? _zz_dataOut_payload_0_6749 : _zz_dataOut_payload_0_6725);
  assign _zz_dataOut_payload_0_6916 = (_zz_dataOut_payload_0_6914 ? _zz_dataOut_payload_0_6725 : _zz_dataOut_payload_0_6749);
  assign _zz_dataOut_payload_0_6917 = (_zz_dataOut_payload_0_6746 < _zz_dataOut_payload_0_6722);
  assign _zz_dataOut_payload_0_6918 = (_zz_dataOut_payload_0_6917 ? _zz_dataOut_payload_0_6746 : _zz_dataOut_payload_0_6722);
  assign _zz_dataOut_payload_0_6919 = (_zz_dataOut_payload_0_6917 ? _zz_dataOut_payload_0_6722 : _zz_dataOut_payload_0_6746);
  assign _zz_dataOut_payload_0_6920 = (_zz_dataOut_payload_0_6897 < _zz_dataOut_payload_0_6909);
  assign _zz_dataOut_payload_0_6921 = (_zz_dataOut_payload_0_6920 ? _zz_dataOut_payload_0_6897 : _zz_dataOut_payload_0_6909);
  assign _zz_dataOut_payload_0_6922 = (_zz_dataOut_payload_0_6920 ? _zz_dataOut_payload_0_6909 : _zz_dataOut_payload_0_6897);
  assign _zz_dataOut_payload_0_6923 = (_zz_dataOut_payload_0_6900 < _zz_dataOut_payload_0_6912);
  assign _zz_dataOut_payload_0_6924 = (_zz_dataOut_payload_0_6923 ? _zz_dataOut_payload_0_6900 : _zz_dataOut_payload_0_6912);
  assign _zz_dataOut_payload_0_6925 = (_zz_dataOut_payload_0_6923 ? _zz_dataOut_payload_0_6912 : _zz_dataOut_payload_0_6900);
  assign _zz_dataOut_payload_0_6926 = (_zz_dataOut_payload_0_6903 < _zz_dataOut_payload_0_6915);
  assign _zz_dataOut_payload_0_6927 = (_zz_dataOut_payload_0_6926 ? _zz_dataOut_payload_0_6903 : _zz_dataOut_payload_0_6915);
  assign _zz_dataOut_payload_0_6928 = (_zz_dataOut_payload_0_6926 ? _zz_dataOut_payload_0_6915 : _zz_dataOut_payload_0_6903);
  assign _zz_dataOut_payload_0_6929 = (_zz_dataOut_payload_0_6906 < _zz_dataOut_payload_0_6918);
  assign _zz_dataOut_payload_0_6930 = (_zz_dataOut_payload_0_6929 ? _zz_dataOut_payload_0_6906 : _zz_dataOut_payload_0_6918);
  assign _zz_dataOut_payload_0_6931 = (_zz_dataOut_payload_0_6929 ? _zz_dataOut_payload_0_6918 : _zz_dataOut_payload_0_6906);
  assign _zz_dataOut_payload_0_6932 = (_zz_dataOut_payload_0_6921 < _zz_dataOut_payload_0_6927);
  assign _zz_dataOut_payload_0_6933 = (_zz_dataOut_payload_0_6932 ? _zz_dataOut_payload_0_6921 : _zz_dataOut_payload_0_6927);
  assign _zz_dataOut_payload_0_6934 = (_zz_dataOut_payload_0_6932 ? _zz_dataOut_payload_0_6927 : _zz_dataOut_payload_0_6921);
  assign _zz_dataOut_payload_0_6935 = (_zz_dataOut_payload_0_6924 < _zz_dataOut_payload_0_6930);
  assign _zz_dataOut_payload_0_6936 = (_zz_dataOut_payload_0_6935 ? _zz_dataOut_payload_0_6924 : _zz_dataOut_payload_0_6930);
  assign _zz_dataOut_payload_0_6937 = (_zz_dataOut_payload_0_6935 ? _zz_dataOut_payload_0_6930 : _zz_dataOut_payload_0_6924);
  assign _zz_dataOut_payload_0_6938 = (_zz_dataOut_payload_0_6933 < _zz_dataOut_payload_0_6936);
  assign _zz_dataOut_payload_0_6939 = (_zz_dataOut_payload_0_6934 < _zz_dataOut_payload_0_6937);
  assign _zz_dataOut_payload_0_6944 = (_zz_dataOut_payload_0_6922 < _zz_dataOut_payload_0_6928);
  assign _zz_dataOut_payload_0_6945 = (_zz_dataOut_payload_0_6944 ? _zz_dataOut_payload_0_6922 : _zz_dataOut_payload_0_6928);
  assign _zz_dataOut_payload_0_6946 = (_zz_dataOut_payload_0_6944 ? _zz_dataOut_payload_0_6928 : _zz_dataOut_payload_0_6922);
  assign _zz_dataOut_payload_0_6947 = (_zz_dataOut_payload_0_6925 < _zz_dataOut_payload_0_6931);
  assign _zz_dataOut_payload_0_6948 = (_zz_dataOut_payload_0_6947 ? _zz_dataOut_payload_0_6925 : _zz_dataOut_payload_0_6931);
  assign _zz_dataOut_payload_0_6949 = (_zz_dataOut_payload_0_6947 ? _zz_dataOut_payload_0_6931 : _zz_dataOut_payload_0_6925);
  assign _zz_dataOut_payload_0_6950 = (_zz_dataOut_payload_0_6945 < _zz_dataOut_payload_0_6948);
  assign _zz_dataOut_payload_0_6951 = (_zz_dataOut_payload_0_6946 < _zz_dataOut_payload_0_6949);
  assign _zz_dataOut_payload_0_6964 = (_zz_dataOut_payload_0_6898 < _zz_dataOut_payload_0_6910);
  assign _zz_dataOut_payload_0_6965 = (_zz_dataOut_payload_0_6964 ? _zz_dataOut_payload_0_6898 : _zz_dataOut_payload_0_6910);
  assign _zz_dataOut_payload_0_6966 = (_zz_dataOut_payload_0_6964 ? _zz_dataOut_payload_0_6910 : _zz_dataOut_payload_0_6898);
  assign _zz_dataOut_payload_0_6967 = (_zz_dataOut_payload_0_6901 < _zz_dataOut_payload_0_6913);
  assign _zz_dataOut_payload_0_6968 = (_zz_dataOut_payload_0_6967 ? _zz_dataOut_payload_0_6901 : _zz_dataOut_payload_0_6913);
  assign _zz_dataOut_payload_0_6969 = (_zz_dataOut_payload_0_6967 ? _zz_dataOut_payload_0_6913 : _zz_dataOut_payload_0_6901);
  assign _zz_dataOut_payload_0_6970 = (_zz_dataOut_payload_0_6904 < _zz_dataOut_payload_0_6916);
  assign _zz_dataOut_payload_0_6971 = (_zz_dataOut_payload_0_6970 ? _zz_dataOut_payload_0_6904 : _zz_dataOut_payload_0_6916);
  assign _zz_dataOut_payload_0_6972 = (_zz_dataOut_payload_0_6970 ? _zz_dataOut_payload_0_6916 : _zz_dataOut_payload_0_6904);
  assign _zz_dataOut_payload_0_6973 = (_zz_dataOut_payload_0_6907 < _zz_dataOut_payload_0_6919);
  assign _zz_dataOut_payload_0_6974 = (_zz_dataOut_payload_0_6973 ? _zz_dataOut_payload_0_6907 : _zz_dataOut_payload_0_6919);
  assign _zz_dataOut_payload_0_6975 = (_zz_dataOut_payload_0_6973 ? _zz_dataOut_payload_0_6919 : _zz_dataOut_payload_0_6907);
  assign _zz_dataOut_payload_0_6976 = (_zz_dataOut_payload_0_6965 < _zz_dataOut_payload_0_6971);
  assign _zz_dataOut_payload_0_6977 = (_zz_dataOut_payload_0_6976 ? _zz_dataOut_payload_0_6965 : _zz_dataOut_payload_0_6971);
  assign _zz_dataOut_payload_0_6978 = (_zz_dataOut_payload_0_6976 ? _zz_dataOut_payload_0_6971 : _zz_dataOut_payload_0_6965);
  assign _zz_dataOut_payload_0_6979 = (_zz_dataOut_payload_0_6968 < _zz_dataOut_payload_0_6974);
  assign _zz_dataOut_payload_0_6980 = (_zz_dataOut_payload_0_6979 ? _zz_dataOut_payload_0_6968 : _zz_dataOut_payload_0_6974);
  assign _zz_dataOut_payload_0_6981 = (_zz_dataOut_payload_0_6979 ? _zz_dataOut_payload_0_6974 : _zz_dataOut_payload_0_6968);
  assign _zz_dataOut_payload_0_6982 = (_zz_dataOut_payload_0_6977 < _zz_dataOut_payload_0_6980);
  assign _zz_dataOut_payload_0_6983 = (_zz_dataOut_payload_0_6978 < _zz_dataOut_payload_0_6981);
  assign _zz_dataOut_payload_0_6988 = (_zz_dataOut_payload_0_6966 < _zz_dataOut_payload_0_6972);
  assign _zz_dataOut_payload_0_6989 = (_zz_dataOut_payload_0_6988 ? _zz_dataOut_payload_0_6966 : _zz_dataOut_payload_0_6972);
  assign _zz_dataOut_payload_0_6990 = (_zz_dataOut_payload_0_6988 ? _zz_dataOut_payload_0_6972 : _zz_dataOut_payload_0_6966);
  assign _zz_dataOut_payload_0_6991 = (_zz_dataOut_payload_0_6969 < _zz_dataOut_payload_0_6975);
  assign _zz_dataOut_payload_0_6992 = (_zz_dataOut_payload_0_6991 ? _zz_dataOut_payload_0_6969 : _zz_dataOut_payload_0_6975);
  assign _zz_dataOut_payload_0_6993 = (_zz_dataOut_payload_0_6991 ? _zz_dataOut_payload_0_6975 : _zz_dataOut_payload_0_6969);
  assign _zz_dataOut_payload_0_6994 = (_zz_dataOut_payload_0_6989 < _zz_dataOut_payload_0_6992);
  assign _zz_dataOut_payload_0_6995 = (_zz_dataOut_payload_0_6990 < _zz_dataOut_payload_0_6993);
  assign _zz_dataOut_payload_0_7056 = (_zz_dataOut_payload_0_5280 < _zz_dataOut_payload_0_5311);
  assign _zz_dataOut_payload_0_7057 = (_zz_dataOut_payload_0_7056 ? _zz_dataOut_payload_0_5280 : _zz_dataOut_payload_0_5311);
  assign _zz_dataOut_payload_0_7058 = (_zz_dataOut_payload_0_7056 ? _zz_dataOut_payload_0_5311 : _zz_dataOut_payload_0_5280);
  assign _zz_dataOut_payload_0_7059 = (_zz_dataOut_payload_0_5281 < _zz_dataOut_payload_0_5310);
  assign _zz_dataOut_payload_0_7060 = (_zz_dataOut_payload_0_7059 ? _zz_dataOut_payload_0_5281 : _zz_dataOut_payload_0_5310);
  assign _zz_dataOut_payload_0_7061 = (_zz_dataOut_payload_0_7059 ? _zz_dataOut_payload_0_5310 : _zz_dataOut_payload_0_5281);
  assign _zz_dataOut_payload_0_7062 = (_zz_dataOut_payload_0_5282 < _zz_dataOut_payload_0_5309);
  assign _zz_dataOut_payload_0_7063 = (_zz_dataOut_payload_0_7062 ? _zz_dataOut_payload_0_5282 : _zz_dataOut_payload_0_5309);
  assign _zz_dataOut_payload_0_7064 = (_zz_dataOut_payload_0_7062 ? _zz_dataOut_payload_0_5309 : _zz_dataOut_payload_0_5282);
  assign _zz_dataOut_payload_0_7065 = (_zz_dataOut_payload_0_5283 < _zz_dataOut_payload_0_5308);
  assign _zz_dataOut_payload_0_7066 = (_zz_dataOut_payload_0_7065 ? _zz_dataOut_payload_0_5283 : _zz_dataOut_payload_0_5308);
  assign _zz_dataOut_payload_0_7067 = (_zz_dataOut_payload_0_7065 ? _zz_dataOut_payload_0_5308 : _zz_dataOut_payload_0_5283);
  assign _zz_dataOut_payload_0_7068 = (_zz_dataOut_payload_0_5284 < _zz_dataOut_payload_0_5307);
  assign _zz_dataOut_payload_0_7069 = (_zz_dataOut_payload_0_7068 ? _zz_dataOut_payload_0_5284 : _zz_dataOut_payload_0_5307);
  assign _zz_dataOut_payload_0_7070 = (_zz_dataOut_payload_0_7068 ? _zz_dataOut_payload_0_5307 : _zz_dataOut_payload_0_5284);
  assign _zz_dataOut_payload_0_7071 = (_zz_dataOut_payload_0_5285 < _zz_dataOut_payload_0_5306);
  assign _zz_dataOut_payload_0_7072 = (_zz_dataOut_payload_0_7071 ? _zz_dataOut_payload_0_5285 : _zz_dataOut_payload_0_5306);
  assign _zz_dataOut_payload_0_7073 = (_zz_dataOut_payload_0_7071 ? _zz_dataOut_payload_0_5306 : _zz_dataOut_payload_0_5285);
  assign _zz_dataOut_payload_0_7074 = (_zz_dataOut_payload_0_5286 < _zz_dataOut_payload_0_5305);
  assign _zz_dataOut_payload_0_7075 = (_zz_dataOut_payload_0_7074 ? _zz_dataOut_payload_0_5286 : _zz_dataOut_payload_0_5305);
  assign _zz_dataOut_payload_0_7076 = (_zz_dataOut_payload_0_7074 ? _zz_dataOut_payload_0_5305 : _zz_dataOut_payload_0_5286);
  assign _zz_dataOut_payload_0_7077 = (_zz_dataOut_payload_0_5287 < _zz_dataOut_payload_0_5304);
  assign _zz_dataOut_payload_0_7078 = (_zz_dataOut_payload_0_7077 ? _zz_dataOut_payload_0_5287 : _zz_dataOut_payload_0_5304);
  assign _zz_dataOut_payload_0_7079 = (_zz_dataOut_payload_0_7077 ? _zz_dataOut_payload_0_5304 : _zz_dataOut_payload_0_5287);
  assign _zz_dataOut_payload_0_7080 = (_zz_dataOut_payload_0_5288 < _zz_dataOut_payload_0_5303);
  assign _zz_dataOut_payload_0_7081 = (_zz_dataOut_payload_0_7080 ? _zz_dataOut_payload_0_5288 : _zz_dataOut_payload_0_5303);
  assign _zz_dataOut_payload_0_7082 = (_zz_dataOut_payload_0_7080 ? _zz_dataOut_payload_0_5303 : _zz_dataOut_payload_0_5288);
  assign _zz_dataOut_payload_0_7083 = (_zz_dataOut_payload_0_5289 < _zz_dataOut_payload_0_5302);
  assign _zz_dataOut_payload_0_7084 = (_zz_dataOut_payload_0_7083 ? _zz_dataOut_payload_0_5289 : _zz_dataOut_payload_0_5302);
  assign _zz_dataOut_payload_0_7085 = (_zz_dataOut_payload_0_7083 ? _zz_dataOut_payload_0_5302 : _zz_dataOut_payload_0_5289);
  assign _zz_dataOut_payload_0_7086 = (_zz_dataOut_payload_0_5290 < _zz_dataOut_payload_0_5301);
  assign _zz_dataOut_payload_0_7087 = (_zz_dataOut_payload_0_7086 ? _zz_dataOut_payload_0_5290 : _zz_dataOut_payload_0_5301);
  assign _zz_dataOut_payload_0_7088 = (_zz_dataOut_payload_0_7086 ? _zz_dataOut_payload_0_5301 : _zz_dataOut_payload_0_5290);
  assign _zz_dataOut_payload_0_7089 = (_zz_dataOut_payload_0_5291 < _zz_dataOut_payload_0_5300);
  assign _zz_dataOut_payload_0_7090 = (_zz_dataOut_payload_0_7089 ? _zz_dataOut_payload_0_5291 : _zz_dataOut_payload_0_5300);
  assign _zz_dataOut_payload_0_7091 = (_zz_dataOut_payload_0_7089 ? _zz_dataOut_payload_0_5300 : _zz_dataOut_payload_0_5291);
  assign _zz_dataOut_payload_0_7092 = (_zz_dataOut_payload_0_5292 < _zz_dataOut_payload_0_5299);
  assign _zz_dataOut_payload_0_7093 = (_zz_dataOut_payload_0_7092 ? _zz_dataOut_payload_0_5292 : _zz_dataOut_payload_0_5299);
  assign _zz_dataOut_payload_0_7094 = (_zz_dataOut_payload_0_7092 ? _zz_dataOut_payload_0_5299 : _zz_dataOut_payload_0_5292);
  assign _zz_dataOut_payload_0_7095 = (_zz_dataOut_payload_0_5293 < _zz_dataOut_payload_0_5298);
  assign _zz_dataOut_payload_0_7096 = (_zz_dataOut_payload_0_7095 ? _zz_dataOut_payload_0_5293 : _zz_dataOut_payload_0_5298);
  assign _zz_dataOut_payload_0_7097 = (_zz_dataOut_payload_0_7095 ? _zz_dataOut_payload_0_5298 : _zz_dataOut_payload_0_5293);
  assign _zz_dataOut_payload_0_7098 = (_zz_dataOut_payload_0_5294 < _zz_dataOut_payload_0_5297);
  assign _zz_dataOut_payload_0_7099 = (_zz_dataOut_payload_0_7098 ? _zz_dataOut_payload_0_5294 : _zz_dataOut_payload_0_5297);
  assign _zz_dataOut_payload_0_7100 = (_zz_dataOut_payload_0_7098 ? _zz_dataOut_payload_0_5297 : _zz_dataOut_payload_0_5294);
  assign _zz_dataOut_payload_0_7101 = (_zz_dataOut_payload_0_5295 < _zz_dataOut_payload_0_5296);
  assign _zz_dataOut_payload_0_7102 = (_zz_dataOut_payload_0_7101 ? _zz_dataOut_payload_0_5295 : _zz_dataOut_payload_0_5296);
  assign _zz_dataOut_payload_0_7103 = (_zz_dataOut_payload_0_7101 ? _zz_dataOut_payload_0_5296 : _zz_dataOut_payload_0_5295);
  assign _zz_dataOut_payload_0_7104 = (_zz_dataOut_payload_0_7057 < _zz_dataOut_payload_0_7081);
  assign _zz_dataOut_payload_0_7105 = (_zz_dataOut_payload_0_7104 ? _zz_dataOut_payload_0_7057 : _zz_dataOut_payload_0_7081);
  assign _zz_dataOut_payload_0_7106 = (_zz_dataOut_payload_0_7104 ? _zz_dataOut_payload_0_7081 : _zz_dataOut_payload_0_7057);
  assign _zz_dataOut_payload_0_7107 = (_zz_dataOut_payload_0_7060 < _zz_dataOut_payload_0_7084);
  assign _zz_dataOut_payload_0_7108 = (_zz_dataOut_payload_0_7107 ? _zz_dataOut_payload_0_7060 : _zz_dataOut_payload_0_7084);
  assign _zz_dataOut_payload_0_7109 = (_zz_dataOut_payload_0_7107 ? _zz_dataOut_payload_0_7084 : _zz_dataOut_payload_0_7060);
  assign _zz_dataOut_payload_0_7110 = (_zz_dataOut_payload_0_7063 < _zz_dataOut_payload_0_7087);
  assign _zz_dataOut_payload_0_7111 = (_zz_dataOut_payload_0_7110 ? _zz_dataOut_payload_0_7063 : _zz_dataOut_payload_0_7087);
  assign _zz_dataOut_payload_0_7112 = (_zz_dataOut_payload_0_7110 ? _zz_dataOut_payload_0_7087 : _zz_dataOut_payload_0_7063);
  assign _zz_dataOut_payload_0_7113 = (_zz_dataOut_payload_0_7066 < _zz_dataOut_payload_0_7090);
  assign _zz_dataOut_payload_0_7114 = (_zz_dataOut_payload_0_7113 ? _zz_dataOut_payload_0_7066 : _zz_dataOut_payload_0_7090);
  assign _zz_dataOut_payload_0_7115 = (_zz_dataOut_payload_0_7113 ? _zz_dataOut_payload_0_7090 : _zz_dataOut_payload_0_7066);
  assign _zz_dataOut_payload_0_7116 = (_zz_dataOut_payload_0_7069 < _zz_dataOut_payload_0_7093);
  assign _zz_dataOut_payload_0_7117 = (_zz_dataOut_payload_0_7116 ? _zz_dataOut_payload_0_7069 : _zz_dataOut_payload_0_7093);
  assign _zz_dataOut_payload_0_7118 = (_zz_dataOut_payload_0_7116 ? _zz_dataOut_payload_0_7093 : _zz_dataOut_payload_0_7069);
  assign _zz_dataOut_payload_0_7119 = (_zz_dataOut_payload_0_7072 < _zz_dataOut_payload_0_7096);
  assign _zz_dataOut_payload_0_7120 = (_zz_dataOut_payload_0_7119 ? _zz_dataOut_payload_0_7072 : _zz_dataOut_payload_0_7096);
  assign _zz_dataOut_payload_0_7121 = (_zz_dataOut_payload_0_7119 ? _zz_dataOut_payload_0_7096 : _zz_dataOut_payload_0_7072);
  assign _zz_dataOut_payload_0_7122 = (_zz_dataOut_payload_0_7075 < _zz_dataOut_payload_0_7099);
  assign _zz_dataOut_payload_0_7123 = (_zz_dataOut_payload_0_7122 ? _zz_dataOut_payload_0_7075 : _zz_dataOut_payload_0_7099);
  assign _zz_dataOut_payload_0_7124 = (_zz_dataOut_payload_0_7122 ? _zz_dataOut_payload_0_7099 : _zz_dataOut_payload_0_7075);
  assign _zz_dataOut_payload_0_7125 = (_zz_dataOut_payload_0_7078 < _zz_dataOut_payload_0_7102);
  assign _zz_dataOut_payload_0_7126 = (_zz_dataOut_payload_0_7125 ? _zz_dataOut_payload_0_7078 : _zz_dataOut_payload_0_7102);
  assign _zz_dataOut_payload_0_7127 = (_zz_dataOut_payload_0_7125 ? _zz_dataOut_payload_0_7102 : _zz_dataOut_payload_0_7078);
  assign _zz_dataOut_payload_0_7128 = (_zz_dataOut_payload_0_7105 < _zz_dataOut_payload_0_7117);
  assign _zz_dataOut_payload_0_7129 = (_zz_dataOut_payload_0_7128 ? _zz_dataOut_payload_0_7105 : _zz_dataOut_payload_0_7117);
  assign _zz_dataOut_payload_0_7130 = (_zz_dataOut_payload_0_7128 ? _zz_dataOut_payload_0_7117 : _zz_dataOut_payload_0_7105);
  assign _zz_dataOut_payload_0_7131 = (_zz_dataOut_payload_0_7108 < _zz_dataOut_payload_0_7120);
  assign _zz_dataOut_payload_0_7132 = (_zz_dataOut_payload_0_7131 ? _zz_dataOut_payload_0_7108 : _zz_dataOut_payload_0_7120);
  assign _zz_dataOut_payload_0_7133 = (_zz_dataOut_payload_0_7131 ? _zz_dataOut_payload_0_7120 : _zz_dataOut_payload_0_7108);
  assign _zz_dataOut_payload_0_7134 = (_zz_dataOut_payload_0_7111 < _zz_dataOut_payload_0_7123);
  assign _zz_dataOut_payload_0_7135 = (_zz_dataOut_payload_0_7134 ? _zz_dataOut_payload_0_7111 : _zz_dataOut_payload_0_7123);
  assign _zz_dataOut_payload_0_7136 = (_zz_dataOut_payload_0_7134 ? _zz_dataOut_payload_0_7123 : _zz_dataOut_payload_0_7111);
  assign _zz_dataOut_payload_0_7137 = (_zz_dataOut_payload_0_7114 < _zz_dataOut_payload_0_7126);
  assign _zz_dataOut_payload_0_7138 = (_zz_dataOut_payload_0_7137 ? _zz_dataOut_payload_0_7114 : _zz_dataOut_payload_0_7126);
  assign _zz_dataOut_payload_0_7139 = (_zz_dataOut_payload_0_7137 ? _zz_dataOut_payload_0_7126 : _zz_dataOut_payload_0_7114);
  assign _zz_dataOut_payload_0_7140 = (_zz_dataOut_payload_0_7129 < _zz_dataOut_payload_0_7135);
  assign _zz_dataOut_payload_0_7141 = (_zz_dataOut_payload_0_7140 ? _zz_dataOut_payload_0_7129 : _zz_dataOut_payload_0_7135);
  assign _zz_dataOut_payload_0_7142 = (_zz_dataOut_payload_0_7140 ? _zz_dataOut_payload_0_7135 : _zz_dataOut_payload_0_7129);
  assign _zz_dataOut_payload_0_7143 = (_zz_dataOut_payload_0_7132 < _zz_dataOut_payload_0_7138);
  assign _zz_dataOut_payload_0_7144 = (_zz_dataOut_payload_0_7143 ? _zz_dataOut_payload_0_7132 : _zz_dataOut_payload_0_7138);
  assign _zz_dataOut_payload_0_7145 = (_zz_dataOut_payload_0_7143 ? _zz_dataOut_payload_0_7138 : _zz_dataOut_payload_0_7132);
  assign _zz_dataOut_payload_0_7146 = (_zz_dataOut_payload_0_7141 < _zz_dataOut_payload_0_7144);
  assign _zz_dataOut_payload_0_7147 = (_zz_dataOut_payload_0_7142 < _zz_dataOut_payload_0_7145);
  assign _zz_dataOut_payload_0_7152 = (_zz_dataOut_payload_0_7130 < _zz_dataOut_payload_0_7136);
  assign _zz_dataOut_payload_0_7153 = (_zz_dataOut_payload_0_7152 ? _zz_dataOut_payload_0_7130 : _zz_dataOut_payload_0_7136);
  assign _zz_dataOut_payload_0_7154 = (_zz_dataOut_payload_0_7152 ? _zz_dataOut_payload_0_7136 : _zz_dataOut_payload_0_7130);
  assign _zz_dataOut_payload_0_7155 = (_zz_dataOut_payload_0_7133 < _zz_dataOut_payload_0_7139);
  assign _zz_dataOut_payload_0_7156 = (_zz_dataOut_payload_0_7155 ? _zz_dataOut_payload_0_7133 : _zz_dataOut_payload_0_7139);
  assign _zz_dataOut_payload_0_7157 = (_zz_dataOut_payload_0_7155 ? _zz_dataOut_payload_0_7139 : _zz_dataOut_payload_0_7133);
  assign _zz_dataOut_payload_0_7158 = (_zz_dataOut_payload_0_7153 < _zz_dataOut_payload_0_7156);
  assign _zz_dataOut_payload_0_7159 = (_zz_dataOut_payload_0_7154 < _zz_dataOut_payload_0_7157);
  assign _zz_dataOut_payload_0_7172 = (_zz_dataOut_payload_0_7106 < _zz_dataOut_payload_0_7118);
  assign _zz_dataOut_payload_0_7173 = (_zz_dataOut_payload_0_7172 ? _zz_dataOut_payload_0_7106 : _zz_dataOut_payload_0_7118);
  assign _zz_dataOut_payload_0_7174 = (_zz_dataOut_payload_0_7172 ? _zz_dataOut_payload_0_7118 : _zz_dataOut_payload_0_7106);
  assign _zz_dataOut_payload_0_7175 = (_zz_dataOut_payload_0_7109 < _zz_dataOut_payload_0_7121);
  assign _zz_dataOut_payload_0_7176 = (_zz_dataOut_payload_0_7175 ? _zz_dataOut_payload_0_7109 : _zz_dataOut_payload_0_7121);
  assign _zz_dataOut_payload_0_7177 = (_zz_dataOut_payload_0_7175 ? _zz_dataOut_payload_0_7121 : _zz_dataOut_payload_0_7109);
  assign _zz_dataOut_payload_0_7178 = (_zz_dataOut_payload_0_7112 < _zz_dataOut_payload_0_7124);
  assign _zz_dataOut_payload_0_7179 = (_zz_dataOut_payload_0_7178 ? _zz_dataOut_payload_0_7112 : _zz_dataOut_payload_0_7124);
  assign _zz_dataOut_payload_0_7180 = (_zz_dataOut_payload_0_7178 ? _zz_dataOut_payload_0_7124 : _zz_dataOut_payload_0_7112);
  assign _zz_dataOut_payload_0_7181 = (_zz_dataOut_payload_0_7115 < _zz_dataOut_payload_0_7127);
  assign _zz_dataOut_payload_0_7182 = (_zz_dataOut_payload_0_7181 ? _zz_dataOut_payload_0_7115 : _zz_dataOut_payload_0_7127);
  assign _zz_dataOut_payload_0_7183 = (_zz_dataOut_payload_0_7181 ? _zz_dataOut_payload_0_7127 : _zz_dataOut_payload_0_7115);
  assign _zz_dataOut_payload_0_7184 = (_zz_dataOut_payload_0_7173 < _zz_dataOut_payload_0_7179);
  assign _zz_dataOut_payload_0_7185 = (_zz_dataOut_payload_0_7184 ? _zz_dataOut_payload_0_7173 : _zz_dataOut_payload_0_7179);
  assign _zz_dataOut_payload_0_7186 = (_zz_dataOut_payload_0_7184 ? _zz_dataOut_payload_0_7179 : _zz_dataOut_payload_0_7173);
  assign _zz_dataOut_payload_0_7187 = (_zz_dataOut_payload_0_7176 < _zz_dataOut_payload_0_7182);
  assign _zz_dataOut_payload_0_7188 = (_zz_dataOut_payload_0_7187 ? _zz_dataOut_payload_0_7176 : _zz_dataOut_payload_0_7182);
  assign _zz_dataOut_payload_0_7189 = (_zz_dataOut_payload_0_7187 ? _zz_dataOut_payload_0_7182 : _zz_dataOut_payload_0_7176);
  assign _zz_dataOut_payload_0_7190 = (_zz_dataOut_payload_0_7185 < _zz_dataOut_payload_0_7188);
  assign _zz_dataOut_payload_0_7191 = (_zz_dataOut_payload_0_7186 < _zz_dataOut_payload_0_7189);
  assign _zz_dataOut_payload_0_7196 = (_zz_dataOut_payload_0_7174 < _zz_dataOut_payload_0_7180);
  assign _zz_dataOut_payload_0_7197 = (_zz_dataOut_payload_0_7196 ? _zz_dataOut_payload_0_7174 : _zz_dataOut_payload_0_7180);
  assign _zz_dataOut_payload_0_7198 = (_zz_dataOut_payload_0_7196 ? _zz_dataOut_payload_0_7180 : _zz_dataOut_payload_0_7174);
  assign _zz_dataOut_payload_0_7199 = (_zz_dataOut_payload_0_7177 < _zz_dataOut_payload_0_7183);
  assign _zz_dataOut_payload_0_7200 = (_zz_dataOut_payload_0_7199 ? _zz_dataOut_payload_0_7177 : _zz_dataOut_payload_0_7183);
  assign _zz_dataOut_payload_0_7201 = (_zz_dataOut_payload_0_7199 ? _zz_dataOut_payload_0_7183 : _zz_dataOut_payload_0_7177);
  assign _zz_dataOut_payload_0_7202 = (_zz_dataOut_payload_0_7197 < _zz_dataOut_payload_0_7200);
  assign _zz_dataOut_payload_0_7203 = (_zz_dataOut_payload_0_7198 < _zz_dataOut_payload_0_7201);
  assign _zz_dataOut_payload_0_7232 = (_zz_dataOut_payload_0_7103 < _zz_dataOut_payload_0_7079);
  assign _zz_dataOut_payload_0_7233 = (_zz_dataOut_payload_0_7232 ? _zz_dataOut_payload_0_7103 : _zz_dataOut_payload_0_7079);
  assign _zz_dataOut_payload_0_7234 = (_zz_dataOut_payload_0_7232 ? _zz_dataOut_payload_0_7079 : _zz_dataOut_payload_0_7103);
  assign _zz_dataOut_payload_0_7235 = (_zz_dataOut_payload_0_7100 < _zz_dataOut_payload_0_7076);
  assign _zz_dataOut_payload_0_7236 = (_zz_dataOut_payload_0_7235 ? _zz_dataOut_payload_0_7100 : _zz_dataOut_payload_0_7076);
  assign _zz_dataOut_payload_0_7237 = (_zz_dataOut_payload_0_7235 ? _zz_dataOut_payload_0_7076 : _zz_dataOut_payload_0_7100);
  assign _zz_dataOut_payload_0_7238 = (_zz_dataOut_payload_0_7097 < _zz_dataOut_payload_0_7073);
  assign _zz_dataOut_payload_0_7239 = (_zz_dataOut_payload_0_7238 ? _zz_dataOut_payload_0_7097 : _zz_dataOut_payload_0_7073);
  assign _zz_dataOut_payload_0_7240 = (_zz_dataOut_payload_0_7238 ? _zz_dataOut_payload_0_7073 : _zz_dataOut_payload_0_7097);
  assign _zz_dataOut_payload_0_7241 = (_zz_dataOut_payload_0_7094 < _zz_dataOut_payload_0_7070);
  assign _zz_dataOut_payload_0_7242 = (_zz_dataOut_payload_0_7241 ? _zz_dataOut_payload_0_7094 : _zz_dataOut_payload_0_7070);
  assign _zz_dataOut_payload_0_7243 = (_zz_dataOut_payload_0_7241 ? _zz_dataOut_payload_0_7070 : _zz_dataOut_payload_0_7094);
  assign _zz_dataOut_payload_0_7244 = (_zz_dataOut_payload_0_7091 < _zz_dataOut_payload_0_7067);
  assign _zz_dataOut_payload_0_7245 = (_zz_dataOut_payload_0_7244 ? _zz_dataOut_payload_0_7091 : _zz_dataOut_payload_0_7067);
  assign _zz_dataOut_payload_0_7246 = (_zz_dataOut_payload_0_7244 ? _zz_dataOut_payload_0_7067 : _zz_dataOut_payload_0_7091);
  assign _zz_dataOut_payload_0_7247 = (_zz_dataOut_payload_0_7088 < _zz_dataOut_payload_0_7064);
  assign _zz_dataOut_payload_0_7248 = (_zz_dataOut_payload_0_7247 ? _zz_dataOut_payload_0_7088 : _zz_dataOut_payload_0_7064);
  assign _zz_dataOut_payload_0_7249 = (_zz_dataOut_payload_0_7247 ? _zz_dataOut_payload_0_7064 : _zz_dataOut_payload_0_7088);
  assign _zz_dataOut_payload_0_7250 = (_zz_dataOut_payload_0_7085 < _zz_dataOut_payload_0_7061);
  assign _zz_dataOut_payload_0_7251 = (_zz_dataOut_payload_0_7250 ? _zz_dataOut_payload_0_7085 : _zz_dataOut_payload_0_7061);
  assign _zz_dataOut_payload_0_7252 = (_zz_dataOut_payload_0_7250 ? _zz_dataOut_payload_0_7061 : _zz_dataOut_payload_0_7085);
  assign _zz_dataOut_payload_0_7253 = (_zz_dataOut_payload_0_7082 < _zz_dataOut_payload_0_7058);
  assign _zz_dataOut_payload_0_7254 = (_zz_dataOut_payload_0_7253 ? _zz_dataOut_payload_0_7082 : _zz_dataOut_payload_0_7058);
  assign _zz_dataOut_payload_0_7255 = (_zz_dataOut_payload_0_7253 ? _zz_dataOut_payload_0_7058 : _zz_dataOut_payload_0_7082);
  assign _zz_dataOut_payload_0_7256 = (_zz_dataOut_payload_0_7233 < _zz_dataOut_payload_0_7245);
  assign _zz_dataOut_payload_0_7257 = (_zz_dataOut_payload_0_7256 ? _zz_dataOut_payload_0_7233 : _zz_dataOut_payload_0_7245);
  assign _zz_dataOut_payload_0_7258 = (_zz_dataOut_payload_0_7256 ? _zz_dataOut_payload_0_7245 : _zz_dataOut_payload_0_7233);
  assign _zz_dataOut_payload_0_7259 = (_zz_dataOut_payload_0_7236 < _zz_dataOut_payload_0_7248);
  assign _zz_dataOut_payload_0_7260 = (_zz_dataOut_payload_0_7259 ? _zz_dataOut_payload_0_7236 : _zz_dataOut_payload_0_7248);
  assign _zz_dataOut_payload_0_7261 = (_zz_dataOut_payload_0_7259 ? _zz_dataOut_payload_0_7248 : _zz_dataOut_payload_0_7236);
  assign _zz_dataOut_payload_0_7262 = (_zz_dataOut_payload_0_7239 < _zz_dataOut_payload_0_7251);
  assign _zz_dataOut_payload_0_7263 = (_zz_dataOut_payload_0_7262 ? _zz_dataOut_payload_0_7239 : _zz_dataOut_payload_0_7251);
  assign _zz_dataOut_payload_0_7264 = (_zz_dataOut_payload_0_7262 ? _zz_dataOut_payload_0_7251 : _zz_dataOut_payload_0_7239);
  assign _zz_dataOut_payload_0_7265 = (_zz_dataOut_payload_0_7242 < _zz_dataOut_payload_0_7254);
  assign _zz_dataOut_payload_0_7266 = (_zz_dataOut_payload_0_7265 ? _zz_dataOut_payload_0_7242 : _zz_dataOut_payload_0_7254);
  assign _zz_dataOut_payload_0_7267 = (_zz_dataOut_payload_0_7265 ? _zz_dataOut_payload_0_7254 : _zz_dataOut_payload_0_7242);
  assign _zz_dataOut_payload_0_7268 = (_zz_dataOut_payload_0_7257 < _zz_dataOut_payload_0_7263);
  assign _zz_dataOut_payload_0_7269 = (_zz_dataOut_payload_0_7268 ? _zz_dataOut_payload_0_7257 : _zz_dataOut_payload_0_7263);
  assign _zz_dataOut_payload_0_7270 = (_zz_dataOut_payload_0_7268 ? _zz_dataOut_payload_0_7263 : _zz_dataOut_payload_0_7257);
  assign _zz_dataOut_payload_0_7271 = (_zz_dataOut_payload_0_7260 < _zz_dataOut_payload_0_7266);
  assign _zz_dataOut_payload_0_7272 = (_zz_dataOut_payload_0_7271 ? _zz_dataOut_payload_0_7260 : _zz_dataOut_payload_0_7266);
  assign _zz_dataOut_payload_0_7273 = (_zz_dataOut_payload_0_7271 ? _zz_dataOut_payload_0_7266 : _zz_dataOut_payload_0_7260);
  assign _zz_dataOut_payload_0_7274 = (_zz_dataOut_payload_0_7269 < _zz_dataOut_payload_0_7272);
  assign _zz_dataOut_payload_0_7275 = (_zz_dataOut_payload_0_7270 < _zz_dataOut_payload_0_7273);
  assign _zz_dataOut_payload_0_7280 = (_zz_dataOut_payload_0_7258 < _zz_dataOut_payload_0_7264);
  assign _zz_dataOut_payload_0_7281 = (_zz_dataOut_payload_0_7280 ? _zz_dataOut_payload_0_7258 : _zz_dataOut_payload_0_7264);
  assign _zz_dataOut_payload_0_7282 = (_zz_dataOut_payload_0_7280 ? _zz_dataOut_payload_0_7264 : _zz_dataOut_payload_0_7258);
  assign _zz_dataOut_payload_0_7283 = (_zz_dataOut_payload_0_7261 < _zz_dataOut_payload_0_7267);
  assign _zz_dataOut_payload_0_7284 = (_zz_dataOut_payload_0_7283 ? _zz_dataOut_payload_0_7261 : _zz_dataOut_payload_0_7267);
  assign _zz_dataOut_payload_0_7285 = (_zz_dataOut_payload_0_7283 ? _zz_dataOut_payload_0_7267 : _zz_dataOut_payload_0_7261);
  assign _zz_dataOut_payload_0_7286 = (_zz_dataOut_payload_0_7281 < _zz_dataOut_payload_0_7284);
  assign _zz_dataOut_payload_0_7287 = (_zz_dataOut_payload_0_7282 < _zz_dataOut_payload_0_7285);
  assign _zz_dataOut_payload_0_7300 = (_zz_dataOut_payload_0_7234 < _zz_dataOut_payload_0_7246);
  assign _zz_dataOut_payload_0_7301 = (_zz_dataOut_payload_0_7300 ? _zz_dataOut_payload_0_7234 : _zz_dataOut_payload_0_7246);
  assign _zz_dataOut_payload_0_7302 = (_zz_dataOut_payload_0_7300 ? _zz_dataOut_payload_0_7246 : _zz_dataOut_payload_0_7234);
  assign _zz_dataOut_payload_0_7303 = (_zz_dataOut_payload_0_7237 < _zz_dataOut_payload_0_7249);
  assign _zz_dataOut_payload_0_7304 = (_zz_dataOut_payload_0_7303 ? _zz_dataOut_payload_0_7237 : _zz_dataOut_payload_0_7249);
  assign _zz_dataOut_payload_0_7305 = (_zz_dataOut_payload_0_7303 ? _zz_dataOut_payload_0_7249 : _zz_dataOut_payload_0_7237);
  assign _zz_dataOut_payload_0_7306 = (_zz_dataOut_payload_0_7240 < _zz_dataOut_payload_0_7252);
  assign _zz_dataOut_payload_0_7307 = (_zz_dataOut_payload_0_7306 ? _zz_dataOut_payload_0_7240 : _zz_dataOut_payload_0_7252);
  assign _zz_dataOut_payload_0_7308 = (_zz_dataOut_payload_0_7306 ? _zz_dataOut_payload_0_7252 : _zz_dataOut_payload_0_7240);
  assign _zz_dataOut_payload_0_7309 = (_zz_dataOut_payload_0_7243 < _zz_dataOut_payload_0_7255);
  assign _zz_dataOut_payload_0_7310 = (_zz_dataOut_payload_0_7309 ? _zz_dataOut_payload_0_7243 : _zz_dataOut_payload_0_7255);
  assign _zz_dataOut_payload_0_7311 = (_zz_dataOut_payload_0_7309 ? _zz_dataOut_payload_0_7255 : _zz_dataOut_payload_0_7243);
  assign _zz_dataOut_payload_0_7312 = (_zz_dataOut_payload_0_7301 < _zz_dataOut_payload_0_7307);
  assign _zz_dataOut_payload_0_7313 = (_zz_dataOut_payload_0_7312 ? _zz_dataOut_payload_0_7301 : _zz_dataOut_payload_0_7307);
  assign _zz_dataOut_payload_0_7314 = (_zz_dataOut_payload_0_7312 ? _zz_dataOut_payload_0_7307 : _zz_dataOut_payload_0_7301);
  assign _zz_dataOut_payload_0_7315 = (_zz_dataOut_payload_0_7304 < _zz_dataOut_payload_0_7310);
  assign _zz_dataOut_payload_0_7316 = (_zz_dataOut_payload_0_7315 ? _zz_dataOut_payload_0_7304 : _zz_dataOut_payload_0_7310);
  assign _zz_dataOut_payload_0_7317 = (_zz_dataOut_payload_0_7315 ? _zz_dataOut_payload_0_7310 : _zz_dataOut_payload_0_7304);
  assign _zz_dataOut_payload_0_7318 = (_zz_dataOut_payload_0_7313 < _zz_dataOut_payload_0_7316);
  assign _zz_dataOut_payload_0_7319 = (_zz_dataOut_payload_0_7314 < _zz_dataOut_payload_0_7317);
  assign _zz_dataOut_payload_0_7324 = (_zz_dataOut_payload_0_7302 < _zz_dataOut_payload_0_7308);
  assign _zz_dataOut_payload_0_7325 = (_zz_dataOut_payload_0_7324 ? _zz_dataOut_payload_0_7302 : _zz_dataOut_payload_0_7308);
  assign _zz_dataOut_payload_0_7326 = (_zz_dataOut_payload_0_7324 ? _zz_dataOut_payload_0_7308 : _zz_dataOut_payload_0_7302);
  assign _zz_dataOut_payload_0_7327 = (_zz_dataOut_payload_0_7305 < _zz_dataOut_payload_0_7311);
  assign _zz_dataOut_payload_0_7328 = (_zz_dataOut_payload_0_7327 ? _zz_dataOut_payload_0_7305 : _zz_dataOut_payload_0_7311);
  assign _zz_dataOut_payload_0_7329 = (_zz_dataOut_payload_0_7327 ? _zz_dataOut_payload_0_7311 : _zz_dataOut_payload_0_7305);
  assign _zz_dataOut_payload_0_7330 = (_zz_dataOut_payload_0_7325 < _zz_dataOut_payload_0_7328);
  assign _zz_dataOut_payload_0_7331 = (_zz_dataOut_payload_0_7326 < _zz_dataOut_payload_0_7329);
  assign _zz_dataOut_payload_0_7392 = (_zz_dataOut_payload_0_5312 < _zz_dataOut_payload_0_5343);
  assign _zz_dataOut_payload_0_7393 = (_zz_dataOut_payload_0_7392 ? _zz_dataOut_payload_0_5312 : _zz_dataOut_payload_0_5343);
  assign _zz_dataOut_payload_0_7394 = (_zz_dataOut_payload_0_7392 ? _zz_dataOut_payload_0_5343 : _zz_dataOut_payload_0_5312);
  assign _zz_dataOut_payload_0_7395 = (_zz_dataOut_payload_0_5313 < _zz_dataOut_payload_0_5342);
  assign _zz_dataOut_payload_0_7396 = (_zz_dataOut_payload_0_7395 ? _zz_dataOut_payload_0_5313 : _zz_dataOut_payload_0_5342);
  assign _zz_dataOut_payload_0_7397 = (_zz_dataOut_payload_0_7395 ? _zz_dataOut_payload_0_5342 : _zz_dataOut_payload_0_5313);
  assign _zz_dataOut_payload_0_7398 = (_zz_dataOut_payload_0_5314 < _zz_dataOut_payload_0_5341);
  assign _zz_dataOut_payload_0_7399 = (_zz_dataOut_payload_0_7398 ? _zz_dataOut_payload_0_5314 : _zz_dataOut_payload_0_5341);
  assign _zz_dataOut_payload_0_7400 = (_zz_dataOut_payload_0_7398 ? _zz_dataOut_payload_0_5341 : _zz_dataOut_payload_0_5314);
  assign _zz_dataOut_payload_0_7401 = (_zz_dataOut_payload_0_5315 < _zz_dataOut_payload_0_5340);
  assign _zz_dataOut_payload_0_7402 = (_zz_dataOut_payload_0_7401 ? _zz_dataOut_payload_0_5315 : _zz_dataOut_payload_0_5340);
  assign _zz_dataOut_payload_0_7403 = (_zz_dataOut_payload_0_7401 ? _zz_dataOut_payload_0_5340 : _zz_dataOut_payload_0_5315);
  assign _zz_dataOut_payload_0_7404 = (_zz_dataOut_payload_0_5316 < _zz_dataOut_payload_0_5339);
  assign _zz_dataOut_payload_0_7405 = (_zz_dataOut_payload_0_7404 ? _zz_dataOut_payload_0_5316 : _zz_dataOut_payload_0_5339);
  assign _zz_dataOut_payload_0_7406 = (_zz_dataOut_payload_0_7404 ? _zz_dataOut_payload_0_5339 : _zz_dataOut_payload_0_5316);
  assign _zz_dataOut_payload_0_7407 = (_zz_dataOut_payload_0_5317 < _zz_dataOut_payload_0_5338);
  assign _zz_dataOut_payload_0_7408 = (_zz_dataOut_payload_0_7407 ? _zz_dataOut_payload_0_5317 : _zz_dataOut_payload_0_5338);
  assign _zz_dataOut_payload_0_7409 = (_zz_dataOut_payload_0_7407 ? _zz_dataOut_payload_0_5338 : _zz_dataOut_payload_0_5317);
  assign _zz_dataOut_payload_0_7410 = (_zz_dataOut_payload_0_5318 < _zz_dataOut_payload_0_5337);
  assign _zz_dataOut_payload_0_7411 = (_zz_dataOut_payload_0_7410 ? _zz_dataOut_payload_0_5318 : _zz_dataOut_payload_0_5337);
  assign _zz_dataOut_payload_0_7412 = (_zz_dataOut_payload_0_7410 ? _zz_dataOut_payload_0_5337 : _zz_dataOut_payload_0_5318);
  assign _zz_dataOut_payload_0_7413 = (_zz_dataOut_payload_0_5319 < _zz_dataOut_payload_0_5336);
  assign _zz_dataOut_payload_0_7414 = (_zz_dataOut_payload_0_7413 ? _zz_dataOut_payload_0_5319 : _zz_dataOut_payload_0_5336);
  assign _zz_dataOut_payload_0_7415 = (_zz_dataOut_payload_0_7413 ? _zz_dataOut_payload_0_5336 : _zz_dataOut_payload_0_5319);
  assign _zz_dataOut_payload_0_7416 = (_zz_dataOut_payload_0_5320 < _zz_dataOut_payload_0_5335);
  assign _zz_dataOut_payload_0_7417 = (_zz_dataOut_payload_0_7416 ? _zz_dataOut_payload_0_5320 : _zz_dataOut_payload_0_5335);
  assign _zz_dataOut_payload_0_7418 = (_zz_dataOut_payload_0_7416 ? _zz_dataOut_payload_0_5335 : _zz_dataOut_payload_0_5320);
  assign _zz_dataOut_payload_0_7419 = (_zz_dataOut_payload_0_5321 < _zz_dataOut_payload_0_5334);
  assign _zz_dataOut_payload_0_7420 = (_zz_dataOut_payload_0_7419 ? _zz_dataOut_payload_0_5321 : _zz_dataOut_payload_0_5334);
  assign _zz_dataOut_payload_0_7421 = (_zz_dataOut_payload_0_7419 ? _zz_dataOut_payload_0_5334 : _zz_dataOut_payload_0_5321);
  assign _zz_dataOut_payload_0_7422 = (_zz_dataOut_payload_0_5322 < _zz_dataOut_payload_0_5333);
  assign _zz_dataOut_payload_0_7423 = (_zz_dataOut_payload_0_7422 ? _zz_dataOut_payload_0_5322 : _zz_dataOut_payload_0_5333);
  assign _zz_dataOut_payload_0_7424 = (_zz_dataOut_payload_0_7422 ? _zz_dataOut_payload_0_5333 : _zz_dataOut_payload_0_5322);
  assign _zz_dataOut_payload_0_7425 = (_zz_dataOut_payload_0_5323 < _zz_dataOut_payload_0_5332);
  assign _zz_dataOut_payload_0_7426 = (_zz_dataOut_payload_0_7425 ? _zz_dataOut_payload_0_5323 : _zz_dataOut_payload_0_5332);
  assign _zz_dataOut_payload_0_7427 = (_zz_dataOut_payload_0_7425 ? _zz_dataOut_payload_0_5332 : _zz_dataOut_payload_0_5323);
  assign _zz_dataOut_payload_0_7428 = (_zz_dataOut_payload_0_5324 < _zz_dataOut_payload_0_5331);
  assign _zz_dataOut_payload_0_7429 = (_zz_dataOut_payload_0_7428 ? _zz_dataOut_payload_0_5324 : _zz_dataOut_payload_0_5331);
  assign _zz_dataOut_payload_0_7430 = (_zz_dataOut_payload_0_7428 ? _zz_dataOut_payload_0_5331 : _zz_dataOut_payload_0_5324);
  assign _zz_dataOut_payload_0_7431 = (_zz_dataOut_payload_0_5325 < _zz_dataOut_payload_0_5330);
  assign _zz_dataOut_payload_0_7432 = (_zz_dataOut_payload_0_7431 ? _zz_dataOut_payload_0_5325 : _zz_dataOut_payload_0_5330);
  assign _zz_dataOut_payload_0_7433 = (_zz_dataOut_payload_0_7431 ? _zz_dataOut_payload_0_5330 : _zz_dataOut_payload_0_5325);
  assign _zz_dataOut_payload_0_7434 = (_zz_dataOut_payload_0_5326 < _zz_dataOut_payload_0_5329);
  assign _zz_dataOut_payload_0_7435 = (_zz_dataOut_payload_0_7434 ? _zz_dataOut_payload_0_5326 : _zz_dataOut_payload_0_5329);
  assign _zz_dataOut_payload_0_7436 = (_zz_dataOut_payload_0_7434 ? _zz_dataOut_payload_0_5329 : _zz_dataOut_payload_0_5326);
  assign _zz_dataOut_payload_0_7437 = (_zz_dataOut_payload_0_5327 < _zz_dataOut_payload_0_5328);
  assign _zz_dataOut_payload_0_7438 = (_zz_dataOut_payload_0_7437 ? _zz_dataOut_payload_0_5327 : _zz_dataOut_payload_0_5328);
  assign _zz_dataOut_payload_0_7439 = (_zz_dataOut_payload_0_7437 ? _zz_dataOut_payload_0_5328 : _zz_dataOut_payload_0_5327);
  assign _zz_dataOut_payload_0_7440 = (_zz_dataOut_payload_0_7393 < _zz_dataOut_payload_0_7417);
  assign _zz_dataOut_payload_0_7441 = (_zz_dataOut_payload_0_7440 ? _zz_dataOut_payload_0_7393 : _zz_dataOut_payload_0_7417);
  assign _zz_dataOut_payload_0_7442 = (_zz_dataOut_payload_0_7440 ? _zz_dataOut_payload_0_7417 : _zz_dataOut_payload_0_7393);
  assign _zz_dataOut_payload_0_7443 = (_zz_dataOut_payload_0_7396 < _zz_dataOut_payload_0_7420);
  assign _zz_dataOut_payload_0_7444 = (_zz_dataOut_payload_0_7443 ? _zz_dataOut_payload_0_7396 : _zz_dataOut_payload_0_7420);
  assign _zz_dataOut_payload_0_7445 = (_zz_dataOut_payload_0_7443 ? _zz_dataOut_payload_0_7420 : _zz_dataOut_payload_0_7396);
  assign _zz_dataOut_payload_0_7446 = (_zz_dataOut_payload_0_7399 < _zz_dataOut_payload_0_7423);
  assign _zz_dataOut_payload_0_7447 = (_zz_dataOut_payload_0_7446 ? _zz_dataOut_payload_0_7399 : _zz_dataOut_payload_0_7423);
  assign _zz_dataOut_payload_0_7448 = (_zz_dataOut_payload_0_7446 ? _zz_dataOut_payload_0_7423 : _zz_dataOut_payload_0_7399);
  assign _zz_dataOut_payload_0_7449 = (_zz_dataOut_payload_0_7402 < _zz_dataOut_payload_0_7426);
  assign _zz_dataOut_payload_0_7450 = (_zz_dataOut_payload_0_7449 ? _zz_dataOut_payload_0_7402 : _zz_dataOut_payload_0_7426);
  assign _zz_dataOut_payload_0_7451 = (_zz_dataOut_payload_0_7449 ? _zz_dataOut_payload_0_7426 : _zz_dataOut_payload_0_7402);
  assign _zz_dataOut_payload_0_7452 = (_zz_dataOut_payload_0_7405 < _zz_dataOut_payload_0_7429);
  assign _zz_dataOut_payload_0_7453 = (_zz_dataOut_payload_0_7452 ? _zz_dataOut_payload_0_7405 : _zz_dataOut_payload_0_7429);
  assign _zz_dataOut_payload_0_7454 = (_zz_dataOut_payload_0_7452 ? _zz_dataOut_payload_0_7429 : _zz_dataOut_payload_0_7405);
  assign _zz_dataOut_payload_0_7455 = (_zz_dataOut_payload_0_7408 < _zz_dataOut_payload_0_7432);
  assign _zz_dataOut_payload_0_7456 = (_zz_dataOut_payload_0_7455 ? _zz_dataOut_payload_0_7408 : _zz_dataOut_payload_0_7432);
  assign _zz_dataOut_payload_0_7457 = (_zz_dataOut_payload_0_7455 ? _zz_dataOut_payload_0_7432 : _zz_dataOut_payload_0_7408);
  assign _zz_dataOut_payload_0_7458 = (_zz_dataOut_payload_0_7411 < _zz_dataOut_payload_0_7435);
  assign _zz_dataOut_payload_0_7459 = (_zz_dataOut_payload_0_7458 ? _zz_dataOut_payload_0_7411 : _zz_dataOut_payload_0_7435);
  assign _zz_dataOut_payload_0_7460 = (_zz_dataOut_payload_0_7458 ? _zz_dataOut_payload_0_7435 : _zz_dataOut_payload_0_7411);
  assign _zz_dataOut_payload_0_7461 = (_zz_dataOut_payload_0_7414 < _zz_dataOut_payload_0_7438);
  assign _zz_dataOut_payload_0_7462 = (_zz_dataOut_payload_0_7461 ? _zz_dataOut_payload_0_7414 : _zz_dataOut_payload_0_7438);
  assign _zz_dataOut_payload_0_7463 = (_zz_dataOut_payload_0_7461 ? _zz_dataOut_payload_0_7438 : _zz_dataOut_payload_0_7414);
  assign _zz_dataOut_payload_0_7464 = (_zz_dataOut_payload_0_7441 < _zz_dataOut_payload_0_7453);
  assign _zz_dataOut_payload_0_7465 = (_zz_dataOut_payload_0_7464 ? _zz_dataOut_payload_0_7441 : _zz_dataOut_payload_0_7453);
  assign _zz_dataOut_payload_0_7466 = (_zz_dataOut_payload_0_7464 ? _zz_dataOut_payload_0_7453 : _zz_dataOut_payload_0_7441);
  assign _zz_dataOut_payload_0_7467 = (_zz_dataOut_payload_0_7444 < _zz_dataOut_payload_0_7456);
  assign _zz_dataOut_payload_0_7468 = (_zz_dataOut_payload_0_7467 ? _zz_dataOut_payload_0_7444 : _zz_dataOut_payload_0_7456);
  assign _zz_dataOut_payload_0_7469 = (_zz_dataOut_payload_0_7467 ? _zz_dataOut_payload_0_7456 : _zz_dataOut_payload_0_7444);
  assign _zz_dataOut_payload_0_7470 = (_zz_dataOut_payload_0_7447 < _zz_dataOut_payload_0_7459);
  assign _zz_dataOut_payload_0_7471 = (_zz_dataOut_payload_0_7470 ? _zz_dataOut_payload_0_7447 : _zz_dataOut_payload_0_7459);
  assign _zz_dataOut_payload_0_7472 = (_zz_dataOut_payload_0_7470 ? _zz_dataOut_payload_0_7459 : _zz_dataOut_payload_0_7447);
  assign _zz_dataOut_payload_0_7473 = (_zz_dataOut_payload_0_7450 < _zz_dataOut_payload_0_7462);
  assign _zz_dataOut_payload_0_7474 = (_zz_dataOut_payload_0_7473 ? _zz_dataOut_payload_0_7450 : _zz_dataOut_payload_0_7462);
  assign _zz_dataOut_payload_0_7475 = (_zz_dataOut_payload_0_7473 ? _zz_dataOut_payload_0_7462 : _zz_dataOut_payload_0_7450);
  assign _zz_dataOut_payload_0_7476 = (_zz_dataOut_payload_0_7465 < _zz_dataOut_payload_0_7471);
  assign _zz_dataOut_payload_0_7477 = (_zz_dataOut_payload_0_7476 ? _zz_dataOut_payload_0_7465 : _zz_dataOut_payload_0_7471);
  assign _zz_dataOut_payload_0_7478 = (_zz_dataOut_payload_0_7476 ? _zz_dataOut_payload_0_7471 : _zz_dataOut_payload_0_7465);
  assign _zz_dataOut_payload_0_7479 = (_zz_dataOut_payload_0_7468 < _zz_dataOut_payload_0_7474);
  assign _zz_dataOut_payload_0_7480 = (_zz_dataOut_payload_0_7479 ? _zz_dataOut_payload_0_7468 : _zz_dataOut_payload_0_7474);
  assign _zz_dataOut_payload_0_7481 = (_zz_dataOut_payload_0_7479 ? _zz_dataOut_payload_0_7474 : _zz_dataOut_payload_0_7468);
  assign _zz_dataOut_payload_0_7482 = (_zz_dataOut_payload_0_7477 < _zz_dataOut_payload_0_7480);
  assign _zz_dataOut_payload_0_7483 = (_zz_dataOut_payload_0_7478 < _zz_dataOut_payload_0_7481);
  assign _zz_dataOut_payload_0_7488 = (_zz_dataOut_payload_0_7466 < _zz_dataOut_payload_0_7472);
  assign _zz_dataOut_payload_0_7489 = (_zz_dataOut_payload_0_7488 ? _zz_dataOut_payload_0_7466 : _zz_dataOut_payload_0_7472);
  assign _zz_dataOut_payload_0_7490 = (_zz_dataOut_payload_0_7488 ? _zz_dataOut_payload_0_7472 : _zz_dataOut_payload_0_7466);
  assign _zz_dataOut_payload_0_7491 = (_zz_dataOut_payload_0_7469 < _zz_dataOut_payload_0_7475);
  assign _zz_dataOut_payload_0_7492 = (_zz_dataOut_payload_0_7491 ? _zz_dataOut_payload_0_7469 : _zz_dataOut_payload_0_7475);
  assign _zz_dataOut_payload_0_7493 = (_zz_dataOut_payload_0_7491 ? _zz_dataOut_payload_0_7475 : _zz_dataOut_payload_0_7469);
  assign _zz_dataOut_payload_0_7494 = (_zz_dataOut_payload_0_7489 < _zz_dataOut_payload_0_7492);
  assign _zz_dataOut_payload_0_7495 = (_zz_dataOut_payload_0_7490 < _zz_dataOut_payload_0_7493);
  assign _zz_dataOut_payload_0_7508 = (_zz_dataOut_payload_0_7442 < _zz_dataOut_payload_0_7454);
  assign _zz_dataOut_payload_0_7509 = (_zz_dataOut_payload_0_7508 ? _zz_dataOut_payload_0_7442 : _zz_dataOut_payload_0_7454);
  assign _zz_dataOut_payload_0_7510 = (_zz_dataOut_payload_0_7508 ? _zz_dataOut_payload_0_7454 : _zz_dataOut_payload_0_7442);
  assign _zz_dataOut_payload_0_7511 = (_zz_dataOut_payload_0_7445 < _zz_dataOut_payload_0_7457);
  assign _zz_dataOut_payload_0_7512 = (_zz_dataOut_payload_0_7511 ? _zz_dataOut_payload_0_7445 : _zz_dataOut_payload_0_7457);
  assign _zz_dataOut_payload_0_7513 = (_zz_dataOut_payload_0_7511 ? _zz_dataOut_payload_0_7457 : _zz_dataOut_payload_0_7445);
  assign _zz_dataOut_payload_0_7514 = (_zz_dataOut_payload_0_7448 < _zz_dataOut_payload_0_7460);
  assign _zz_dataOut_payload_0_7515 = (_zz_dataOut_payload_0_7514 ? _zz_dataOut_payload_0_7448 : _zz_dataOut_payload_0_7460);
  assign _zz_dataOut_payload_0_7516 = (_zz_dataOut_payload_0_7514 ? _zz_dataOut_payload_0_7460 : _zz_dataOut_payload_0_7448);
  assign _zz_dataOut_payload_0_7517 = (_zz_dataOut_payload_0_7451 < _zz_dataOut_payload_0_7463);
  assign _zz_dataOut_payload_0_7518 = (_zz_dataOut_payload_0_7517 ? _zz_dataOut_payload_0_7451 : _zz_dataOut_payload_0_7463);
  assign _zz_dataOut_payload_0_7519 = (_zz_dataOut_payload_0_7517 ? _zz_dataOut_payload_0_7463 : _zz_dataOut_payload_0_7451);
  assign _zz_dataOut_payload_0_7520 = (_zz_dataOut_payload_0_7509 < _zz_dataOut_payload_0_7515);
  assign _zz_dataOut_payload_0_7521 = (_zz_dataOut_payload_0_7520 ? _zz_dataOut_payload_0_7509 : _zz_dataOut_payload_0_7515);
  assign _zz_dataOut_payload_0_7522 = (_zz_dataOut_payload_0_7520 ? _zz_dataOut_payload_0_7515 : _zz_dataOut_payload_0_7509);
  assign _zz_dataOut_payload_0_7523 = (_zz_dataOut_payload_0_7512 < _zz_dataOut_payload_0_7518);
  assign _zz_dataOut_payload_0_7524 = (_zz_dataOut_payload_0_7523 ? _zz_dataOut_payload_0_7512 : _zz_dataOut_payload_0_7518);
  assign _zz_dataOut_payload_0_7525 = (_zz_dataOut_payload_0_7523 ? _zz_dataOut_payload_0_7518 : _zz_dataOut_payload_0_7512);
  assign _zz_dataOut_payload_0_7526 = (_zz_dataOut_payload_0_7521 < _zz_dataOut_payload_0_7524);
  assign _zz_dataOut_payload_0_7527 = (_zz_dataOut_payload_0_7522 < _zz_dataOut_payload_0_7525);
  assign _zz_dataOut_payload_0_7532 = (_zz_dataOut_payload_0_7510 < _zz_dataOut_payload_0_7516);
  assign _zz_dataOut_payload_0_7533 = (_zz_dataOut_payload_0_7532 ? _zz_dataOut_payload_0_7510 : _zz_dataOut_payload_0_7516);
  assign _zz_dataOut_payload_0_7534 = (_zz_dataOut_payload_0_7532 ? _zz_dataOut_payload_0_7516 : _zz_dataOut_payload_0_7510);
  assign _zz_dataOut_payload_0_7535 = (_zz_dataOut_payload_0_7513 < _zz_dataOut_payload_0_7519);
  assign _zz_dataOut_payload_0_7536 = (_zz_dataOut_payload_0_7535 ? _zz_dataOut_payload_0_7513 : _zz_dataOut_payload_0_7519);
  assign _zz_dataOut_payload_0_7537 = (_zz_dataOut_payload_0_7535 ? _zz_dataOut_payload_0_7519 : _zz_dataOut_payload_0_7513);
  assign _zz_dataOut_payload_0_7538 = (_zz_dataOut_payload_0_7533 < _zz_dataOut_payload_0_7536);
  assign _zz_dataOut_payload_0_7539 = (_zz_dataOut_payload_0_7534 < _zz_dataOut_payload_0_7537);
  assign _zz_dataOut_payload_0_7568 = (_zz_dataOut_payload_0_7439 < _zz_dataOut_payload_0_7415);
  assign _zz_dataOut_payload_0_7569 = (_zz_dataOut_payload_0_7568 ? _zz_dataOut_payload_0_7439 : _zz_dataOut_payload_0_7415);
  assign _zz_dataOut_payload_0_7570 = (_zz_dataOut_payload_0_7568 ? _zz_dataOut_payload_0_7415 : _zz_dataOut_payload_0_7439);
  assign _zz_dataOut_payload_0_7571 = (_zz_dataOut_payload_0_7436 < _zz_dataOut_payload_0_7412);
  assign _zz_dataOut_payload_0_7572 = (_zz_dataOut_payload_0_7571 ? _zz_dataOut_payload_0_7436 : _zz_dataOut_payload_0_7412);
  assign _zz_dataOut_payload_0_7573 = (_zz_dataOut_payload_0_7571 ? _zz_dataOut_payload_0_7412 : _zz_dataOut_payload_0_7436);
  assign _zz_dataOut_payload_0_7574 = (_zz_dataOut_payload_0_7433 < _zz_dataOut_payload_0_7409);
  assign _zz_dataOut_payload_0_7575 = (_zz_dataOut_payload_0_7574 ? _zz_dataOut_payload_0_7433 : _zz_dataOut_payload_0_7409);
  assign _zz_dataOut_payload_0_7576 = (_zz_dataOut_payload_0_7574 ? _zz_dataOut_payload_0_7409 : _zz_dataOut_payload_0_7433);
  assign _zz_dataOut_payload_0_7577 = (_zz_dataOut_payload_0_7430 < _zz_dataOut_payload_0_7406);
  assign _zz_dataOut_payload_0_7578 = (_zz_dataOut_payload_0_7577 ? _zz_dataOut_payload_0_7430 : _zz_dataOut_payload_0_7406);
  assign _zz_dataOut_payload_0_7579 = (_zz_dataOut_payload_0_7577 ? _zz_dataOut_payload_0_7406 : _zz_dataOut_payload_0_7430);
  assign _zz_dataOut_payload_0_7580 = (_zz_dataOut_payload_0_7427 < _zz_dataOut_payload_0_7403);
  assign _zz_dataOut_payload_0_7581 = (_zz_dataOut_payload_0_7580 ? _zz_dataOut_payload_0_7427 : _zz_dataOut_payload_0_7403);
  assign _zz_dataOut_payload_0_7582 = (_zz_dataOut_payload_0_7580 ? _zz_dataOut_payload_0_7403 : _zz_dataOut_payload_0_7427);
  assign _zz_dataOut_payload_0_7583 = (_zz_dataOut_payload_0_7424 < _zz_dataOut_payload_0_7400);
  assign _zz_dataOut_payload_0_7584 = (_zz_dataOut_payload_0_7583 ? _zz_dataOut_payload_0_7424 : _zz_dataOut_payload_0_7400);
  assign _zz_dataOut_payload_0_7585 = (_zz_dataOut_payload_0_7583 ? _zz_dataOut_payload_0_7400 : _zz_dataOut_payload_0_7424);
  assign _zz_dataOut_payload_0_7586 = (_zz_dataOut_payload_0_7421 < _zz_dataOut_payload_0_7397);
  assign _zz_dataOut_payload_0_7587 = (_zz_dataOut_payload_0_7586 ? _zz_dataOut_payload_0_7421 : _zz_dataOut_payload_0_7397);
  assign _zz_dataOut_payload_0_7588 = (_zz_dataOut_payload_0_7586 ? _zz_dataOut_payload_0_7397 : _zz_dataOut_payload_0_7421);
  assign _zz_dataOut_payload_0_7589 = (_zz_dataOut_payload_0_7418 < _zz_dataOut_payload_0_7394);
  assign _zz_dataOut_payload_0_7590 = (_zz_dataOut_payload_0_7589 ? _zz_dataOut_payload_0_7418 : _zz_dataOut_payload_0_7394);
  assign _zz_dataOut_payload_0_7591 = (_zz_dataOut_payload_0_7589 ? _zz_dataOut_payload_0_7394 : _zz_dataOut_payload_0_7418);
  assign _zz_dataOut_payload_0_7592 = (_zz_dataOut_payload_0_7569 < _zz_dataOut_payload_0_7581);
  assign _zz_dataOut_payload_0_7593 = (_zz_dataOut_payload_0_7592 ? _zz_dataOut_payload_0_7569 : _zz_dataOut_payload_0_7581);
  assign _zz_dataOut_payload_0_7594 = (_zz_dataOut_payload_0_7592 ? _zz_dataOut_payload_0_7581 : _zz_dataOut_payload_0_7569);
  assign _zz_dataOut_payload_0_7595 = (_zz_dataOut_payload_0_7572 < _zz_dataOut_payload_0_7584);
  assign _zz_dataOut_payload_0_7596 = (_zz_dataOut_payload_0_7595 ? _zz_dataOut_payload_0_7572 : _zz_dataOut_payload_0_7584);
  assign _zz_dataOut_payload_0_7597 = (_zz_dataOut_payload_0_7595 ? _zz_dataOut_payload_0_7584 : _zz_dataOut_payload_0_7572);
  assign _zz_dataOut_payload_0_7598 = (_zz_dataOut_payload_0_7575 < _zz_dataOut_payload_0_7587);
  assign _zz_dataOut_payload_0_7599 = (_zz_dataOut_payload_0_7598 ? _zz_dataOut_payload_0_7575 : _zz_dataOut_payload_0_7587);
  assign _zz_dataOut_payload_0_7600 = (_zz_dataOut_payload_0_7598 ? _zz_dataOut_payload_0_7587 : _zz_dataOut_payload_0_7575);
  assign _zz_dataOut_payload_0_7601 = (_zz_dataOut_payload_0_7578 < _zz_dataOut_payload_0_7590);
  assign _zz_dataOut_payload_0_7602 = (_zz_dataOut_payload_0_7601 ? _zz_dataOut_payload_0_7578 : _zz_dataOut_payload_0_7590);
  assign _zz_dataOut_payload_0_7603 = (_zz_dataOut_payload_0_7601 ? _zz_dataOut_payload_0_7590 : _zz_dataOut_payload_0_7578);
  assign _zz_dataOut_payload_0_7604 = (_zz_dataOut_payload_0_7593 < _zz_dataOut_payload_0_7599);
  assign _zz_dataOut_payload_0_7605 = (_zz_dataOut_payload_0_7604 ? _zz_dataOut_payload_0_7593 : _zz_dataOut_payload_0_7599);
  assign _zz_dataOut_payload_0_7606 = (_zz_dataOut_payload_0_7604 ? _zz_dataOut_payload_0_7599 : _zz_dataOut_payload_0_7593);
  assign _zz_dataOut_payload_0_7607 = (_zz_dataOut_payload_0_7596 < _zz_dataOut_payload_0_7602);
  assign _zz_dataOut_payload_0_7608 = (_zz_dataOut_payload_0_7607 ? _zz_dataOut_payload_0_7596 : _zz_dataOut_payload_0_7602);
  assign _zz_dataOut_payload_0_7609 = (_zz_dataOut_payload_0_7607 ? _zz_dataOut_payload_0_7602 : _zz_dataOut_payload_0_7596);
  assign _zz_dataOut_payload_0_7610 = (_zz_dataOut_payload_0_7605 < _zz_dataOut_payload_0_7608);
  assign _zz_dataOut_payload_0_7611 = (_zz_dataOut_payload_0_7606 < _zz_dataOut_payload_0_7609);
  assign _zz_dataOut_payload_0_7616 = (_zz_dataOut_payload_0_7594 < _zz_dataOut_payload_0_7600);
  assign _zz_dataOut_payload_0_7617 = (_zz_dataOut_payload_0_7616 ? _zz_dataOut_payload_0_7594 : _zz_dataOut_payload_0_7600);
  assign _zz_dataOut_payload_0_7618 = (_zz_dataOut_payload_0_7616 ? _zz_dataOut_payload_0_7600 : _zz_dataOut_payload_0_7594);
  assign _zz_dataOut_payload_0_7619 = (_zz_dataOut_payload_0_7597 < _zz_dataOut_payload_0_7603);
  assign _zz_dataOut_payload_0_7620 = (_zz_dataOut_payload_0_7619 ? _zz_dataOut_payload_0_7597 : _zz_dataOut_payload_0_7603);
  assign _zz_dataOut_payload_0_7621 = (_zz_dataOut_payload_0_7619 ? _zz_dataOut_payload_0_7603 : _zz_dataOut_payload_0_7597);
  assign _zz_dataOut_payload_0_7622 = (_zz_dataOut_payload_0_7617 < _zz_dataOut_payload_0_7620);
  assign _zz_dataOut_payload_0_7623 = (_zz_dataOut_payload_0_7618 < _zz_dataOut_payload_0_7621);
  assign _zz_dataOut_payload_0_7636 = (_zz_dataOut_payload_0_7570 < _zz_dataOut_payload_0_7582);
  assign _zz_dataOut_payload_0_7637 = (_zz_dataOut_payload_0_7636 ? _zz_dataOut_payload_0_7570 : _zz_dataOut_payload_0_7582);
  assign _zz_dataOut_payload_0_7638 = (_zz_dataOut_payload_0_7636 ? _zz_dataOut_payload_0_7582 : _zz_dataOut_payload_0_7570);
  assign _zz_dataOut_payload_0_7639 = (_zz_dataOut_payload_0_7573 < _zz_dataOut_payload_0_7585);
  assign _zz_dataOut_payload_0_7640 = (_zz_dataOut_payload_0_7639 ? _zz_dataOut_payload_0_7573 : _zz_dataOut_payload_0_7585);
  assign _zz_dataOut_payload_0_7641 = (_zz_dataOut_payload_0_7639 ? _zz_dataOut_payload_0_7585 : _zz_dataOut_payload_0_7573);
  assign _zz_dataOut_payload_0_7642 = (_zz_dataOut_payload_0_7576 < _zz_dataOut_payload_0_7588);
  assign _zz_dataOut_payload_0_7643 = (_zz_dataOut_payload_0_7642 ? _zz_dataOut_payload_0_7576 : _zz_dataOut_payload_0_7588);
  assign _zz_dataOut_payload_0_7644 = (_zz_dataOut_payload_0_7642 ? _zz_dataOut_payload_0_7588 : _zz_dataOut_payload_0_7576);
  assign _zz_dataOut_payload_0_7645 = (_zz_dataOut_payload_0_7579 < _zz_dataOut_payload_0_7591);
  assign _zz_dataOut_payload_0_7646 = (_zz_dataOut_payload_0_7645 ? _zz_dataOut_payload_0_7579 : _zz_dataOut_payload_0_7591);
  assign _zz_dataOut_payload_0_7647 = (_zz_dataOut_payload_0_7645 ? _zz_dataOut_payload_0_7591 : _zz_dataOut_payload_0_7579);
  assign _zz_dataOut_payload_0_7648 = (_zz_dataOut_payload_0_7637 < _zz_dataOut_payload_0_7643);
  assign _zz_dataOut_payload_0_7649 = (_zz_dataOut_payload_0_7648 ? _zz_dataOut_payload_0_7637 : _zz_dataOut_payload_0_7643);
  assign _zz_dataOut_payload_0_7650 = (_zz_dataOut_payload_0_7648 ? _zz_dataOut_payload_0_7643 : _zz_dataOut_payload_0_7637);
  assign _zz_dataOut_payload_0_7651 = (_zz_dataOut_payload_0_7640 < _zz_dataOut_payload_0_7646);
  assign _zz_dataOut_payload_0_7652 = (_zz_dataOut_payload_0_7651 ? _zz_dataOut_payload_0_7640 : _zz_dataOut_payload_0_7646);
  assign _zz_dataOut_payload_0_7653 = (_zz_dataOut_payload_0_7651 ? _zz_dataOut_payload_0_7646 : _zz_dataOut_payload_0_7640);
  assign _zz_dataOut_payload_0_7654 = (_zz_dataOut_payload_0_7649 < _zz_dataOut_payload_0_7652);
  assign _zz_dataOut_payload_0_7655 = (_zz_dataOut_payload_0_7650 < _zz_dataOut_payload_0_7653);
  assign _zz_dataOut_payload_0_7660 = (_zz_dataOut_payload_0_7638 < _zz_dataOut_payload_0_7644);
  assign _zz_dataOut_payload_0_7661 = (_zz_dataOut_payload_0_7660 ? _zz_dataOut_payload_0_7638 : _zz_dataOut_payload_0_7644);
  assign _zz_dataOut_payload_0_7662 = (_zz_dataOut_payload_0_7660 ? _zz_dataOut_payload_0_7644 : _zz_dataOut_payload_0_7638);
  assign _zz_dataOut_payload_0_7663 = (_zz_dataOut_payload_0_7641 < _zz_dataOut_payload_0_7647);
  assign _zz_dataOut_payload_0_7664 = (_zz_dataOut_payload_0_7663 ? _zz_dataOut_payload_0_7641 : _zz_dataOut_payload_0_7647);
  assign _zz_dataOut_payload_0_7665 = (_zz_dataOut_payload_0_7663 ? _zz_dataOut_payload_0_7647 : _zz_dataOut_payload_0_7641);
  assign _zz_dataOut_payload_0_7666 = (_zz_dataOut_payload_0_7661 < _zz_dataOut_payload_0_7664);
  assign _zz_dataOut_payload_0_7667 = (_zz_dataOut_payload_0_7662 < _zz_dataOut_payload_0_7665);
  assign _zz_dataOut_payload_0_7728 = (_zz_dataOut_payload_0_5344 < _zz_dataOut_payload_0_5375);
  assign _zz_dataOut_payload_0_7729 = (_zz_dataOut_payload_0_7728 ? _zz_dataOut_payload_0_5344 : _zz_dataOut_payload_0_5375);
  assign _zz_dataOut_payload_0_7730 = (_zz_dataOut_payload_0_7728 ? _zz_dataOut_payload_0_5375 : _zz_dataOut_payload_0_5344);
  assign _zz_dataOut_payload_0_7731 = (_zz_dataOut_payload_0_5345 < _zz_dataOut_payload_0_5374);
  assign _zz_dataOut_payload_0_7732 = (_zz_dataOut_payload_0_7731 ? _zz_dataOut_payload_0_5345 : _zz_dataOut_payload_0_5374);
  assign _zz_dataOut_payload_0_7733 = (_zz_dataOut_payload_0_7731 ? _zz_dataOut_payload_0_5374 : _zz_dataOut_payload_0_5345);
  assign _zz_dataOut_payload_0_7734 = (_zz_dataOut_payload_0_5346 < _zz_dataOut_payload_0_5373);
  assign _zz_dataOut_payload_0_7735 = (_zz_dataOut_payload_0_7734 ? _zz_dataOut_payload_0_5346 : _zz_dataOut_payload_0_5373);
  assign _zz_dataOut_payload_0_7736 = (_zz_dataOut_payload_0_7734 ? _zz_dataOut_payload_0_5373 : _zz_dataOut_payload_0_5346);
  assign _zz_dataOut_payload_0_7737 = (_zz_dataOut_payload_0_5347 < _zz_dataOut_payload_0_5372);
  assign _zz_dataOut_payload_0_7738 = (_zz_dataOut_payload_0_7737 ? _zz_dataOut_payload_0_5347 : _zz_dataOut_payload_0_5372);
  assign _zz_dataOut_payload_0_7739 = (_zz_dataOut_payload_0_7737 ? _zz_dataOut_payload_0_5372 : _zz_dataOut_payload_0_5347);
  assign _zz_dataOut_payload_0_7740 = (_zz_dataOut_payload_0_5348 < _zz_dataOut_payload_0_5371);
  assign _zz_dataOut_payload_0_7741 = (_zz_dataOut_payload_0_7740 ? _zz_dataOut_payload_0_5348 : _zz_dataOut_payload_0_5371);
  assign _zz_dataOut_payload_0_7742 = (_zz_dataOut_payload_0_7740 ? _zz_dataOut_payload_0_5371 : _zz_dataOut_payload_0_5348);
  assign _zz_dataOut_payload_0_7743 = (_zz_dataOut_payload_0_5349 < _zz_dataOut_payload_0_5370);
  assign _zz_dataOut_payload_0_7744 = (_zz_dataOut_payload_0_7743 ? _zz_dataOut_payload_0_5349 : _zz_dataOut_payload_0_5370);
  assign _zz_dataOut_payload_0_7745 = (_zz_dataOut_payload_0_7743 ? _zz_dataOut_payload_0_5370 : _zz_dataOut_payload_0_5349);
  assign _zz_dataOut_payload_0_7746 = (_zz_dataOut_payload_0_5350 < _zz_dataOut_payload_0_5369);
  assign _zz_dataOut_payload_0_7747 = (_zz_dataOut_payload_0_7746 ? _zz_dataOut_payload_0_5350 : _zz_dataOut_payload_0_5369);
  assign _zz_dataOut_payload_0_7748 = (_zz_dataOut_payload_0_7746 ? _zz_dataOut_payload_0_5369 : _zz_dataOut_payload_0_5350);
  assign _zz_dataOut_payload_0_7749 = (_zz_dataOut_payload_0_5351 < _zz_dataOut_payload_0_5368);
  assign _zz_dataOut_payload_0_7750 = (_zz_dataOut_payload_0_7749 ? _zz_dataOut_payload_0_5351 : _zz_dataOut_payload_0_5368);
  assign _zz_dataOut_payload_0_7751 = (_zz_dataOut_payload_0_7749 ? _zz_dataOut_payload_0_5368 : _zz_dataOut_payload_0_5351);
  assign _zz_dataOut_payload_0_7752 = (_zz_dataOut_payload_0_5352 < _zz_dataOut_payload_0_5367);
  assign _zz_dataOut_payload_0_7753 = (_zz_dataOut_payload_0_7752 ? _zz_dataOut_payload_0_5352 : _zz_dataOut_payload_0_5367);
  assign _zz_dataOut_payload_0_7754 = (_zz_dataOut_payload_0_7752 ? _zz_dataOut_payload_0_5367 : _zz_dataOut_payload_0_5352);
  assign _zz_dataOut_payload_0_7755 = (_zz_dataOut_payload_0_5353 < _zz_dataOut_payload_0_5366);
  assign _zz_dataOut_payload_0_7756 = (_zz_dataOut_payload_0_7755 ? _zz_dataOut_payload_0_5353 : _zz_dataOut_payload_0_5366);
  assign _zz_dataOut_payload_0_7757 = (_zz_dataOut_payload_0_7755 ? _zz_dataOut_payload_0_5366 : _zz_dataOut_payload_0_5353);
  assign _zz_dataOut_payload_0_7758 = (_zz_dataOut_payload_0_5354 < _zz_dataOut_payload_0_5365);
  assign _zz_dataOut_payload_0_7759 = (_zz_dataOut_payload_0_7758 ? _zz_dataOut_payload_0_5354 : _zz_dataOut_payload_0_5365);
  assign _zz_dataOut_payload_0_7760 = (_zz_dataOut_payload_0_7758 ? _zz_dataOut_payload_0_5365 : _zz_dataOut_payload_0_5354);
  assign _zz_dataOut_payload_0_7761 = (_zz_dataOut_payload_0_5355 < _zz_dataOut_payload_0_5364);
  assign _zz_dataOut_payload_0_7762 = (_zz_dataOut_payload_0_7761 ? _zz_dataOut_payload_0_5355 : _zz_dataOut_payload_0_5364);
  assign _zz_dataOut_payload_0_7763 = (_zz_dataOut_payload_0_7761 ? _zz_dataOut_payload_0_5364 : _zz_dataOut_payload_0_5355);
  assign _zz_dataOut_payload_0_7764 = (_zz_dataOut_payload_0_5356 < _zz_dataOut_payload_0_5363);
  assign _zz_dataOut_payload_0_7765 = (_zz_dataOut_payload_0_7764 ? _zz_dataOut_payload_0_5356 : _zz_dataOut_payload_0_5363);
  assign _zz_dataOut_payload_0_7766 = (_zz_dataOut_payload_0_7764 ? _zz_dataOut_payload_0_5363 : _zz_dataOut_payload_0_5356);
  assign _zz_dataOut_payload_0_7767 = (_zz_dataOut_payload_0_5357 < _zz_dataOut_payload_0_5362);
  assign _zz_dataOut_payload_0_7768 = (_zz_dataOut_payload_0_7767 ? _zz_dataOut_payload_0_5357 : _zz_dataOut_payload_0_5362);
  assign _zz_dataOut_payload_0_7769 = (_zz_dataOut_payload_0_7767 ? _zz_dataOut_payload_0_5362 : _zz_dataOut_payload_0_5357);
  assign _zz_dataOut_payload_0_7770 = (_zz_dataOut_payload_0_5358 < _zz_dataOut_payload_0_5361);
  assign _zz_dataOut_payload_0_7771 = (_zz_dataOut_payload_0_7770 ? _zz_dataOut_payload_0_5358 : _zz_dataOut_payload_0_5361);
  assign _zz_dataOut_payload_0_7772 = (_zz_dataOut_payload_0_7770 ? _zz_dataOut_payload_0_5361 : _zz_dataOut_payload_0_5358);
  assign _zz_dataOut_payload_0_7773 = (_zz_dataOut_payload_0_5359 < _zz_dataOut_payload_0_5360);
  assign _zz_dataOut_payload_0_7774 = (_zz_dataOut_payload_0_7773 ? _zz_dataOut_payload_0_5359 : _zz_dataOut_payload_0_5360);
  assign _zz_dataOut_payload_0_7775 = (_zz_dataOut_payload_0_7773 ? _zz_dataOut_payload_0_5360 : _zz_dataOut_payload_0_5359);
  assign _zz_dataOut_payload_0_7776 = (_zz_dataOut_payload_0_7729 < _zz_dataOut_payload_0_7753);
  assign _zz_dataOut_payload_0_7777 = (_zz_dataOut_payload_0_7776 ? _zz_dataOut_payload_0_7729 : _zz_dataOut_payload_0_7753);
  assign _zz_dataOut_payload_0_7778 = (_zz_dataOut_payload_0_7776 ? _zz_dataOut_payload_0_7753 : _zz_dataOut_payload_0_7729);
  assign _zz_dataOut_payload_0_7779 = (_zz_dataOut_payload_0_7732 < _zz_dataOut_payload_0_7756);
  assign _zz_dataOut_payload_0_7780 = (_zz_dataOut_payload_0_7779 ? _zz_dataOut_payload_0_7732 : _zz_dataOut_payload_0_7756);
  assign _zz_dataOut_payload_0_7781 = (_zz_dataOut_payload_0_7779 ? _zz_dataOut_payload_0_7756 : _zz_dataOut_payload_0_7732);
  assign _zz_dataOut_payload_0_7782 = (_zz_dataOut_payload_0_7735 < _zz_dataOut_payload_0_7759);
  assign _zz_dataOut_payload_0_7783 = (_zz_dataOut_payload_0_7782 ? _zz_dataOut_payload_0_7735 : _zz_dataOut_payload_0_7759);
  assign _zz_dataOut_payload_0_7784 = (_zz_dataOut_payload_0_7782 ? _zz_dataOut_payload_0_7759 : _zz_dataOut_payload_0_7735);
  assign _zz_dataOut_payload_0_7785 = (_zz_dataOut_payload_0_7738 < _zz_dataOut_payload_0_7762);
  assign _zz_dataOut_payload_0_7786 = (_zz_dataOut_payload_0_7785 ? _zz_dataOut_payload_0_7738 : _zz_dataOut_payload_0_7762);
  assign _zz_dataOut_payload_0_7787 = (_zz_dataOut_payload_0_7785 ? _zz_dataOut_payload_0_7762 : _zz_dataOut_payload_0_7738);
  assign _zz_dataOut_payload_0_7788 = (_zz_dataOut_payload_0_7741 < _zz_dataOut_payload_0_7765);
  assign _zz_dataOut_payload_0_7789 = (_zz_dataOut_payload_0_7788 ? _zz_dataOut_payload_0_7741 : _zz_dataOut_payload_0_7765);
  assign _zz_dataOut_payload_0_7790 = (_zz_dataOut_payload_0_7788 ? _zz_dataOut_payload_0_7765 : _zz_dataOut_payload_0_7741);
  assign _zz_dataOut_payload_0_7791 = (_zz_dataOut_payload_0_7744 < _zz_dataOut_payload_0_7768);
  assign _zz_dataOut_payload_0_7792 = (_zz_dataOut_payload_0_7791 ? _zz_dataOut_payload_0_7744 : _zz_dataOut_payload_0_7768);
  assign _zz_dataOut_payload_0_7793 = (_zz_dataOut_payload_0_7791 ? _zz_dataOut_payload_0_7768 : _zz_dataOut_payload_0_7744);
  assign _zz_dataOut_payload_0_7794 = (_zz_dataOut_payload_0_7747 < _zz_dataOut_payload_0_7771);
  assign _zz_dataOut_payload_0_7795 = (_zz_dataOut_payload_0_7794 ? _zz_dataOut_payload_0_7747 : _zz_dataOut_payload_0_7771);
  assign _zz_dataOut_payload_0_7796 = (_zz_dataOut_payload_0_7794 ? _zz_dataOut_payload_0_7771 : _zz_dataOut_payload_0_7747);
  assign _zz_dataOut_payload_0_7797 = (_zz_dataOut_payload_0_7750 < _zz_dataOut_payload_0_7774);
  assign _zz_dataOut_payload_0_7798 = (_zz_dataOut_payload_0_7797 ? _zz_dataOut_payload_0_7750 : _zz_dataOut_payload_0_7774);
  assign _zz_dataOut_payload_0_7799 = (_zz_dataOut_payload_0_7797 ? _zz_dataOut_payload_0_7774 : _zz_dataOut_payload_0_7750);
  assign _zz_dataOut_payload_0_7800 = (_zz_dataOut_payload_0_7777 < _zz_dataOut_payload_0_7789);
  assign _zz_dataOut_payload_0_7801 = (_zz_dataOut_payload_0_7800 ? _zz_dataOut_payload_0_7777 : _zz_dataOut_payload_0_7789);
  assign _zz_dataOut_payload_0_7802 = (_zz_dataOut_payload_0_7800 ? _zz_dataOut_payload_0_7789 : _zz_dataOut_payload_0_7777);
  assign _zz_dataOut_payload_0_7803 = (_zz_dataOut_payload_0_7780 < _zz_dataOut_payload_0_7792);
  assign _zz_dataOut_payload_0_7804 = (_zz_dataOut_payload_0_7803 ? _zz_dataOut_payload_0_7780 : _zz_dataOut_payload_0_7792);
  assign _zz_dataOut_payload_0_7805 = (_zz_dataOut_payload_0_7803 ? _zz_dataOut_payload_0_7792 : _zz_dataOut_payload_0_7780);
  assign _zz_dataOut_payload_0_7806 = (_zz_dataOut_payload_0_7783 < _zz_dataOut_payload_0_7795);
  assign _zz_dataOut_payload_0_7807 = (_zz_dataOut_payload_0_7806 ? _zz_dataOut_payload_0_7783 : _zz_dataOut_payload_0_7795);
  assign _zz_dataOut_payload_0_7808 = (_zz_dataOut_payload_0_7806 ? _zz_dataOut_payload_0_7795 : _zz_dataOut_payload_0_7783);
  assign _zz_dataOut_payload_0_7809 = (_zz_dataOut_payload_0_7786 < _zz_dataOut_payload_0_7798);
  assign _zz_dataOut_payload_0_7810 = (_zz_dataOut_payload_0_7809 ? _zz_dataOut_payload_0_7786 : _zz_dataOut_payload_0_7798);
  assign _zz_dataOut_payload_0_7811 = (_zz_dataOut_payload_0_7809 ? _zz_dataOut_payload_0_7798 : _zz_dataOut_payload_0_7786);
  assign _zz_dataOut_payload_0_7812 = (_zz_dataOut_payload_0_7801 < _zz_dataOut_payload_0_7807);
  assign _zz_dataOut_payload_0_7813 = (_zz_dataOut_payload_0_7812 ? _zz_dataOut_payload_0_7801 : _zz_dataOut_payload_0_7807);
  assign _zz_dataOut_payload_0_7814 = (_zz_dataOut_payload_0_7812 ? _zz_dataOut_payload_0_7807 : _zz_dataOut_payload_0_7801);
  assign _zz_dataOut_payload_0_7815 = (_zz_dataOut_payload_0_7804 < _zz_dataOut_payload_0_7810);
  assign _zz_dataOut_payload_0_7816 = (_zz_dataOut_payload_0_7815 ? _zz_dataOut_payload_0_7804 : _zz_dataOut_payload_0_7810);
  assign _zz_dataOut_payload_0_7817 = (_zz_dataOut_payload_0_7815 ? _zz_dataOut_payload_0_7810 : _zz_dataOut_payload_0_7804);
  assign _zz_dataOut_payload_0_7818 = (_zz_dataOut_payload_0_7813 < _zz_dataOut_payload_0_7816);
  assign _zz_dataOut_payload_0_7819 = (_zz_dataOut_payload_0_7814 < _zz_dataOut_payload_0_7817);
  assign _zz_dataOut_payload_0_7824 = (_zz_dataOut_payload_0_7802 < _zz_dataOut_payload_0_7808);
  assign _zz_dataOut_payload_0_7825 = (_zz_dataOut_payload_0_7824 ? _zz_dataOut_payload_0_7802 : _zz_dataOut_payload_0_7808);
  assign _zz_dataOut_payload_0_7826 = (_zz_dataOut_payload_0_7824 ? _zz_dataOut_payload_0_7808 : _zz_dataOut_payload_0_7802);
  assign _zz_dataOut_payload_0_7827 = (_zz_dataOut_payload_0_7805 < _zz_dataOut_payload_0_7811);
  assign _zz_dataOut_payload_0_7828 = (_zz_dataOut_payload_0_7827 ? _zz_dataOut_payload_0_7805 : _zz_dataOut_payload_0_7811);
  assign _zz_dataOut_payload_0_7829 = (_zz_dataOut_payload_0_7827 ? _zz_dataOut_payload_0_7811 : _zz_dataOut_payload_0_7805);
  assign _zz_dataOut_payload_0_7830 = (_zz_dataOut_payload_0_7825 < _zz_dataOut_payload_0_7828);
  assign _zz_dataOut_payload_0_7831 = (_zz_dataOut_payload_0_7826 < _zz_dataOut_payload_0_7829);
  assign _zz_dataOut_payload_0_7844 = (_zz_dataOut_payload_0_7778 < _zz_dataOut_payload_0_7790);
  assign _zz_dataOut_payload_0_7845 = (_zz_dataOut_payload_0_7844 ? _zz_dataOut_payload_0_7778 : _zz_dataOut_payload_0_7790);
  assign _zz_dataOut_payload_0_7846 = (_zz_dataOut_payload_0_7844 ? _zz_dataOut_payload_0_7790 : _zz_dataOut_payload_0_7778);
  assign _zz_dataOut_payload_0_7847 = (_zz_dataOut_payload_0_7781 < _zz_dataOut_payload_0_7793);
  assign _zz_dataOut_payload_0_7848 = (_zz_dataOut_payload_0_7847 ? _zz_dataOut_payload_0_7781 : _zz_dataOut_payload_0_7793);
  assign _zz_dataOut_payload_0_7849 = (_zz_dataOut_payload_0_7847 ? _zz_dataOut_payload_0_7793 : _zz_dataOut_payload_0_7781);
  assign _zz_dataOut_payload_0_7850 = (_zz_dataOut_payload_0_7784 < _zz_dataOut_payload_0_7796);
  assign _zz_dataOut_payload_0_7851 = (_zz_dataOut_payload_0_7850 ? _zz_dataOut_payload_0_7784 : _zz_dataOut_payload_0_7796);
  assign _zz_dataOut_payload_0_7852 = (_zz_dataOut_payload_0_7850 ? _zz_dataOut_payload_0_7796 : _zz_dataOut_payload_0_7784);
  assign _zz_dataOut_payload_0_7853 = (_zz_dataOut_payload_0_7787 < _zz_dataOut_payload_0_7799);
  assign _zz_dataOut_payload_0_7854 = (_zz_dataOut_payload_0_7853 ? _zz_dataOut_payload_0_7787 : _zz_dataOut_payload_0_7799);
  assign _zz_dataOut_payload_0_7855 = (_zz_dataOut_payload_0_7853 ? _zz_dataOut_payload_0_7799 : _zz_dataOut_payload_0_7787);
  assign _zz_dataOut_payload_0_7856 = (_zz_dataOut_payload_0_7845 < _zz_dataOut_payload_0_7851);
  assign _zz_dataOut_payload_0_7857 = (_zz_dataOut_payload_0_7856 ? _zz_dataOut_payload_0_7845 : _zz_dataOut_payload_0_7851);
  assign _zz_dataOut_payload_0_7858 = (_zz_dataOut_payload_0_7856 ? _zz_dataOut_payload_0_7851 : _zz_dataOut_payload_0_7845);
  assign _zz_dataOut_payload_0_7859 = (_zz_dataOut_payload_0_7848 < _zz_dataOut_payload_0_7854);
  assign _zz_dataOut_payload_0_7860 = (_zz_dataOut_payload_0_7859 ? _zz_dataOut_payload_0_7848 : _zz_dataOut_payload_0_7854);
  assign _zz_dataOut_payload_0_7861 = (_zz_dataOut_payload_0_7859 ? _zz_dataOut_payload_0_7854 : _zz_dataOut_payload_0_7848);
  assign _zz_dataOut_payload_0_7862 = (_zz_dataOut_payload_0_7857 < _zz_dataOut_payload_0_7860);
  assign _zz_dataOut_payload_0_7863 = (_zz_dataOut_payload_0_7858 < _zz_dataOut_payload_0_7861);
  assign _zz_dataOut_payload_0_7868 = (_zz_dataOut_payload_0_7846 < _zz_dataOut_payload_0_7852);
  assign _zz_dataOut_payload_0_7869 = (_zz_dataOut_payload_0_7868 ? _zz_dataOut_payload_0_7846 : _zz_dataOut_payload_0_7852);
  assign _zz_dataOut_payload_0_7870 = (_zz_dataOut_payload_0_7868 ? _zz_dataOut_payload_0_7852 : _zz_dataOut_payload_0_7846);
  assign _zz_dataOut_payload_0_7871 = (_zz_dataOut_payload_0_7849 < _zz_dataOut_payload_0_7855);
  assign _zz_dataOut_payload_0_7872 = (_zz_dataOut_payload_0_7871 ? _zz_dataOut_payload_0_7849 : _zz_dataOut_payload_0_7855);
  assign _zz_dataOut_payload_0_7873 = (_zz_dataOut_payload_0_7871 ? _zz_dataOut_payload_0_7855 : _zz_dataOut_payload_0_7849);
  assign _zz_dataOut_payload_0_7874 = (_zz_dataOut_payload_0_7869 < _zz_dataOut_payload_0_7872);
  assign _zz_dataOut_payload_0_7875 = (_zz_dataOut_payload_0_7870 < _zz_dataOut_payload_0_7873);
  assign _zz_dataOut_payload_0_7904 = (_zz_dataOut_payload_0_7775 < _zz_dataOut_payload_0_7751);
  assign _zz_dataOut_payload_0_7905 = (_zz_dataOut_payload_0_7904 ? _zz_dataOut_payload_0_7775 : _zz_dataOut_payload_0_7751);
  assign _zz_dataOut_payload_0_7906 = (_zz_dataOut_payload_0_7904 ? _zz_dataOut_payload_0_7751 : _zz_dataOut_payload_0_7775);
  assign _zz_dataOut_payload_0_7907 = (_zz_dataOut_payload_0_7772 < _zz_dataOut_payload_0_7748);
  assign _zz_dataOut_payload_0_7908 = (_zz_dataOut_payload_0_7907 ? _zz_dataOut_payload_0_7772 : _zz_dataOut_payload_0_7748);
  assign _zz_dataOut_payload_0_7909 = (_zz_dataOut_payload_0_7907 ? _zz_dataOut_payload_0_7748 : _zz_dataOut_payload_0_7772);
  assign _zz_dataOut_payload_0_7910 = (_zz_dataOut_payload_0_7769 < _zz_dataOut_payload_0_7745);
  assign _zz_dataOut_payload_0_7911 = (_zz_dataOut_payload_0_7910 ? _zz_dataOut_payload_0_7769 : _zz_dataOut_payload_0_7745);
  assign _zz_dataOut_payload_0_7912 = (_zz_dataOut_payload_0_7910 ? _zz_dataOut_payload_0_7745 : _zz_dataOut_payload_0_7769);
  assign _zz_dataOut_payload_0_7913 = (_zz_dataOut_payload_0_7766 < _zz_dataOut_payload_0_7742);
  assign _zz_dataOut_payload_0_7914 = (_zz_dataOut_payload_0_7913 ? _zz_dataOut_payload_0_7766 : _zz_dataOut_payload_0_7742);
  assign _zz_dataOut_payload_0_7915 = (_zz_dataOut_payload_0_7913 ? _zz_dataOut_payload_0_7742 : _zz_dataOut_payload_0_7766);
  assign _zz_dataOut_payload_0_7916 = (_zz_dataOut_payload_0_7763 < _zz_dataOut_payload_0_7739);
  assign _zz_dataOut_payload_0_7917 = (_zz_dataOut_payload_0_7916 ? _zz_dataOut_payload_0_7763 : _zz_dataOut_payload_0_7739);
  assign _zz_dataOut_payload_0_7918 = (_zz_dataOut_payload_0_7916 ? _zz_dataOut_payload_0_7739 : _zz_dataOut_payload_0_7763);
  assign _zz_dataOut_payload_0_7919 = (_zz_dataOut_payload_0_7760 < _zz_dataOut_payload_0_7736);
  assign _zz_dataOut_payload_0_7920 = (_zz_dataOut_payload_0_7919 ? _zz_dataOut_payload_0_7760 : _zz_dataOut_payload_0_7736);
  assign _zz_dataOut_payload_0_7921 = (_zz_dataOut_payload_0_7919 ? _zz_dataOut_payload_0_7736 : _zz_dataOut_payload_0_7760);
  assign _zz_dataOut_payload_0_7922 = (_zz_dataOut_payload_0_7757 < _zz_dataOut_payload_0_7733);
  assign _zz_dataOut_payload_0_7923 = (_zz_dataOut_payload_0_7922 ? _zz_dataOut_payload_0_7757 : _zz_dataOut_payload_0_7733);
  assign _zz_dataOut_payload_0_7924 = (_zz_dataOut_payload_0_7922 ? _zz_dataOut_payload_0_7733 : _zz_dataOut_payload_0_7757);
  assign _zz_dataOut_payload_0_7925 = (_zz_dataOut_payload_0_7754 < _zz_dataOut_payload_0_7730);
  assign _zz_dataOut_payload_0_7926 = (_zz_dataOut_payload_0_7925 ? _zz_dataOut_payload_0_7754 : _zz_dataOut_payload_0_7730);
  assign _zz_dataOut_payload_0_7927 = (_zz_dataOut_payload_0_7925 ? _zz_dataOut_payload_0_7730 : _zz_dataOut_payload_0_7754);
  assign _zz_dataOut_payload_0_7928 = (_zz_dataOut_payload_0_7905 < _zz_dataOut_payload_0_7917);
  assign _zz_dataOut_payload_0_7929 = (_zz_dataOut_payload_0_7928 ? _zz_dataOut_payload_0_7905 : _zz_dataOut_payload_0_7917);
  assign _zz_dataOut_payload_0_7930 = (_zz_dataOut_payload_0_7928 ? _zz_dataOut_payload_0_7917 : _zz_dataOut_payload_0_7905);
  assign _zz_dataOut_payload_0_7931 = (_zz_dataOut_payload_0_7908 < _zz_dataOut_payload_0_7920);
  assign _zz_dataOut_payload_0_7932 = (_zz_dataOut_payload_0_7931 ? _zz_dataOut_payload_0_7908 : _zz_dataOut_payload_0_7920);
  assign _zz_dataOut_payload_0_7933 = (_zz_dataOut_payload_0_7931 ? _zz_dataOut_payload_0_7920 : _zz_dataOut_payload_0_7908);
  assign _zz_dataOut_payload_0_7934 = (_zz_dataOut_payload_0_7911 < _zz_dataOut_payload_0_7923);
  assign _zz_dataOut_payload_0_7935 = (_zz_dataOut_payload_0_7934 ? _zz_dataOut_payload_0_7911 : _zz_dataOut_payload_0_7923);
  assign _zz_dataOut_payload_0_7936 = (_zz_dataOut_payload_0_7934 ? _zz_dataOut_payload_0_7923 : _zz_dataOut_payload_0_7911);
  assign _zz_dataOut_payload_0_7937 = (_zz_dataOut_payload_0_7914 < _zz_dataOut_payload_0_7926);
  assign _zz_dataOut_payload_0_7938 = (_zz_dataOut_payload_0_7937 ? _zz_dataOut_payload_0_7914 : _zz_dataOut_payload_0_7926);
  assign _zz_dataOut_payload_0_7939 = (_zz_dataOut_payload_0_7937 ? _zz_dataOut_payload_0_7926 : _zz_dataOut_payload_0_7914);
  assign _zz_dataOut_payload_0_7940 = (_zz_dataOut_payload_0_7929 < _zz_dataOut_payload_0_7935);
  assign _zz_dataOut_payload_0_7941 = (_zz_dataOut_payload_0_7940 ? _zz_dataOut_payload_0_7929 : _zz_dataOut_payload_0_7935);
  assign _zz_dataOut_payload_0_7942 = (_zz_dataOut_payload_0_7940 ? _zz_dataOut_payload_0_7935 : _zz_dataOut_payload_0_7929);
  assign _zz_dataOut_payload_0_7943 = (_zz_dataOut_payload_0_7932 < _zz_dataOut_payload_0_7938);
  assign _zz_dataOut_payload_0_7944 = (_zz_dataOut_payload_0_7943 ? _zz_dataOut_payload_0_7932 : _zz_dataOut_payload_0_7938);
  assign _zz_dataOut_payload_0_7945 = (_zz_dataOut_payload_0_7943 ? _zz_dataOut_payload_0_7938 : _zz_dataOut_payload_0_7932);
  assign _zz_dataOut_payload_0_7946 = (_zz_dataOut_payload_0_7941 < _zz_dataOut_payload_0_7944);
  assign _zz_dataOut_payload_0_7947 = (_zz_dataOut_payload_0_7942 < _zz_dataOut_payload_0_7945);
  assign _zz_dataOut_payload_0_7952 = (_zz_dataOut_payload_0_7930 < _zz_dataOut_payload_0_7936);
  assign _zz_dataOut_payload_0_7953 = (_zz_dataOut_payload_0_7952 ? _zz_dataOut_payload_0_7930 : _zz_dataOut_payload_0_7936);
  assign _zz_dataOut_payload_0_7954 = (_zz_dataOut_payload_0_7952 ? _zz_dataOut_payload_0_7936 : _zz_dataOut_payload_0_7930);
  assign _zz_dataOut_payload_0_7955 = (_zz_dataOut_payload_0_7933 < _zz_dataOut_payload_0_7939);
  assign _zz_dataOut_payload_0_7956 = (_zz_dataOut_payload_0_7955 ? _zz_dataOut_payload_0_7933 : _zz_dataOut_payload_0_7939);
  assign _zz_dataOut_payload_0_7957 = (_zz_dataOut_payload_0_7955 ? _zz_dataOut_payload_0_7939 : _zz_dataOut_payload_0_7933);
  assign _zz_dataOut_payload_0_7958 = (_zz_dataOut_payload_0_7953 < _zz_dataOut_payload_0_7956);
  assign _zz_dataOut_payload_0_7959 = (_zz_dataOut_payload_0_7954 < _zz_dataOut_payload_0_7957);
  assign _zz_dataOut_payload_0_7972 = (_zz_dataOut_payload_0_7906 < _zz_dataOut_payload_0_7918);
  assign _zz_dataOut_payload_0_7973 = (_zz_dataOut_payload_0_7972 ? _zz_dataOut_payload_0_7906 : _zz_dataOut_payload_0_7918);
  assign _zz_dataOut_payload_0_7974 = (_zz_dataOut_payload_0_7972 ? _zz_dataOut_payload_0_7918 : _zz_dataOut_payload_0_7906);
  assign _zz_dataOut_payload_0_7975 = (_zz_dataOut_payload_0_7909 < _zz_dataOut_payload_0_7921);
  assign _zz_dataOut_payload_0_7976 = (_zz_dataOut_payload_0_7975 ? _zz_dataOut_payload_0_7909 : _zz_dataOut_payload_0_7921);
  assign _zz_dataOut_payload_0_7977 = (_zz_dataOut_payload_0_7975 ? _zz_dataOut_payload_0_7921 : _zz_dataOut_payload_0_7909);
  assign _zz_dataOut_payload_0_7978 = (_zz_dataOut_payload_0_7912 < _zz_dataOut_payload_0_7924);
  assign _zz_dataOut_payload_0_7979 = (_zz_dataOut_payload_0_7978 ? _zz_dataOut_payload_0_7912 : _zz_dataOut_payload_0_7924);
  assign _zz_dataOut_payload_0_7980 = (_zz_dataOut_payload_0_7978 ? _zz_dataOut_payload_0_7924 : _zz_dataOut_payload_0_7912);
  assign _zz_dataOut_payload_0_7981 = (_zz_dataOut_payload_0_7915 < _zz_dataOut_payload_0_7927);
  assign _zz_dataOut_payload_0_7982 = (_zz_dataOut_payload_0_7981 ? _zz_dataOut_payload_0_7915 : _zz_dataOut_payload_0_7927);
  assign _zz_dataOut_payload_0_7983 = (_zz_dataOut_payload_0_7981 ? _zz_dataOut_payload_0_7927 : _zz_dataOut_payload_0_7915);
  assign _zz_dataOut_payload_0_7984 = (_zz_dataOut_payload_0_7973 < _zz_dataOut_payload_0_7979);
  assign _zz_dataOut_payload_0_7985 = (_zz_dataOut_payload_0_7984 ? _zz_dataOut_payload_0_7973 : _zz_dataOut_payload_0_7979);
  assign _zz_dataOut_payload_0_7986 = (_zz_dataOut_payload_0_7984 ? _zz_dataOut_payload_0_7979 : _zz_dataOut_payload_0_7973);
  assign _zz_dataOut_payload_0_7987 = (_zz_dataOut_payload_0_7976 < _zz_dataOut_payload_0_7982);
  assign _zz_dataOut_payload_0_7988 = (_zz_dataOut_payload_0_7987 ? _zz_dataOut_payload_0_7976 : _zz_dataOut_payload_0_7982);
  assign _zz_dataOut_payload_0_7989 = (_zz_dataOut_payload_0_7987 ? _zz_dataOut_payload_0_7982 : _zz_dataOut_payload_0_7976);
  assign _zz_dataOut_payload_0_7990 = (_zz_dataOut_payload_0_7985 < _zz_dataOut_payload_0_7988);
  assign _zz_dataOut_payload_0_7991 = (_zz_dataOut_payload_0_7986 < _zz_dataOut_payload_0_7989);
  assign _zz_dataOut_payload_0_7996 = (_zz_dataOut_payload_0_7974 < _zz_dataOut_payload_0_7980);
  assign _zz_dataOut_payload_0_7997 = (_zz_dataOut_payload_0_7996 ? _zz_dataOut_payload_0_7974 : _zz_dataOut_payload_0_7980);
  assign _zz_dataOut_payload_0_7998 = (_zz_dataOut_payload_0_7996 ? _zz_dataOut_payload_0_7980 : _zz_dataOut_payload_0_7974);
  assign _zz_dataOut_payload_0_7999 = (_zz_dataOut_payload_0_7977 < _zz_dataOut_payload_0_7983);
  assign _zz_dataOut_payload_0_8000 = (_zz_dataOut_payload_0_7999 ? _zz_dataOut_payload_0_7977 : _zz_dataOut_payload_0_7983);
  assign _zz_dataOut_payload_0_8001 = (_zz_dataOut_payload_0_7999 ? _zz_dataOut_payload_0_7983 : _zz_dataOut_payload_0_7977);
  assign _zz_dataOut_payload_0_8002 = (_zz_dataOut_payload_0_7997 < _zz_dataOut_payload_0_8000);
  assign _zz_dataOut_payload_0_8003 = (_zz_dataOut_payload_0_7998 < _zz_dataOut_payload_0_8001);
  assign _zz_dataOut_payload_0_8320 = (_zz_dataOut_payload_0_8064 < _zz_dataOut_payload_0_8127);
  assign _zz_dataOut_payload_0_8321 = (_zz_dataOut_payload_0_8320 ? _zz_dataOut_payload_0_8064 : _zz_dataOut_payload_0_8127);
  assign _zz_dataOut_payload_0_8322 = (_zz_dataOut_payload_0_8320 ? _zz_dataOut_payload_0_8127 : _zz_dataOut_payload_0_8064);
  assign _zz_dataOut_payload_0_8323 = (_zz_dataOut_payload_0_8065 < _zz_dataOut_payload_0_8126);
  assign _zz_dataOut_payload_0_8324 = (_zz_dataOut_payload_0_8323 ? _zz_dataOut_payload_0_8065 : _zz_dataOut_payload_0_8126);
  assign _zz_dataOut_payload_0_8325 = (_zz_dataOut_payload_0_8323 ? _zz_dataOut_payload_0_8126 : _zz_dataOut_payload_0_8065);
  assign _zz_dataOut_payload_0_8326 = (_zz_dataOut_payload_0_8066 < _zz_dataOut_payload_0_8125);
  assign _zz_dataOut_payload_0_8327 = (_zz_dataOut_payload_0_8326 ? _zz_dataOut_payload_0_8066 : _zz_dataOut_payload_0_8125);
  assign _zz_dataOut_payload_0_8328 = (_zz_dataOut_payload_0_8326 ? _zz_dataOut_payload_0_8125 : _zz_dataOut_payload_0_8066);
  assign _zz_dataOut_payload_0_8329 = (_zz_dataOut_payload_0_8067 < _zz_dataOut_payload_0_8124);
  assign _zz_dataOut_payload_0_8330 = (_zz_dataOut_payload_0_8329 ? _zz_dataOut_payload_0_8067 : _zz_dataOut_payload_0_8124);
  assign _zz_dataOut_payload_0_8331 = (_zz_dataOut_payload_0_8329 ? _zz_dataOut_payload_0_8124 : _zz_dataOut_payload_0_8067);
  assign _zz_dataOut_payload_0_8332 = (_zz_dataOut_payload_0_8068 < _zz_dataOut_payload_0_8123);
  assign _zz_dataOut_payload_0_8333 = (_zz_dataOut_payload_0_8332 ? _zz_dataOut_payload_0_8068 : _zz_dataOut_payload_0_8123);
  assign _zz_dataOut_payload_0_8334 = (_zz_dataOut_payload_0_8332 ? _zz_dataOut_payload_0_8123 : _zz_dataOut_payload_0_8068);
  assign _zz_dataOut_payload_0_8335 = (_zz_dataOut_payload_0_8069 < _zz_dataOut_payload_0_8122);
  assign _zz_dataOut_payload_0_8336 = (_zz_dataOut_payload_0_8335 ? _zz_dataOut_payload_0_8069 : _zz_dataOut_payload_0_8122);
  assign _zz_dataOut_payload_0_8337 = (_zz_dataOut_payload_0_8335 ? _zz_dataOut_payload_0_8122 : _zz_dataOut_payload_0_8069);
  assign _zz_dataOut_payload_0_8338 = (_zz_dataOut_payload_0_8070 < _zz_dataOut_payload_0_8121);
  assign _zz_dataOut_payload_0_8339 = (_zz_dataOut_payload_0_8338 ? _zz_dataOut_payload_0_8070 : _zz_dataOut_payload_0_8121);
  assign _zz_dataOut_payload_0_8340 = (_zz_dataOut_payload_0_8338 ? _zz_dataOut_payload_0_8121 : _zz_dataOut_payload_0_8070);
  assign _zz_dataOut_payload_0_8341 = (_zz_dataOut_payload_0_8071 < _zz_dataOut_payload_0_8120);
  assign _zz_dataOut_payload_0_8342 = (_zz_dataOut_payload_0_8341 ? _zz_dataOut_payload_0_8071 : _zz_dataOut_payload_0_8120);
  assign _zz_dataOut_payload_0_8343 = (_zz_dataOut_payload_0_8341 ? _zz_dataOut_payload_0_8120 : _zz_dataOut_payload_0_8071);
  assign _zz_dataOut_payload_0_8344 = (_zz_dataOut_payload_0_8072 < _zz_dataOut_payload_0_8119);
  assign _zz_dataOut_payload_0_8345 = (_zz_dataOut_payload_0_8344 ? _zz_dataOut_payload_0_8072 : _zz_dataOut_payload_0_8119);
  assign _zz_dataOut_payload_0_8346 = (_zz_dataOut_payload_0_8344 ? _zz_dataOut_payload_0_8119 : _zz_dataOut_payload_0_8072);
  assign _zz_dataOut_payload_0_8347 = (_zz_dataOut_payload_0_8073 < _zz_dataOut_payload_0_8118);
  assign _zz_dataOut_payload_0_8348 = (_zz_dataOut_payload_0_8347 ? _zz_dataOut_payload_0_8073 : _zz_dataOut_payload_0_8118);
  assign _zz_dataOut_payload_0_8349 = (_zz_dataOut_payload_0_8347 ? _zz_dataOut_payload_0_8118 : _zz_dataOut_payload_0_8073);
  assign _zz_dataOut_payload_0_8350 = (_zz_dataOut_payload_0_8074 < _zz_dataOut_payload_0_8117);
  assign _zz_dataOut_payload_0_8351 = (_zz_dataOut_payload_0_8350 ? _zz_dataOut_payload_0_8074 : _zz_dataOut_payload_0_8117);
  assign _zz_dataOut_payload_0_8352 = (_zz_dataOut_payload_0_8350 ? _zz_dataOut_payload_0_8117 : _zz_dataOut_payload_0_8074);
  assign _zz_dataOut_payload_0_8353 = (_zz_dataOut_payload_0_8075 < _zz_dataOut_payload_0_8116);
  assign _zz_dataOut_payload_0_8354 = (_zz_dataOut_payload_0_8353 ? _zz_dataOut_payload_0_8075 : _zz_dataOut_payload_0_8116);
  assign _zz_dataOut_payload_0_8355 = (_zz_dataOut_payload_0_8353 ? _zz_dataOut_payload_0_8116 : _zz_dataOut_payload_0_8075);
  assign _zz_dataOut_payload_0_8356 = (_zz_dataOut_payload_0_8076 < _zz_dataOut_payload_0_8115);
  assign _zz_dataOut_payload_0_8357 = (_zz_dataOut_payload_0_8356 ? _zz_dataOut_payload_0_8076 : _zz_dataOut_payload_0_8115);
  assign _zz_dataOut_payload_0_8358 = (_zz_dataOut_payload_0_8356 ? _zz_dataOut_payload_0_8115 : _zz_dataOut_payload_0_8076);
  assign _zz_dataOut_payload_0_8359 = (_zz_dataOut_payload_0_8077 < _zz_dataOut_payload_0_8114);
  assign _zz_dataOut_payload_0_8360 = (_zz_dataOut_payload_0_8359 ? _zz_dataOut_payload_0_8077 : _zz_dataOut_payload_0_8114);
  assign _zz_dataOut_payload_0_8361 = (_zz_dataOut_payload_0_8359 ? _zz_dataOut_payload_0_8114 : _zz_dataOut_payload_0_8077);
  assign _zz_dataOut_payload_0_8362 = (_zz_dataOut_payload_0_8078 < _zz_dataOut_payload_0_8113);
  assign _zz_dataOut_payload_0_8363 = (_zz_dataOut_payload_0_8362 ? _zz_dataOut_payload_0_8078 : _zz_dataOut_payload_0_8113);
  assign _zz_dataOut_payload_0_8364 = (_zz_dataOut_payload_0_8362 ? _zz_dataOut_payload_0_8113 : _zz_dataOut_payload_0_8078);
  assign _zz_dataOut_payload_0_8365 = (_zz_dataOut_payload_0_8079 < _zz_dataOut_payload_0_8112);
  assign _zz_dataOut_payload_0_8366 = (_zz_dataOut_payload_0_8365 ? _zz_dataOut_payload_0_8079 : _zz_dataOut_payload_0_8112);
  assign _zz_dataOut_payload_0_8367 = (_zz_dataOut_payload_0_8365 ? _zz_dataOut_payload_0_8112 : _zz_dataOut_payload_0_8079);
  assign _zz_dataOut_payload_0_8368 = (_zz_dataOut_payload_0_8080 < _zz_dataOut_payload_0_8111);
  assign _zz_dataOut_payload_0_8369 = (_zz_dataOut_payload_0_8368 ? _zz_dataOut_payload_0_8080 : _zz_dataOut_payload_0_8111);
  assign _zz_dataOut_payload_0_8370 = (_zz_dataOut_payload_0_8368 ? _zz_dataOut_payload_0_8111 : _zz_dataOut_payload_0_8080);
  assign _zz_dataOut_payload_0_8371 = (_zz_dataOut_payload_0_8081 < _zz_dataOut_payload_0_8110);
  assign _zz_dataOut_payload_0_8372 = (_zz_dataOut_payload_0_8371 ? _zz_dataOut_payload_0_8081 : _zz_dataOut_payload_0_8110);
  assign _zz_dataOut_payload_0_8373 = (_zz_dataOut_payload_0_8371 ? _zz_dataOut_payload_0_8110 : _zz_dataOut_payload_0_8081);
  assign _zz_dataOut_payload_0_8374 = (_zz_dataOut_payload_0_8082 < _zz_dataOut_payload_0_8109);
  assign _zz_dataOut_payload_0_8375 = (_zz_dataOut_payload_0_8374 ? _zz_dataOut_payload_0_8082 : _zz_dataOut_payload_0_8109);
  assign _zz_dataOut_payload_0_8376 = (_zz_dataOut_payload_0_8374 ? _zz_dataOut_payload_0_8109 : _zz_dataOut_payload_0_8082);
  assign _zz_dataOut_payload_0_8377 = (_zz_dataOut_payload_0_8083 < _zz_dataOut_payload_0_8108);
  assign _zz_dataOut_payload_0_8378 = (_zz_dataOut_payload_0_8377 ? _zz_dataOut_payload_0_8083 : _zz_dataOut_payload_0_8108);
  assign _zz_dataOut_payload_0_8379 = (_zz_dataOut_payload_0_8377 ? _zz_dataOut_payload_0_8108 : _zz_dataOut_payload_0_8083);
  assign _zz_dataOut_payload_0_8380 = (_zz_dataOut_payload_0_8084 < _zz_dataOut_payload_0_8107);
  assign _zz_dataOut_payload_0_8381 = (_zz_dataOut_payload_0_8380 ? _zz_dataOut_payload_0_8084 : _zz_dataOut_payload_0_8107);
  assign _zz_dataOut_payload_0_8382 = (_zz_dataOut_payload_0_8380 ? _zz_dataOut_payload_0_8107 : _zz_dataOut_payload_0_8084);
  assign _zz_dataOut_payload_0_8383 = (_zz_dataOut_payload_0_8085 < _zz_dataOut_payload_0_8106);
  assign _zz_dataOut_payload_0_8384 = (_zz_dataOut_payload_0_8383 ? _zz_dataOut_payload_0_8085 : _zz_dataOut_payload_0_8106);
  assign _zz_dataOut_payload_0_8385 = (_zz_dataOut_payload_0_8383 ? _zz_dataOut_payload_0_8106 : _zz_dataOut_payload_0_8085);
  assign _zz_dataOut_payload_0_8386 = (_zz_dataOut_payload_0_8086 < _zz_dataOut_payload_0_8105);
  assign _zz_dataOut_payload_0_8387 = (_zz_dataOut_payload_0_8386 ? _zz_dataOut_payload_0_8086 : _zz_dataOut_payload_0_8105);
  assign _zz_dataOut_payload_0_8388 = (_zz_dataOut_payload_0_8386 ? _zz_dataOut_payload_0_8105 : _zz_dataOut_payload_0_8086);
  assign _zz_dataOut_payload_0_8389 = (_zz_dataOut_payload_0_8087 < _zz_dataOut_payload_0_8104);
  assign _zz_dataOut_payload_0_8390 = (_zz_dataOut_payload_0_8389 ? _zz_dataOut_payload_0_8087 : _zz_dataOut_payload_0_8104);
  assign _zz_dataOut_payload_0_8391 = (_zz_dataOut_payload_0_8389 ? _zz_dataOut_payload_0_8104 : _zz_dataOut_payload_0_8087);
  assign _zz_dataOut_payload_0_8392 = (_zz_dataOut_payload_0_8088 < _zz_dataOut_payload_0_8103);
  assign _zz_dataOut_payload_0_8393 = (_zz_dataOut_payload_0_8392 ? _zz_dataOut_payload_0_8088 : _zz_dataOut_payload_0_8103);
  assign _zz_dataOut_payload_0_8394 = (_zz_dataOut_payload_0_8392 ? _zz_dataOut_payload_0_8103 : _zz_dataOut_payload_0_8088);
  assign _zz_dataOut_payload_0_8395 = (_zz_dataOut_payload_0_8089 < _zz_dataOut_payload_0_8102);
  assign _zz_dataOut_payload_0_8396 = (_zz_dataOut_payload_0_8395 ? _zz_dataOut_payload_0_8089 : _zz_dataOut_payload_0_8102);
  assign _zz_dataOut_payload_0_8397 = (_zz_dataOut_payload_0_8395 ? _zz_dataOut_payload_0_8102 : _zz_dataOut_payload_0_8089);
  assign _zz_dataOut_payload_0_8398 = (_zz_dataOut_payload_0_8090 < _zz_dataOut_payload_0_8101);
  assign _zz_dataOut_payload_0_8399 = (_zz_dataOut_payload_0_8398 ? _zz_dataOut_payload_0_8090 : _zz_dataOut_payload_0_8101);
  assign _zz_dataOut_payload_0_8400 = (_zz_dataOut_payload_0_8398 ? _zz_dataOut_payload_0_8101 : _zz_dataOut_payload_0_8090);
  assign _zz_dataOut_payload_0_8401 = (_zz_dataOut_payload_0_8091 < _zz_dataOut_payload_0_8100);
  assign _zz_dataOut_payload_0_8402 = (_zz_dataOut_payload_0_8401 ? _zz_dataOut_payload_0_8091 : _zz_dataOut_payload_0_8100);
  assign _zz_dataOut_payload_0_8403 = (_zz_dataOut_payload_0_8401 ? _zz_dataOut_payload_0_8100 : _zz_dataOut_payload_0_8091);
  assign _zz_dataOut_payload_0_8404 = (_zz_dataOut_payload_0_8092 < _zz_dataOut_payload_0_8099);
  assign _zz_dataOut_payload_0_8405 = (_zz_dataOut_payload_0_8404 ? _zz_dataOut_payload_0_8092 : _zz_dataOut_payload_0_8099);
  assign _zz_dataOut_payload_0_8406 = (_zz_dataOut_payload_0_8404 ? _zz_dataOut_payload_0_8099 : _zz_dataOut_payload_0_8092);
  assign _zz_dataOut_payload_0_8407 = (_zz_dataOut_payload_0_8093 < _zz_dataOut_payload_0_8098);
  assign _zz_dataOut_payload_0_8408 = (_zz_dataOut_payload_0_8407 ? _zz_dataOut_payload_0_8093 : _zz_dataOut_payload_0_8098);
  assign _zz_dataOut_payload_0_8409 = (_zz_dataOut_payload_0_8407 ? _zz_dataOut_payload_0_8098 : _zz_dataOut_payload_0_8093);
  assign _zz_dataOut_payload_0_8410 = (_zz_dataOut_payload_0_8094 < _zz_dataOut_payload_0_8097);
  assign _zz_dataOut_payload_0_8411 = (_zz_dataOut_payload_0_8410 ? _zz_dataOut_payload_0_8094 : _zz_dataOut_payload_0_8097);
  assign _zz_dataOut_payload_0_8412 = (_zz_dataOut_payload_0_8410 ? _zz_dataOut_payload_0_8097 : _zz_dataOut_payload_0_8094);
  assign _zz_dataOut_payload_0_8413 = (_zz_dataOut_payload_0_8095 < _zz_dataOut_payload_0_8096);
  assign _zz_dataOut_payload_0_8414 = (_zz_dataOut_payload_0_8413 ? _zz_dataOut_payload_0_8095 : _zz_dataOut_payload_0_8096);
  assign _zz_dataOut_payload_0_8415 = (_zz_dataOut_payload_0_8413 ? _zz_dataOut_payload_0_8096 : _zz_dataOut_payload_0_8095);
  assign _zz_dataOut_payload_0_8416 = (_zz_dataOut_payload_0_8321 < _zz_dataOut_payload_0_8369);
  assign _zz_dataOut_payload_0_8417 = (_zz_dataOut_payload_0_8416 ? _zz_dataOut_payload_0_8321 : _zz_dataOut_payload_0_8369);
  assign _zz_dataOut_payload_0_8418 = (_zz_dataOut_payload_0_8416 ? _zz_dataOut_payload_0_8369 : _zz_dataOut_payload_0_8321);
  assign _zz_dataOut_payload_0_8419 = (_zz_dataOut_payload_0_8324 < _zz_dataOut_payload_0_8372);
  assign _zz_dataOut_payload_0_8420 = (_zz_dataOut_payload_0_8419 ? _zz_dataOut_payload_0_8324 : _zz_dataOut_payload_0_8372);
  assign _zz_dataOut_payload_0_8421 = (_zz_dataOut_payload_0_8419 ? _zz_dataOut_payload_0_8372 : _zz_dataOut_payload_0_8324);
  assign _zz_dataOut_payload_0_8422 = (_zz_dataOut_payload_0_8327 < _zz_dataOut_payload_0_8375);
  assign _zz_dataOut_payload_0_8423 = (_zz_dataOut_payload_0_8422 ? _zz_dataOut_payload_0_8327 : _zz_dataOut_payload_0_8375);
  assign _zz_dataOut_payload_0_8424 = (_zz_dataOut_payload_0_8422 ? _zz_dataOut_payload_0_8375 : _zz_dataOut_payload_0_8327);
  assign _zz_dataOut_payload_0_8425 = (_zz_dataOut_payload_0_8330 < _zz_dataOut_payload_0_8378);
  assign _zz_dataOut_payload_0_8426 = (_zz_dataOut_payload_0_8425 ? _zz_dataOut_payload_0_8330 : _zz_dataOut_payload_0_8378);
  assign _zz_dataOut_payload_0_8427 = (_zz_dataOut_payload_0_8425 ? _zz_dataOut_payload_0_8378 : _zz_dataOut_payload_0_8330);
  assign _zz_dataOut_payload_0_8428 = (_zz_dataOut_payload_0_8333 < _zz_dataOut_payload_0_8381);
  assign _zz_dataOut_payload_0_8429 = (_zz_dataOut_payload_0_8428 ? _zz_dataOut_payload_0_8333 : _zz_dataOut_payload_0_8381);
  assign _zz_dataOut_payload_0_8430 = (_zz_dataOut_payload_0_8428 ? _zz_dataOut_payload_0_8381 : _zz_dataOut_payload_0_8333);
  assign _zz_dataOut_payload_0_8431 = (_zz_dataOut_payload_0_8336 < _zz_dataOut_payload_0_8384);
  assign _zz_dataOut_payload_0_8432 = (_zz_dataOut_payload_0_8431 ? _zz_dataOut_payload_0_8336 : _zz_dataOut_payload_0_8384);
  assign _zz_dataOut_payload_0_8433 = (_zz_dataOut_payload_0_8431 ? _zz_dataOut_payload_0_8384 : _zz_dataOut_payload_0_8336);
  assign _zz_dataOut_payload_0_8434 = (_zz_dataOut_payload_0_8339 < _zz_dataOut_payload_0_8387);
  assign _zz_dataOut_payload_0_8435 = (_zz_dataOut_payload_0_8434 ? _zz_dataOut_payload_0_8339 : _zz_dataOut_payload_0_8387);
  assign _zz_dataOut_payload_0_8436 = (_zz_dataOut_payload_0_8434 ? _zz_dataOut_payload_0_8387 : _zz_dataOut_payload_0_8339);
  assign _zz_dataOut_payload_0_8437 = (_zz_dataOut_payload_0_8342 < _zz_dataOut_payload_0_8390);
  assign _zz_dataOut_payload_0_8438 = (_zz_dataOut_payload_0_8437 ? _zz_dataOut_payload_0_8342 : _zz_dataOut_payload_0_8390);
  assign _zz_dataOut_payload_0_8439 = (_zz_dataOut_payload_0_8437 ? _zz_dataOut_payload_0_8390 : _zz_dataOut_payload_0_8342);
  assign _zz_dataOut_payload_0_8440 = (_zz_dataOut_payload_0_8345 < _zz_dataOut_payload_0_8393);
  assign _zz_dataOut_payload_0_8441 = (_zz_dataOut_payload_0_8440 ? _zz_dataOut_payload_0_8345 : _zz_dataOut_payload_0_8393);
  assign _zz_dataOut_payload_0_8442 = (_zz_dataOut_payload_0_8440 ? _zz_dataOut_payload_0_8393 : _zz_dataOut_payload_0_8345);
  assign _zz_dataOut_payload_0_8443 = (_zz_dataOut_payload_0_8348 < _zz_dataOut_payload_0_8396);
  assign _zz_dataOut_payload_0_8444 = (_zz_dataOut_payload_0_8443 ? _zz_dataOut_payload_0_8348 : _zz_dataOut_payload_0_8396);
  assign _zz_dataOut_payload_0_8445 = (_zz_dataOut_payload_0_8443 ? _zz_dataOut_payload_0_8396 : _zz_dataOut_payload_0_8348);
  assign _zz_dataOut_payload_0_8446 = (_zz_dataOut_payload_0_8351 < _zz_dataOut_payload_0_8399);
  assign _zz_dataOut_payload_0_8447 = (_zz_dataOut_payload_0_8446 ? _zz_dataOut_payload_0_8351 : _zz_dataOut_payload_0_8399);
  assign _zz_dataOut_payload_0_8448 = (_zz_dataOut_payload_0_8446 ? _zz_dataOut_payload_0_8399 : _zz_dataOut_payload_0_8351);
  assign _zz_dataOut_payload_0_8449 = (_zz_dataOut_payload_0_8354 < _zz_dataOut_payload_0_8402);
  assign _zz_dataOut_payload_0_8450 = (_zz_dataOut_payload_0_8449 ? _zz_dataOut_payload_0_8354 : _zz_dataOut_payload_0_8402);
  assign _zz_dataOut_payload_0_8451 = (_zz_dataOut_payload_0_8449 ? _zz_dataOut_payload_0_8402 : _zz_dataOut_payload_0_8354);
  assign _zz_dataOut_payload_0_8452 = (_zz_dataOut_payload_0_8357 < _zz_dataOut_payload_0_8405);
  assign _zz_dataOut_payload_0_8453 = (_zz_dataOut_payload_0_8452 ? _zz_dataOut_payload_0_8357 : _zz_dataOut_payload_0_8405);
  assign _zz_dataOut_payload_0_8454 = (_zz_dataOut_payload_0_8452 ? _zz_dataOut_payload_0_8405 : _zz_dataOut_payload_0_8357);
  assign _zz_dataOut_payload_0_8455 = (_zz_dataOut_payload_0_8360 < _zz_dataOut_payload_0_8408);
  assign _zz_dataOut_payload_0_8456 = (_zz_dataOut_payload_0_8455 ? _zz_dataOut_payload_0_8360 : _zz_dataOut_payload_0_8408);
  assign _zz_dataOut_payload_0_8457 = (_zz_dataOut_payload_0_8455 ? _zz_dataOut_payload_0_8408 : _zz_dataOut_payload_0_8360);
  assign _zz_dataOut_payload_0_8458 = (_zz_dataOut_payload_0_8363 < _zz_dataOut_payload_0_8411);
  assign _zz_dataOut_payload_0_8459 = (_zz_dataOut_payload_0_8458 ? _zz_dataOut_payload_0_8363 : _zz_dataOut_payload_0_8411);
  assign _zz_dataOut_payload_0_8460 = (_zz_dataOut_payload_0_8458 ? _zz_dataOut_payload_0_8411 : _zz_dataOut_payload_0_8363);
  assign _zz_dataOut_payload_0_8461 = (_zz_dataOut_payload_0_8366 < _zz_dataOut_payload_0_8414);
  assign _zz_dataOut_payload_0_8462 = (_zz_dataOut_payload_0_8461 ? _zz_dataOut_payload_0_8366 : _zz_dataOut_payload_0_8414);
  assign _zz_dataOut_payload_0_8463 = (_zz_dataOut_payload_0_8461 ? _zz_dataOut_payload_0_8414 : _zz_dataOut_payload_0_8366);
  assign _zz_dataOut_payload_0_8464 = (_zz_dataOut_payload_0_8417 < _zz_dataOut_payload_0_8441);
  assign _zz_dataOut_payload_0_8465 = (_zz_dataOut_payload_0_8464 ? _zz_dataOut_payload_0_8417 : _zz_dataOut_payload_0_8441);
  assign _zz_dataOut_payload_0_8466 = (_zz_dataOut_payload_0_8464 ? _zz_dataOut_payload_0_8441 : _zz_dataOut_payload_0_8417);
  assign _zz_dataOut_payload_0_8467 = (_zz_dataOut_payload_0_8420 < _zz_dataOut_payload_0_8444);
  assign _zz_dataOut_payload_0_8468 = (_zz_dataOut_payload_0_8467 ? _zz_dataOut_payload_0_8420 : _zz_dataOut_payload_0_8444);
  assign _zz_dataOut_payload_0_8469 = (_zz_dataOut_payload_0_8467 ? _zz_dataOut_payload_0_8444 : _zz_dataOut_payload_0_8420);
  assign _zz_dataOut_payload_0_8470 = (_zz_dataOut_payload_0_8423 < _zz_dataOut_payload_0_8447);
  assign _zz_dataOut_payload_0_8471 = (_zz_dataOut_payload_0_8470 ? _zz_dataOut_payload_0_8423 : _zz_dataOut_payload_0_8447);
  assign _zz_dataOut_payload_0_8472 = (_zz_dataOut_payload_0_8470 ? _zz_dataOut_payload_0_8447 : _zz_dataOut_payload_0_8423);
  assign _zz_dataOut_payload_0_8473 = (_zz_dataOut_payload_0_8426 < _zz_dataOut_payload_0_8450);
  assign _zz_dataOut_payload_0_8474 = (_zz_dataOut_payload_0_8473 ? _zz_dataOut_payload_0_8426 : _zz_dataOut_payload_0_8450);
  assign _zz_dataOut_payload_0_8475 = (_zz_dataOut_payload_0_8473 ? _zz_dataOut_payload_0_8450 : _zz_dataOut_payload_0_8426);
  assign _zz_dataOut_payload_0_8476 = (_zz_dataOut_payload_0_8429 < _zz_dataOut_payload_0_8453);
  assign _zz_dataOut_payload_0_8477 = (_zz_dataOut_payload_0_8476 ? _zz_dataOut_payload_0_8429 : _zz_dataOut_payload_0_8453);
  assign _zz_dataOut_payload_0_8478 = (_zz_dataOut_payload_0_8476 ? _zz_dataOut_payload_0_8453 : _zz_dataOut_payload_0_8429);
  assign _zz_dataOut_payload_0_8479 = (_zz_dataOut_payload_0_8432 < _zz_dataOut_payload_0_8456);
  assign _zz_dataOut_payload_0_8480 = (_zz_dataOut_payload_0_8479 ? _zz_dataOut_payload_0_8432 : _zz_dataOut_payload_0_8456);
  assign _zz_dataOut_payload_0_8481 = (_zz_dataOut_payload_0_8479 ? _zz_dataOut_payload_0_8456 : _zz_dataOut_payload_0_8432);
  assign _zz_dataOut_payload_0_8482 = (_zz_dataOut_payload_0_8435 < _zz_dataOut_payload_0_8459);
  assign _zz_dataOut_payload_0_8483 = (_zz_dataOut_payload_0_8482 ? _zz_dataOut_payload_0_8435 : _zz_dataOut_payload_0_8459);
  assign _zz_dataOut_payload_0_8484 = (_zz_dataOut_payload_0_8482 ? _zz_dataOut_payload_0_8459 : _zz_dataOut_payload_0_8435);
  assign _zz_dataOut_payload_0_8485 = (_zz_dataOut_payload_0_8438 < _zz_dataOut_payload_0_8462);
  assign _zz_dataOut_payload_0_8486 = (_zz_dataOut_payload_0_8485 ? _zz_dataOut_payload_0_8438 : _zz_dataOut_payload_0_8462);
  assign _zz_dataOut_payload_0_8487 = (_zz_dataOut_payload_0_8485 ? _zz_dataOut_payload_0_8462 : _zz_dataOut_payload_0_8438);
  assign _zz_dataOut_payload_0_8488 = (_zz_dataOut_payload_0_8465 < _zz_dataOut_payload_0_8477);
  assign _zz_dataOut_payload_0_8489 = (_zz_dataOut_payload_0_8488 ? _zz_dataOut_payload_0_8465 : _zz_dataOut_payload_0_8477);
  assign _zz_dataOut_payload_0_8490 = (_zz_dataOut_payload_0_8488 ? _zz_dataOut_payload_0_8477 : _zz_dataOut_payload_0_8465);
  assign _zz_dataOut_payload_0_8491 = (_zz_dataOut_payload_0_8468 < _zz_dataOut_payload_0_8480);
  assign _zz_dataOut_payload_0_8492 = (_zz_dataOut_payload_0_8491 ? _zz_dataOut_payload_0_8468 : _zz_dataOut_payload_0_8480);
  assign _zz_dataOut_payload_0_8493 = (_zz_dataOut_payload_0_8491 ? _zz_dataOut_payload_0_8480 : _zz_dataOut_payload_0_8468);
  assign _zz_dataOut_payload_0_8494 = (_zz_dataOut_payload_0_8471 < _zz_dataOut_payload_0_8483);
  assign _zz_dataOut_payload_0_8495 = (_zz_dataOut_payload_0_8494 ? _zz_dataOut_payload_0_8471 : _zz_dataOut_payload_0_8483);
  assign _zz_dataOut_payload_0_8496 = (_zz_dataOut_payload_0_8494 ? _zz_dataOut_payload_0_8483 : _zz_dataOut_payload_0_8471);
  assign _zz_dataOut_payload_0_8497 = (_zz_dataOut_payload_0_8474 < _zz_dataOut_payload_0_8486);
  assign _zz_dataOut_payload_0_8498 = (_zz_dataOut_payload_0_8497 ? _zz_dataOut_payload_0_8474 : _zz_dataOut_payload_0_8486);
  assign _zz_dataOut_payload_0_8499 = (_zz_dataOut_payload_0_8497 ? _zz_dataOut_payload_0_8486 : _zz_dataOut_payload_0_8474);
  assign _zz_dataOut_payload_0_8500 = (_zz_dataOut_payload_0_8489 < _zz_dataOut_payload_0_8495);
  assign _zz_dataOut_payload_0_8501 = (_zz_dataOut_payload_0_8500 ? _zz_dataOut_payload_0_8489 : _zz_dataOut_payload_0_8495);
  assign _zz_dataOut_payload_0_8502 = (_zz_dataOut_payload_0_8500 ? _zz_dataOut_payload_0_8495 : _zz_dataOut_payload_0_8489);
  assign _zz_dataOut_payload_0_8503 = (_zz_dataOut_payload_0_8492 < _zz_dataOut_payload_0_8498);
  assign _zz_dataOut_payload_0_8504 = (_zz_dataOut_payload_0_8503 ? _zz_dataOut_payload_0_8492 : _zz_dataOut_payload_0_8498);
  assign _zz_dataOut_payload_0_8505 = (_zz_dataOut_payload_0_8503 ? _zz_dataOut_payload_0_8498 : _zz_dataOut_payload_0_8492);
  assign _zz_dataOut_payload_0_8506 = (_zz_dataOut_payload_0_8501 < _zz_dataOut_payload_0_8504);
  assign _zz_dataOut_payload_0_8507 = (_zz_dataOut_payload_0_8502 < _zz_dataOut_payload_0_8505);
  assign _zz_dataOut_payload_0_8512 = (_zz_dataOut_payload_0_8490 < _zz_dataOut_payload_0_8496);
  assign _zz_dataOut_payload_0_8513 = (_zz_dataOut_payload_0_8512 ? _zz_dataOut_payload_0_8490 : _zz_dataOut_payload_0_8496);
  assign _zz_dataOut_payload_0_8514 = (_zz_dataOut_payload_0_8512 ? _zz_dataOut_payload_0_8496 : _zz_dataOut_payload_0_8490);
  assign _zz_dataOut_payload_0_8515 = (_zz_dataOut_payload_0_8493 < _zz_dataOut_payload_0_8499);
  assign _zz_dataOut_payload_0_8516 = (_zz_dataOut_payload_0_8515 ? _zz_dataOut_payload_0_8493 : _zz_dataOut_payload_0_8499);
  assign _zz_dataOut_payload_0_8517 = (_zz_dataOut_payload_0_8515 ? _zz_dataOut_payload_0_8499 : _zz_dataOut_payload_0_8493);
  assign _zz_dataOut_payload_0_8518 = (_zz_dataOut_payload_0_8513 < _zz_dataOut_payload_0_8516);
  assign _zz_dataOut_payload_0_8519 = (_zz_dataOut_payload_0_8514 < _zz_dataOut_payload_0_8517);
  assign _zz_dataOut_payload_0_8532 = (_zz_dataOut_payload_0_8466 < _zz_dataOut_payload_0_8478);
  assign _zz_dataOut_payload_0_8533 = (_zz_dataOut_payload_0_8532 ? _zz_dataOut_payload_0_8466 : _zz_dataOut_payload_0_8478);
  assign _zz_dataOut_payload_0_8534 = (_zz_dataOut_payload_0_8532 ? _zz_dataOut_payload_0_8478 : _zz_dataOut_payload_0_8466);
  assign _zz_dataOut_payload_0_8535 = (_zz_dataOut_payload_0_8469 < _zz_dataOut_payload_0_8481);
  assign _zz_dataOut_payload_0_8536 = (_zz_dataOut_payload_0_8535 ? _zz_dataOut_payload_0_8469 : _zz_dataOut_payload_0_8481);
  assign _zz_dataOut_payload_0_8537 = (_zz_dataOut_payload_0_8535 ? _zz_dataOut_payload_0_8481 : _zz_dataOut_payload_0_8469);
  assign _zz_dataOut_payload_0_8538 = (_zz_dataOut_payload_0_8472 < _zz_dataOut_payload_0_8484);
  assign _zz_dataOut_payload_0_8539 = (_zz_dataOut_payload_0_8538 ? _zz_dataOut_payload_0_8472 : _zz_dataOut_payload_0_8484);
  assign _zz_dataOut_payload_0_8540 = (_zz_dataOut_payload_0_8538 ? _zz_dataOut_payload_0_8484 : _zz_dataOut_payload_0_8472);
  assign _zz_dataOut_payload_0_8541 = (_zz_dataOut_payload_0_8475 < _zz_dataOut_payload_0_8487);
  assign _zz_dataOut_payload_0_8542 = (_zz_dataOut_payload_0_8541 ? _zz_dataOut_payload_0_8475 : _zz_dataOut_payload_0_8487);
  assign _zz_dataOut_payload_0_8543 = (_zz_dataOut_payload_0_8541 ? _zz_dataOut_payload_0_8487 : _zz_dataOut_payload_0_8475);
  assign _zz_dataOut_payload_0_8544 = (_zz_dataOut_payload_0_8533 < _zz_dataOut_payload_0_8539);
  assign _zz_dataOut_payload_0_8545 = (_zz_dataOut_payload_0_8544 ? _zz_dataOut_payload_0_8533 : _zz_dataOut_payload_0_8539);
  assign _zz_dataOut_payload_0_8546 = (_zz_dataOut_payload_0_8544 ? _zz_dataOut_payload_0_8539 : _zz_dataOut_payload_0_8533);
  assign _zz_dataOut_payload_0_8547 = (_zz_dataOut_payload_0_8536 < _zz_dataOut_payload_0_8542);
  assign _zz_dataOut_payload_0_8548 = (_zz_dataOut_payload_0_8547 ? _zz_dataOut_payload_0_8536 : _zz_dataOut_payload_0_8542);
  assign _zz_dataOut_payload_0_8549 = (_zz_dataOut_payload_0_8547 ? _zz_dataOut_payload_0_8542 : _zz_dataOut_payload_0_8536);
  assign _zz_dataOut_payload_0_8550 = (_zz_dataOut_payload_0_8545 < _zz_dataOut_payload_0_8548);
  assign _zz_dataOut_payload_0_8551 = (_zz_dataOut_payload_0_8546 < _zz_dataOut_payload_0_8549);
  assign _zz_dataOut_payload_0_8556 = (_zz_dataOut_payload_0_8534 < _zz_dataOut_payload_0_8540);
  assign _zz_dataOut_payload_0_8557 = (_zz_dataOut_payload_0_8556 ? _zz_dataOut_payload_0_8534 : _zz_dataOut_payload_0_8540);
  assign _zz_dataOut_payload_0_8558 = (_zz_dataOut_payload_0_8556 ? _zz_dataOut_payload_0_8540 : _zz_dataOut_payload_0_8534);
  assign _zz_dataOut_payload_0_8559 = (_zz_dataOut_payload_0_8537 < _zz_dataOut_payload_0_8543);
  assign _zz_dataOut_payload_0_8560 = (_zz_dataOut_payload_0_8559 ? _zz_dataOut_payload_0_8537 : _zz_dataOut_payload_0_8543);
  assign _zz_dataOut_payload_0_8561 = (_zz_dataOut_payload_0_8559 ? _zz_dataOut_payload_0_8543 : _zz_dataOut_payload_0_8537);
  assign _zz_dataOut_payload_0_8562 = (_zz_dataOut_payload_0_8557 < _zz_dataOut_payload_0_8560);
  assign _zz_dataOut_payload_0_8563 = (_zz_dataOut_payload_0_8558 < _zz_dataOut_payload_0_8561);
  assign _zz_dataOut_payload_0_8592 = (_zz_dataOut_payload_0_8418 < _zz_dataOut_payload_0_8442);
  assign _zz_dataOut_payload_0_8593 = (_zz_dataOut_payload_0_8592 ? _zz_dataOut_payload_0_8418 : _zz_dataOut_payload_0_8442);
  assign _zz_dataOut_payload_0_8594 = (_zz_dataOut_payload_0_8592 ? _zz_dataOut_payload_0_8442 : _zz_dataOut_payload_0_8418);
  assign _zz_dataOut_payload_0_8595 = (_zz_dataOut_payload_0_8421 < _zz_dataOut_payload_0_8445);
  assign _zz_dataOut_payload_0_8596 = (_zz_dataOut_payload_0_8595 ? _zz_dataOut_payload_0_8421 : _zz_dataOut_payload_0_8445);
  assign _zz_dataOut_payload_0_8597 = (_zz_dataOut_payload_0_8595 ? _zz_dataOut_payload_0_8445 : _zz_dataOut_payload_0_8421);
  assign _zz_dataOut_payload_0_8598 = (_zz_dataOut_payload_0_8424 < _zz_dataOut_payload_0_8448);
  assign _zz_dataOut_payload_0_8599 = (_zz_dataOut_payload_0_8598 ? _zz_dataOut_payload_0_8424 : _zz_dataOut_payload_0_8448);
  assign _zz_dataOut_payload_0_8600 = (_zz_dataOut_payload_0_8598 ? _zz_dataOut_payload_0_8448 : _zz_dataOut_payload_0_8424);
  assign _zz_dataOut_payload_0_8601 = (_zz_dataOut_payload_0_8427 < _zz_dataOut_payload_0_8451);
  assign _zz_dataOut_payload_0_8602 = (_zz_dataOut_payload_0_8601 ? _zz_dataOut_payload_0_8427 : _zz_dataOut_payload_0_8451);
  assign _zz_dataOut_payload_0_8603 = (_zz_dataOut_payload_0_8601 ? _zz_dataOut_payload_0_8451 : _zz_dataOut_payload_0_8427);
  assign _zz_dataOut_payload_0_8604 = (_zz_dataOut_payload_0_8430 < _zz_dataOut_payload_0_8454);
  assign _zz_dataOut_payload_0_8605 = (_zz_dataOut_payload_0_8604 ? _zz_dataOut_payload_0_8430 : _zz_dataOut_payload_0_8454);
  assign _zz_dataOut_payload_0_8606 = (_zz_dataOut_payload_0_8604 ? _zz_dataOut_payload_0_8454 : _zz_dataOut_payload_0_8430);
  assign _zz_dataOut_payload_0_8607 = (_zz_dataOut_payload_0_8433 < _zz_dataOut_payload_0_8457);
  assign _zz_dataOut_payload_0_8608 = (_zz_dataOut_payload_0_8607 ? _zz_dataOut_payload_0_8433 : _zz_dataOut_payload_0_8457);
  assign _zz_dataOut_payload_0_8609 = (_zz_dataOut_payload_0_8607 ? _zz_dataOut_payload_0_8457 : _zz_dataOut_payload_0_8433);
  assign _zz_dataOut_payload_0_8610 = (_zz_dataOut_payload_0_8436 < _zz_dataOut_payload_0_8460);
  assign _zz_dataOut_payload_0_8611 = (_zz_dataOut_payload_0_8610 ? _zz_dataOut_payload_0_8436 : _zz_dataOut_payload_0_8460);
  assign _zz_dataOut_payload_0_8612 = (_zz_dataOut_payload_0_8610 ? _zz_dataOut_payload_0_8460 : _zz_dataOut_payload_0_8436);
  assign _zz_dataOut_payload_0_8613 = (_zz_dataOut_payload_0_8439 < _zz_dataOut_payload_0_8463);
  assign _zz_dataOut_payload_0_8614 = (_zz_dataOut_payload_0_8613 ? _zz_dataOut_payload_0_8439 : _zz_dataOut_payload_0_8463);
  assign _zz_dataOut_payload_0_8615 = (_zz_dataOut_payload_0_8613 ? _zz_dataOut_payload_0_8463 : _zz_dataOut_payload_0_8439);
  assign _zz_dataOut_payload_0_8616 = (_zz_dataOut_payload_0_8593 < _zz_dataOut_payload_0_8605);
  assign _zz_dataOut_payload_0_8617 = (_zz_dataOut_payload_0_8616 ? _zz_dataOut_payload_0_8593 : _zz_dataOut_payload_0_8605);
  assign _zz_dataOut_payload_0_8618 = (_zz_dataOut_payload_0_8616 ? _zz_dataOut_payload_0_8605 : _zz_dataOut_payload_0_8593);
  assign _zz_dataOut_payload_0_8619 = (_zz_dataOut_payload_0_8596 < _zz_dataOut_payload_0_8608);
  assign _zz_dataOut_payload_0_8620 = (_zz_dataOut_payload_0_8619 ? _zz_dataOut_payload_0_8596 : _zz_dataOut_payload_0_8608);
  assign _zz_dataOut_payload_0_8621 = (_zz_dataOut_payload_0_8619 ? _zz_dataOut_payload_0_8608 : _zz_dataOut_payload_0_8596);
  assign _zz_dataOut_payload_0_8622 = (_zz_dataOut_payload_0_8599 < _zz_dataOut_payload_0_8611);
  assign _zz_dataOut_payload_0_8623 = (_zz_dataOut_payload_0_8622 ? _zz_dataOut_payload_0_8599 : _zz_dataOut_payload_0_8611);
  assign _zz_dataOut_payload_0_8624 = (_zz_dataOut_payload_0_8622 ? _zz_dataOut_payload_0_8611 : _zz_dataOut_payload_0_8599);
  assign _zz_dataOut_payload_0_8625 = (_zz_dataOut_payload_0_8602 < _zz_dataOut_payload_0_8614);
  assign _zz_dataOut_payload_0_8626 = (_zz_dataOut_payload_0_8625 ? _zz_dataOut_payload_0_8602 : _zz_dataOut_payload_0_8614);
  assign _zz_dataOut_payload_0_8627 = (_zz_dataOut_payload_0_8625 ? _zz_dataOut_payload_0_8614 : _zz_dataOut_payload_0_8602);
  assign _zz_dataOut_payload_0_8628 = (_zz_dataOut_payload_0_8617 < _zz_dataOut_payload_0_8623);
  assign _zz_dataOut_payload_0_8629 = (_zz_dataOut_payload_0_8628 ? _zz_dataOut_payload_0_8617 : _zz_dataOut_payload_0_8623);
  assign _zz_dataOut_payload_0_8630 = (_zz_dataOut_payload_0_8628 ? _zz_dataOut_payload_0_8623 : _zz_dataOut_payload_0_8617);
  assign _zz_dataOut_payload_0_8631 = (_zz_dataOut_payload_0_8620 < _zz_dataOut_payload_0_8626);
  assign _zz_dataOut_payload_0_8632 = (_zz_dataOut_payload_0_8631 ? _zz_dataOut_payload_0_8620 : _zz_dataOut_payload_0_8626);
  assign _zz_dataOut_payload_0_8633 = (_zz_dataOut_payload_0_8631 ? _zz_dataOut_payload_0_8626 : _zz_dataOut_payload_0_8620);
  assign _zz_dataOut_payload_0_8634 = (_zz_dataOut_payload_0_8629 < _zz_dataOut_payload_0_8632);
  assign _zz_dataOut_payload_0_8635 = (_zz_dataOut_payload_0_8630 < _zz_dataOut_payload_0_8633);
  assign _zz_dataOut_payload_0_8640 = (_zz_dataOut_payload_0_8618 < _zz_dataOut_payload_0_8624);
  assign _zz_dataOut_payload_0_8641 = (_zz_dataOut_payload_0_8640 ? _zz_dataOut_payload_0_8618 : _zz_dataOut_payload_0_8624);
  assign _zz_dataOut_payload_0_8642 = (_zz_dataOut_payload_0_8640 ? _zz_dataOut_payload_0_8624 : _zz_dataOut_payload_0_8618);
  assign _zz_dataOut_payload_0_8643 = (_zz_dataOut_payload_0_8621 < _zz_dataOut_payload_0_8627);
  assign _zz_dataOut_payload_0_8644 = (_zz_dataOut_payload_0_8643 ? _zz_dataOut_payload_0_8621 : _zz_dataOut_payload_0_8627);
  assign _zz_dataOut_payload_0_8645 = (_zz_dataOut_payload_0_8643 ? _zz_dataOut_payload_0_8627 : _zz_dataOut_payload_0_8621);
  assign _zz_dataOut_payload_0_8646 = (_zz_dataOut_payload_0_8641 < _zz_dataOut_payload_0_8644);
  assign _zz_dataOut_payload_0_8647 = (_zz_dataOut_payload_0_8642 < _zz_dataOut_payload_0_8645);
  assign _zz_dataOut_payload_0_8660 = (_zz_dataOut_payload_0_8594 < _zz_dataOut_payload_0_8606);
  assign _zz_dataOut_payload_0_8661 = (_zz_dataOut_payload_0_8660 ? _zz_dataOut_payload_0_8594 : _zz_dataOut_payload_0_8606);
  assign _zz_dataOut_payload_0_8662 = (_zz_dataOut_payload_0_8660 ? _zz_dataOut_payload_0_8606 : _zz_dataOut_payload_0_8594);
  assign _zz_dataOut_payload_0_8663 = (_zz_dataOut_payload_0_8597 < _zz_dataOut_payload_0_8609);
  assign _zz_dataOut_payload_0_8664 = (_zz_dataOut_payload_0_8663 ? _zz_dataOut_payload_0_8597 : _zz_dataOut_payload_0_8609);
  assign _zz_dataOut_payload_0_8665 = (_zz_dataOut_payload_0_8663 ? _zz_dataOut_payload_0_8609 : _zz_dataOut_payload_0_8597);
  assign _zz_dataOut_payload_0_8666 = (_zz_dataOut_payload_0_8600 < _zz_dataOut_payload_0_8612);
  assign _zz_dataOut_payload_0_8667 = (_zz_dataOut_payload_0_8666 ? _zz_dataOut_payload_0_8600 : _zz_dataOut_payload_0_8612);
  assign _zz_dataOut_payload_0_8668 = (_zz_dataOut_payload_0_8666 ? _zz_dataOut_payload_0_8612 : _zz_dataOut_payload_0_8600);
  assign _zz_dataOut_payload_0_8669 = (_zz_dataOut_payload_0_8603 < _zz_dataOut_payload_0_8615);
  assign _zz_dataOut_payload_0_8670 = (_zz_dataOut_payload_0_8669 ? _zz_dataOut_payload_0_8603 : _zz_dataOut_payload_0_8615);
  assign _zz_dataOut_payload_0_8671 = (_zz_dataOut_payload_0_8669 ? _zz_dataOut_payload_0_8615 : _zz_dataOut_payload_0_8603);
  assign _zz_dataOut_payload_0_8672 = (_zz_dataOut_payload_0_8661 < _zz_dataOut_payload_0_8667);
  assign _zz_dataOut_payload_0_8673 = (_zz_dataOut_payload_0_8672 ? _zz_dataOut_payload_0_8661 : _zz_dataOut_payload_0_8667);
  assign _zz_dataOut_payload_0_8674 = (_zz_dataOut_payload_0_8672 ? _zz_dataOut_payload_0_8667 : _zz_dataOut_payload_0_8661);
  assign _zz_dataOut_payload_0_8675 = (_zz_dataOut_payload_0_8664 < _zz_dataOut_payload_0_8670);
  assign _zz_dataOut_payload_0_8676 = (_zz_dataOut_payload_0_8675 ? _zz_dataOut_payload_0_8664 : _zz_dataOut_payload_0_8670);
  assign _zz_dataOut_payload_0_8677 = (_zz_dataOut_payload_0_8675 ? _zz_dataOut_payload_0_8670 : _zz_dataOut_payload_0_8664);
  assign _zz_dataOut_payload_0_8678 = (_zz_dataOut_payload_0_8673 < _zz_dataOut_payload_0_8676);
  assign _zz_dataOut_payload_0_8679 = (_zz_dataOut_payload_0_8674 < _zz_dataOut_payload_0_8677);
  assign _zz_dataOut_payload_0_8684 = (_zz_dataOut_payload_0_8662 < _zz_dataOut_payload_0_8668);
  assign _zz_dataOut_payload_0_8685 = (_zz_dataOut_payload_0_8684 ? _zz_dataOut_payload_0_8662 : _zz_dataOut_payload_0_8668);
  assign _zz_dataOut_payload_0_8686 = (_zz_dataOut_payload_0_8684 ? _zz_dataOut_payload_0_8668 : _zz_dataOut_payload_0_8662);
  assign _zz_dataOut_payload_0_8687 = (_zz_dataOut_payload_0_8665 < _zz_dataOut_payload_0_8671);
  assign _zz_dataOut_payload_0_8688 = (_zz_dataOut_payload_0_8687 ? _zz_dataOut_payload_0_8665 : _zz_dataOut_payload_0_8671);
  assign _zz_dataOut_payload_0_8689 = (_zz_dataOut_payload_0_8687 ? _zz_dataOut_payload_0_8671 : _zz_dataOut_payload_0_8665);
  assign _zz_dataOut_payload_0_8690 = (_zz_dataOut_payload_0_8685 < _zz_dataOut_payload_0_8688);
  assign _zz_dataOut_payload_0_8691 = (_zz_dataOut_payload_0_8686 < _zz_dataOut_payload_0_8689);
  assign _zz_dataOut_payload_0_8752 = (_zz_dataOut_payload_0_8415 < _zz_dataOut_payload_0_8367);
  assign _zz_dataOut_payload_0_8753 = (_zz_dataOut_payload_0_8752 ? _zz_dataOut_payload_0_8415 : _zz_dataOut_payload_0_8367);
  assign _zz_dataOut_payload_0_8754 = (_zz_dataOut_payload_0_8752 ? _zz_dataOut_payload_0_8367 : _zz_dataOut_payload_0_8415);
  assign _zz_dataOut_payload_0_8755 = (_zz_dataOut_payload_0_8412 < _zz_dataOut_payload_0_8364);
  assign _zz_dataOut_payload_0_8756 = (_zz_dataOut_payload_0_8755 ? _zz_dataOut_payload_0_8412 : _zz_dataOut_payload_0_8364);
  assign _zz_dataOut_payload_0_8757 = (_zz_dataOut_payload_0_8755 ? _zz_dataOut_payload_0_8364 : _zz_dataOut_payload_0_8412);
  assign _zz_dataOut_payload_0_8758 = (_zz_dataOut_payload_0_8409 < _zz_dataOut_payload_0_8361);
  assign _zz_dataOut_payload_0_8759 = (_zz_dataOut_payload_0_8758 ? _zz_dataOut_payload_0_8409 : _zz_dataOut_payload_0_8361);
  assign _zz_dataOut_payload_0_8760 = (_zz_dataOut_payload_0_8758 ? _zz_dataOut_payload_0_8361 : _zz_dataOut_payload_0_8409);
  assign _zz_dataOut_payload_0_8761 = (_zz_dataOut_payload_0_8406 < _zz_dataOut_payload_0_8358);
  assign _zz_dataOut_payload_0_8762 = (_zz_dataOut_payload_0_8761 ? _zz_dataOut_payload_0_8406 : _zz_dataOut_payload_0_8358);
  assign _zz_dataOut_payload_0_8763 = (_zz_dataOut_payload_0_8761 ? _zz_dataOut_payload_0_8358 : _zz_dataOut_payload_0_8406);
  assign _zz_dataOut_payload_0_8764 = (_zz_dataOut_payload_0_8403 < _zz_dataOut_payload_0_8355);
  assign _zz_dataOut_payload_0_8765 = (_zz_dataOut_payload_0_8764 ? _zz_dataOut_payload_0_8403 : _zz_dataOut_payload_0_8355);
  assign _zz_dataOut_payload_0_8766 = (_zz_dataOut_payload_0_8764 ? _zz_dataOut_payload_0_8355 : _zz_dataOut_payload_0_8403);
  assign _zz_dataOut_payload_0_8767 = (_zz_dataOut_payload_0_8400 < _zz_dataOut_payload_0_8352);
  assign _zz_dataOut_payload_0_8768 = (_zz_dataOut_payload_0_8767 ? _zz_dataOut_payload_0_8400 : _zz_dataOut_payload_0_8352);
  assign _zz_dataOut_payload_0_8769 = (_zz_dataOut_payload_0_8767 ? _zz_dataOut_payload_0_8352 : _zz_dataOut_payload_0_8400);
  assign _zz_dataOut_payload_0_8770 = (_zz_dataOut_payload_0_8397 < _zz_dataOut_payload_0_8349);
  assign _zz_dataOut_payload_0_8771 = (_zz_dataOut_payload_0_8770 ? _zz_dataOut_payload_0_8397 : _zz_dataOut_payload_0_8349);
  assign _zz_dataOut_payload_0_8772 = (_zz_dataOut_payload_0_8770 ? _zz_dataOut_payload_0_8349 : _zz_dataOut_payload_0_8397);
  assign _zz_dataOut_payload_0_8773 = (_zz_dataOut_payload_0_8394 < _zz_dataOut_payload_0_8346);
  assign _zz_dataOut_payload_0_8774 = (_zz_dataOut_payload_0_8773 ? _zz_dataOut_payload_0_8394 : _zz_dataOut_payload_0_8346);
  assign _zz_dataOut_payload_0_8775 = (_zz_dataOut_payload_0_8773 ? _zz_dataOut_payload_0_8346 : _zz_dataOut_payload_0_8394);
  assign _zz_dataOut_payload_0_8776 = (_zz_dataOut_payload_0_8391 < _zz_dataOut_payload_0_8343);
  assign _zz_dataOut_payload_0_8777 = (_zz_dataOut_payload_0_8776 ? _zz_dataOut_payload_0_8391 : _zz_dataOut_payload_0_8343);
  assign _zz_dataOut_payload_0_8778 = (_zz_dataOut_payload_0_8776 ? _zz_dataOut_payload_0_8343 : _zz_dataOut_payload_0_8391);
  assign _zz_dataOut_payload_0_8779 = (_zz_dataOut_payload_0_8388 < _zz_dataOut_payload_0_8340);
  assign _zz_dataOut_payload_0_8780 = (_zz_dataOut_payload_0_8779 ? _zz_dataOut_payload_0_8388 : _zz_dataOut_payload_0_8340);
  assign _zz_dataOut_payload_0_8781 = (_zz_dataOut_payload_0_8779 ? _zz_dataOut_payload_0_8340 : _zz_dataOut_payload_0_8388);
  assign _zz_dataOut_payload_0_8782 = (_zz_dataOut_payload_0_8385 < _zz_dataOut_payload_0_8337);
  assign _zz_dataOut_payload_0_8783 = (_zz_dataOut_payload_0_8782 ? _zz_dataOut_payload_0_8385 : _zz_dataOut_payload_0_8337);
  assign _zz_dataOut_payload_0_8784 = (_zz_dataOut_payload_0_8782 ? _zz_dataOut_payload_0_8337 : _zz_dataOut_payload_0_8385);
  assign _zz_dataOut_payload_0_8785 = (_zz_dataOut_payload_0_8382 < _zz_dataOut_payload_0_8334);
  assign _zz_dataOut_payload_0_8786 = (_zz_dataOut_payload_0_8785 ? _zz_dataOut_payload_0_8382 : _zz_dataOut_payload_0_8334);
  assign _zz_dataOut_payload_0_8787 = (_zz_dataOut_payload_0_8785 ? _zz_dataOut_payload_0_8334 : _zz_dataOut_payload_0_8382);
  assign _zz_dataOut_payload_0_8788 = (_zz_dataOut_payload_0_8379 < _zz_dataOut_payload_0_8331);
  assign _zz_dataOut_payload_0_8789 = (_zz_dataOut_payload_0_8788 ? _zz_dataOut_payload_0_8379 : _zz_dataOut_payload_0_8331);
  assign _zz_dataOut_payload_0_8790 = (_zz_dataOut_payload_0_8788 ? _zz_dataOut_payload_0_8331 : _zz_dataOut_payload_0_8379);
  assign _zz_dataOut_payload_0_8791 = (_zz_dataOut_payload_0_8376 < _zz_dataOut_payload_0_8328);
  assign _zz_dataOut_payload_0_8792 = (_zz_dataOut_payload_0_8791 ? _zz_dataOut_payload_0_8376 : _zz_dataOut_payload_0_8328);
  assign _zz_dataOut_payload_0_8793 = (_zz_dataOut_payload_0_8791 ? _zz_dataOut_payload_0_8328 : _zz_dataOut_payload_0_8376);
  assign _zz_dataOut_payload_0_8794 = (_zz_dataOut_payload_0_8373 < _zz_dataOut_payload_0_8325);
  assign _zz_dataOut_payload_0_8795 = (_zz_dataOut_payload_0_8794 ? _zz_dataOut_payload_0_8373 : _zz_dataOut_payload_0_8325);
  assign _zz_dataOut_payload_0_8796 = (_zz_dataOut_payload_0_8794 ? _zz_dataOut_payload_0_8325 : _zz_dataOut_payload_0_8373);
  assign _zz_dataOut_payload_0_8797 = (_zz_dataOut_payload_0_8370 < _zz_dataOut_payload_0_8322);
  assign _zz_dataOut_payload_0_8798 = (_zz_dataOut_payload_0_8797 ? _zz_dataOut_payload_0_8370 : _zz_dataOut_payload_0_8322);
  assign _zz_dataOut_payload_0_8799 = (_zz_dataOut_payload_0_8797 ? _zz_dataOut_payload_0_8322 : _zz_dataOut_payload_0_8370);
  assign _zz_dataOut_payload_0_8800 = (_zz_dataOut_payload_0_8753 < _zz_dataOut_payload_0_8777);
  assign _zz_dataOut_payload_0_8801 = (_zz_dataOut_payload_0_8800 ? _zz_dataOut_payload_0_8753 : _zz_dataOut_payload_0_8777);
  assign _zz_dataOut_payload_0_8802 = (_zz_dataOut_payload_0_8800 ? _zz_dataOut_payload_0_8777 : _zz_dataOut_payload_0_8753);
  assign _zz_dataOut_payload_0_8803 = (_zz_dataOut_payload_0_8756 < _zz_dataOut_payload_0_8780);
  assign _zz_dataOut_payload_0_8804 = (_zz_dataOut_payload_0_8803 ? _zz_dataOut_payload_0_8756 : _zz_dataOut_payload_0_8780);
  assign _zz_dataOut_payload_0_8805 = (_zz_dataOut_payload_0_8803 ? _zz_dataOut_payload_0_8780 : _zz_dataOut_payload_0_8756);
  assign _zz_dataOut_payload_0_8806 = (_zz_dataOut_payload_0_8759 < _zz_dataOut_payload_0_8783);
  assign _zz_dataOut_payload_0_8807 = (_zz_dataOut_payload_0_8806 ? _zz_dataOut_payload_0_8759 : _zz_dataOut_payload_0_8783);
  assign _zz_dataOut_payload_0_8808 = (_zz_dataOut_payload_0_8806 ? _zz_dataOut_payload_0_8783 : _zz_dataOut_payload_0_8759);
  assign _zz_dataOut_payload_0_8809 = (_zz_dataOut_payload_0_8762 < _zz_dataOut_payload_0_8786);
  assign _zz_dataOut_payload_0_8810 = (_zz_dataOut_payload_0_8809 ? _zz_dataOut_payload_0_8762 : _zz_dataOut_payload_0_8786);
  assign _zz_dataOut_payload_0_8811 = (_zz_dataOut_payload_0_8809 ? _zz_dataOut_payload_0_8786 : _zz_dataOut_payload_0_8762);
  assign _zz_dataOut_payload_0_8812 = (_zz_dataOut_payload_0_8765 < _zz_dataOut_payload_0_8789);
  assign _zz_dataOut_payload_0_8813 = (_zz_dataOut_payload_0_8812 ? _zz_dataOut_payload_0_8765 : _zz_dataOut_payload_0_8789);
  assign _zz_dataOut_payload_0_8814 = (_zz_dataOut_payload_0_8812 ? _zz_dataOut_payload_0_8789 : _zz_dataOut_payload_0_8765);
  assign _zz_dataOut_payload_0_8815 = (_zz_dataOut_payload_0_8768 < _zz_dataOut_payload_0_8792);
  assign _zz_dataOut_payload_0_8816 = (_zz_dataOut_payload_0_8815 ? _zz_dataOut_payload_0_8768 : _zz_dataOut_payload_0_8792);
  assign _zz_dataOut_payload_0_8817 = (_zz_dataOut_payload_0_8815 ? _zz_dataOut_payload_0_8792 : _zz_dataOut_payload_0_8768);
  assign _zz_dataOut_payload_0_8818 = (_zz_dataOut_payload_0_8771 < _zz_dataOut_payload_0_8795);
  assign _zz_dataOut_payload_0_8819 = (_zz_dataOut_payload_0_8818 ? _zz_dataOut_payload_0_8771 : _zz_dataOut_payload_0_8795);
  assign _zz_dataOut_payload_0_8820 = (_zz_dataOut_payload_0_8818 ? _zz_dataOut_payload_0_8795 : _zz_dataOut_payload_0_8771);
  assign _zz_dataOut_payload_0_8821 = (_zz_dataOut_payload_0_8774 < _zz_dataOut_payload_0_8798);
  assign _zz_dataOut_payload_0_8822 = (_zz_dataOut_payload_0_8821 ? _zz_dataOut_payload_0_8774 : _zz_dataOut_payload_0_8798);
  assign _zz_dataOut_payload_0_8823 = (_zz_dataOut_payload_0_8821 ? _zz_dataOut_payload_0_8798 : _zz_dataOut_payload_0_8774);
  assign _zz_dataOut_payload_0_8824 = (_zz_dataOut_payload_0_8801 < _zz_dataOut_payload_0_8813);
  assign _zz_dataOut_payload_0_8825 = (_zz_dataOut_payload_0_8824 ? _zz_dataOut_payload_0_8801 : _zz_dataOut_payload_0_8813);
  assign _zz_dataOut_payload_0_8826 = (_zz_dataOut_payload_0_8824 ? _zz_dataOut_payload_0_8813 : _zz_dataOut_payload_0_8801);
  assign _zz_dataOut_payload_0_8827 = (_zz_dataOut_payload_0_8804 < _zz_dataOut_payload_0_8816);
  assign _zz_dataOut_payload_0_8828 = (_zz_dataOut_payload_0_8827 ? _zz_dataOut_payload_0_8804 : _zz_dataOut_payload_0_8816);
  assign _zz_dataOut_payload_0_8829 = (_zz_dataOut_payload_0_8827 ? _zz_dataOut_payload_0_8816 : _zz_dataOut_payload_0_8804);
  assign _zz_dataOut_payload_0_8830 = (_zz_dataOut_payload_0_8807 < _zz_dataOut_payload_0_8819);
  assign _zz_dataOut_payload_0_8831 = (_zz_dataOut_payload_0_8830 ? _zz_dataOut_payload_0_8807 : _zz_dataOut_payload_0_8819);
  assign _zz_dataOut_payload_0_8832 = (_zz_dataOut_payload_0_8830 ? _zz_dataOut_payload_0_8819 : _zz_dataOut_payload_0_8807);
  assign _zz_dataOut_payload_0_8833 = (_zz_dataOut_payload_0_8810 < _zz_dataOut_payload_0_8822);
  assign _zz_dataOut_payload_0_8834 = (_zz_dataOut_payload_0_8833 ? _zz_dataOut_payload_0_8810 : _zz_dataOut_payload_0_8822);
  assign _zz_dataOut_payload_0_8835 = (_zz_dataOut_payload_0_8833 ? _zz_dataOut_payload_0_8822 : _zz_dataOut_payload_0_8810);
  assign _zz_dataOut_payload_0_8836 = (_zz_dataOut_payload_0_8825 < _zz_dataOut_payload_0_8831);
  assign _zz_dataOut_payload_0_8837 = (_zz_dataOut_payload_0_8836 ? _zz_dataOut_payload_0_8825 : _zz_dataOut_payload_0_8831);
  assign _zz_dataOut_payload_0_8838 = (_zz_dataOut_payload_0_8836 ? _zz_dataOut_payload_0_8831 : _zz_dataOut_payload_0_8825);
  assign _zz_dataOut_payload_0_8839 = (_zz_dataOut_payload_0_8828 < _zz_dataOut_payload_0_8834);
  assign _zz_dataOut_payload_0_8840 = (_zz_dataOut_payload_0_8839 ? _zz_dataOut_payload_0_8828 : _zz_dataOut_payload_0_8834);
  assign _zz_dataOut_payload_0_8841 = (_zz_dataOut_payload_0_8839 ? _zz_dataOut_payload_0_8834 : _zz_dataOut_payload_0_8828);
  assign _zz_dataOut_payload_0_8842 = (_zz_dataOut_payload_0_8837 < _zz_dataOut_payload_0_8840);
  assign _zz_dataOut_payload_0_8843 = (_zz_dataOut_payload_0_8838 < _zz_dataOut_payload_0_8841);
  assign _zz_dataOut_payload_0_8848 = (_zz_dataOut_payload_0_8826 < _zz_dataOut_payload_0_8832);
  assign _zz_dataOut_payload_0_8849 = (_zz_dataOut_payload_0_8848 ? _zz_dataOut_payload_0_8826 : _zz_dataOut_payload_0_8832);
  assign _zz_dataOut_payload_0_8850 = (_zz_dataOut_payload_0_8848 ? _zz_dataOut_payload_0_8832 : _zz_dataOut_payload_0_8826);
  assign _zz_dataOut_payload_0_8851 = (_zz_dataOut_payload_0_8829 < _zz_dataOut_payload_0_8835);
  assign _zz_dataOut_payload_0_8852 = (_zz_dataOut_payload_0_8851 ? _zz_dataOut_payload_0_8829 : _zz_dataOut_payload_0_8835);
  assign _zz_dataOut_payload_0_8853 = (_zz_dataOut_payload_0_8851 ? _zz_dataOut_payload_0_8835 : _zz_dataOut_payload_0_8829);
  assign _zz_dataOut_payload_0_8854 = (_zz_dataOut_payload_0_8849 < _zz_dataOut_payload_0_8852);
  assign _zz_dataOut_payload_0_8855 = (_zz_dataOut_payload_0_8850 < _zz_dataOut_payload_0_8853);
  assign _zz_dataOut_payload_0_8868 = (_zz_dataOut_payload_0_8802 < _zz_dataOut_payload_0_8814);
  assign _zz_dataOut_payload_0_8869 = (_zz_dataOut_payload_0_8868 ? _zz_dataOut_payload_0_8802 : _zz_dataOut_payload_0_8814);
  assign _zz_dataOut_payload_0_8870 = (_zz_dataOut_payload_0_8868 ? _zz_dataOut_payload_0_8814 : _zz_dataOut_payload_0_8802);
  assign _zz_dataOut_payload_0_8871 = (_zz_dataOut_payload_0_8805 < _zz_dataOut_payload_0_8817);
  assign _zz_dataOut_payload_0_8872 = (_zz_dataOut_payload_0_8871 ? _zz_dataOut_payload_0_8805 : _zz_dataOut_payload_0_8817);
  assign _zz_dataOut_payload_0_8873 = (_zz_dataOut_payload_0_8871 ? _zz_dataOut_payload_0_8817 : _zz_dataOut_payload_0_8805);
  assign _zz_dataOut_payload_0_8874 = (_zz_dataOut_payload_0_8808 < _zz_dataOut_payload_0_8820);
  assign _zz_dataOut_payload_0_8875 = (_zz_dataOut_payload_0_8874 ? _zz_dataOut_payload_0_8808 : _zz_dataOut_payload_0_8820);
  assign _zz_dataOut_payload_0_8876 = (_zz_dataOut_payload_0_8874 ? _zz_dataOut_payload_0_8820 : _zz_dataOut_payload_0_8808);
  assign _zz_dataOut_payload_0_8877 = (_zz_dataOut_payload_0_8811 < _zz_dataOut_payload_0_8823);
  assign _zz_dataOut_payload_0_8878 = (_zz_dataOut_payload_0_8877 ? _zz_dataOut_payload_0_8811 : _zz_dataOut_payload_0_8823);
  assign _zz_dataOut_payload_0_8879 = (_zz_dataOut_payload_0_8877 ? _zz_dataOut_payload_0_8823 : _zz_dataOut_payload_0_8811);
  assign _zz_dataOut_payload_0_8880 = (_zz_dataOut_payload_0_8869 < _zz_dataOut_payload_0_8875);
  assign _zz_dataOut_payload_0_8881 = (_zz_dataOut_payload_0_8880 ? _zz_dataOut_payload_0_8869 : _zz_dataOut_payload_0_8875);
  assign _zz_dataOut_payload_0_8882 = (_zz_dataOut_payload_0_8880 ? _zz_dataOut_payload_0_8875 : _zz_dataOut_payload_0_8869);
  assign _zz_dataOut_payload_0_8883 = (_zz_dataOut_payload_0_8872 < _zz_dataOut_payload_0_8878);
  assign _zz_dataOut_payload_0_8884 = (_zz_dataOut_payload_0_8883 ? _zz_dataOut_payload_0_8872 : _zz_dataOut_payload_0_8878);
  assign _zz_dataOut_payload_0_8885 = (_zz_dataOut_payload_0_8883 ? _zz_dataOut_payload_0_8878 : _zz_dataOut_payload_0_8872);
  assign _zz_dataOut_payload_0_8886 = (_zz_dataOut_payload_0_8881 < _zz_dataOut_payload_0_8884);
  assign _zz_dataOut_payload_0_8887 = (_zz_dataOut_payload_0_8882 < _zz_dataOut_payload_0_8885);
  assign _zz_dataOut_payload_0_8892 = (_zz_dataOut_payload_0_8870 < _zz_dataOut_payload_0_8876);
  assign _zz_dataOut_payload_0_8893 = (_zz_dataOut_payload_0_8892 ? _zz_dataOut_payload_0_8870 : _zz_dataOut_payload_0_8876);
  assign _zz_dataOut_payload_0_8894 = (_zz_dataOut_payload_0_8892 ? _zz_dataOut_payload_0_8876 : _zz_dataOut_payload_0_8870);
  assign _zz_dataOut_payload_0_8895 = (_zz_dataOut_payload_0_8873 < _zz_dataOut_payload_0_8879);
  assign _zz_dataOut_payload_0_8896 = (_zz_dataOut_payload_0_8895 ? _zz_dataOut_payload_0_8873 : _zz_dataOut_payload_0_8879);
  assign _zz_dataOut_payload_0_8897 = (_zz_dataOut_payload_0_8895 ? _zz_dataOut_payload_0_8879 : _zz_dataOut_payload_0_8873);
  assign _zz_dataOut_payload_0_8898 = (_zz_dataOut_payload_0_8893 < _zz_dataOut_payload_0_8896);
  assign _zz_dataOut_payload_0_8899 = (_zz_dataOut_payload_0_8894 < _zz_dataOut_payload_0_8897);
  assign _zz_dataOut_payload_0_8928 = (_zz_dataOut_payload_0_8754 < _zz_dataOut_payload_0_8778);
  assign _zz_dataOut_payload_0_8929 = (_zz_dataOut_payload_0_8928 ? _zz_dataOut_payload_0_8754 : _zz_dataOut_payload_0_8778);
  assign _zz_dataOut_payload_0_8930 = (_zz_dataOut_payload_0_8928 ? _zz_dataOut_payload_0_8778 : _zz_dataOut_payload_0_8754);
  assign _zz_dataOut_payload_0_8931 = (_zz_dataOut_payload_0_8757 < _zz_dataOut_payload_0_8781);
  assign _zz_dataOut_payload_0_8932 = (_zz_dataOut_payload_0_8931 ? _zz_dataOut_payload_0_8757 : _zz_dataOut_payload_0_8781);
  assign _zz_dataOut_payload_0_8933 = (_zz_dataOut_payload_0_8931 ? _zz_dataOut_payload_0_8781 : _zz_dataOut_payload_0_8757);
  assign _zz_dataOut_payload_0_8934 = (_zz_dataOut_payload_0_8760 < _zz_dataOut_payload_0_8784);
  assign _zz_dataOut_payload_0_8935 = (_zz_dataOut_payload_0_8934 ? _zz_dataOut_payload_0_8760 : _zz_dataOut_payload_0_8784);
  assign _zz_dataOut_payload_0_8936 = (_zz_dataOut_payload_0_8934 ? _zz_dataOut_payload_0_8784 : _zz_dataOut_payload_0_8760);
  assign _zz_dataOut_payload_0_8937 = (_zz_dataOut_payload_0_8763 < _zz_dataOut_payload_0_8787);
  assign _zz_dataOut_payload_0_8938 = (_zz_dataOut_payload_0_8937 ? _zz_dataOut_payload_0_8763 : _zz_dataOut_payload_0_8787);
  assign _zz_dataOut_payload_0_8939 = (_zz_dataOut_payload_0_8937 ? _zz_dataOut_payload_0_8787 : _zz_dataOut_payload_0_8763);
  assign _zz_dataOut_payload_0_8940 = (_zz_dataOut_payload_0_8766 < _zz_dataOut_payload_0_8790);
  assign _zz_dataOut_payload_0_8941 = (_zz_dataOut_payload_0_8940 ? _zz_dataOut_payload_0_8766 : _zz_dataOut_payload_0_8790);
  assign _zz_dataOut_payload_0_8942 = (_zz_dataOut_payload_0_8940 ? _zz_dataOut_payload_0_8790 : _zz_dataOut_payload_0_8766);
  assign _zz_dataOut_payload_0_8943 = (_zz_dataOut_payload_0_8769 < _zz_dataOut_payload_0_8793);
  assign _zz_dataOut_payload_0_8944 = (_zz_dataOut_payload_0_8943 ? _zz_dataOut_payload_0_8769 : _zz_dataOut_payload_0_8793);
  assign _zz_dataOut_payload_0_8945 = (_zz_dataOut_payload_0_8943 ? _zz_dataOut_payload_0_8793 : _zz_dataOut_payload_0_8769);
  assign _zz_dataOut_payload_0_8946 = (_zz_dataOut_payload_0_8772 < _zz_dataOut_payload_0_8796);
  assign _zz_dataOut_payload_0_8947 = (_zz_dataOut_payload_0_8946 ? _zz_dataOut_payload_0_8772 : _zz_dataOut_payload_0_8796);
  assign _zz_dataOut_payload_0_8948 = (_zz_dataOut_payload_0_8946 ? _zz_dataOut_payload_0_8796 : _zz_dataOut_payload_0_8772);
  assign _zz_dataOut_payload_0_8949 = (_zz_dataOut_payload_0_8775 < _zz_dataOut_payload_0_8799);
  assign _zz_dataOut_payload_0_8950 = (_zz_dataOut_payload_0_8949 ? _zz_dataOut_payload_0_8775 : _zz_dataOut_payload_0_8799);
  assign _zz_dataOut_payload_0_8951 = (_zz_dataOut_payload_0_8949 ? _zz_dataOut_payload_0_8799 : _zz_dataOut_payload_0_8775);
  assign _zz_dataOut_payload_0_8952 = (_zz_dataOut_payload_0_8929 < _zz_dataOut_payload_0_8941);
  assign _zz_dataOut_payload_0_8953 = (_zz_dataOut_payload_0_8952 ? _zz_dataOut_payload_0_8929 : _zz_dataOut_payload_0_8941);
  assign _zz_dataOut_payload_0_8954 = (_zz_dataOut_payload_0_8952 ? _zz_dataOut_payload_0_8941 : _zz_dataOut_payload_0_8929);
  assign _zz_dataOut_payload_0_8955 = (_zz_dataOut_payload_0_8932 < _zz_dataOut_payload_0_8944);
  assign _zz_dataOut_payload_0_8956 = (_zz_dataOut_payload_0_8955 ? _zz_dataOut_payload_0_8932 : _zz_dataOut_payload_0_8944);
  assign _zz_dataOut_payload_0_8957 = (_zz_dataOut_payload_0_8955 ? _zz_dataOut_payload_0_8944 : _zz_dataOut_payload_0_8932);
  assign _zz_dataOut_payload_0_8958 = (_zz_dataOut_payload_0_8935 < _zz_dataOut_payload_0_8947);
  assign _zz_dataOut_payload_0_8959 = (_zz_dataOut_payload_0_8958 ? _zz_dataOut_payload_0_8935 : _zz_dataOut_payload_0_8947);
  assign _zz_dataOut_payload_0_8960 = (_zz_dataOut_payload_0_8958 ? _zz_dataOut_payload_0_8947 : _zz_dataOut_payload_0_8935);
  assign _zz_dataOut_payload_0_8961 = (_zz_dataOut_payload_0_8938 < _zz_dataOut_payload_0_8950);
  assign _zz_dataOut_payload_0_8962 = (_zz_dataOut_payload_0_8961 ? _zz_dataOut_payload_0_8938 : _zz_dataOut_payload_0_8950);
  assign _zz_dataOut_payload_0_8963 = (_zz_dataOut_payload_0_8961 ? _zz_dataOut_payload_0_8950 : _zz_dataOut_payload_0_8938);
  assign _zz_dataOut_payload_0_8964 = (_zz_dataOut_payload_0_8953 < _zz_dataOut_payload_0_8959);
  assign _zz_dataOut_payload_0_8965 = (_zz_dataOut_payload_0_8964 ? _zz_dataOut_payload_0_8953 : _zz_dataOut_payload_0_8959);
  assign _zz_dataOut_payload_0_8966 = (_zz_dataOut_payload_0_8964 ? _zz_dataOut_payload_0_8959 : _zz_dataOut_payload_0_8953);
  assign _zz_dataOut_payload_0_8967 = (_zz_dataOut_payload_0_8956 < _zz_dataOut_payload_0_8962);
  assign _zz_dataOut_payload_0_8968 = (_zz_dataOut_payload_0_8967 ? _zz_dataOut_payload_0_8956 : _zz_dataOut_payload_0_8962);
  assign _zz_dataOut_payload_0_8969 = (_zz_dataOut_payload_0_8967 ? _zz_dataOut_payload_0_8962 : _zz_dataOut_payload_0_8956);
  assign _zz_dataOut_payload_0_8970 = (_zz_dataOut_payload_0_8965 < _zz_dataOut_payload_0_8968);
  assign _zz_dataOut_payload_0_8971 = (_zz_dataOut_payload_0_8966 < _zz_dataOut_payload_0_8969);
  assign _zz_dataOut_payload_0_8976 = (_zz_dataOut_payload_0_8954 < _zz_dataOut_payload_0_8960);
  assign _zz_dataOut_payload_0_8977 = (_zz_dataOut_payload_0_8976 ? _zz_dataOut_payload_0_8954 : _zz_dataOut_payload_0_8960);
  assign _zz_dataOut_payload_0_8978 = (_zz_dataOut_payload_0_8976 ? _zz_dataOut_payload_0_8960 : _zz_dataOut_payload_0_8954);
  assign _zz_dataOut_payload_0_8979 = (_zz_dataOut_payload_0_8957 < _zz_dataOut_payload_0_8963);
  assign _zz_dataOut_payload_0_8980 = (_zz_dataOut_payload_0_8979 ? _zz_dataOut_payload_0_8957 : _zz_dataOut_payload_0_8963);
  assign _zz_dataOut_payload_0_8981 = (_zz_dataOut_payload_0_8979 ? _zz_dataOut_payload_0_8963 : _zz_dataOut_payload_0_8957);
  assign _zz_dataOut_payload_0_8982 = (_zz_dataOut_payload_0_8977 < _zz_dataOut_payload_0_8980);
  assign _zz_dataOut_payload_0_8983 = (_zz_dataOut_payload_0_8978 < _zz_dataOut_payload_0_8981);
  assign _zz_dataOut_payload_0_8996 = (_zz_dataOut_payload_0_8930 < _zz_dataOut_payload_0_8942);
  assign _zz_dataOut_payload_0_8997 = (_zz_dataOut_payload_0_8996 ? _zz_dataOut_payload_0_8930 : _zz_dataOut_payload_0_8942);
  assign _zz_dataOut_payload_0_8998 = (_zz_dataOut_payload_0_8996 ? _zz_dataOut_payload_0_8942 : _zz_dataOut_payload_0_8930);
  assign _zz_dataOut_payload_0_8999 = (_zz_dataOut_payload_0_8933 < _zz_dataOut_payload_0_8945);
  assign _zz_dataOut_payload_0_9000 = (_zz_dataOut_payload_0_8999 ? _zz_dataOut_payload_0_8933 : _zz_dataOut_payload_0_8945);
  assign _zz_dataOut_payload_0_9001 = (_zz_dataOut_payload_0_8999 ? _zz_dataOut_payload_0_8945 : _zz_dataOut_payload_0_8933);
  assign _zz_dataOut_payload_0_9002 = (_zz_dataOut_payload_0_8936 < _zz_dataOut_payload_0_8948);
  assign _zz_dataOut_payload_0_9003 = (_zz_dataOut_payload_0_9002 ? _zz_dataOut_payload_0_8936 : _zz_dataOut_payload_0_8948);
  assign _zz_dataOut_payload_0_9004 = (_zz_dataOut_payload_0_9002 ? _zz_dataOut_payload_0_8948 : _zz_dataOut_payload_0_8936);
  assign _zz_dataOut_payload_0_9005 = (_zz_dataOut_payload_0_8939 < _zz_dataOut_payload_0_8951);
  assign _zz_dataOut_payload_0_9006 = (_zz_dataOut_payload_0_9005 ? _zz_dataOut_payload_0_8939 : _zz_dataOut_payload_0_8951);
  assign _zz_dataOut_payload_0_9007 = (_zz_dataOut_payload_0_9005 ? _zz_dataOut_payload_0_8951 : _zz_dataOut_payload_0_8939);
  assign _zz_dataOut_payload_0_9008 = (_zz_dataOut_payload_0_8997 < _zz_dataOut_payload_0_9003);
  assign _zz_dataOut_payload_0_9009 = (_zz_dataOut_payload_0_9008 ? _zz_dataOut_payload_0_8997 : _zz_dataOut_payload_0_9003);
  assign _zz_dataOut_payload_0_9010 = (_zz_dataOut_payload_0_9008 ? _zz_dataOut_payload_0_9003 : _zz_dataOut_payload_0_8997);
  assign _zz_dataOut_payload_0_9011 = (_zz_dataOut_payload_0_9000 < _zz_dataOut_payload_0_9006);
  assign _zz_dataOut_payload_0_9012 = (_zz_dataOut_payload_0_9011 ? _zz_dataOut_payload_0_9000 : _zz_dataOut_payload_0_9006);
  assign _zz_dataOut_payload_0_9013 = (_zz_dataOut_payload_0_9011 ? _zz_dataOut_payload_0_9006 : _zz_dataOut_payload_0_9000);
  assign _zz_dataOut_payload_0_9014 = (_zz_dataOut_payload_0_9009 < _zz_dataOut_payload_0_9012);
  assign _zz_dataOut_payload_0_9015 = (_zz_dataOut_payload_0_9010 < _zz_dataOut_payload_0_9013);
  assign _zz_dataOut_payload_0_9020 = (_zz_dataOut_payload_0_8998 < _zz_dataOut_payload_0_9004);
  assign _zz_dataOut_payload_0_9021 = (_zz_dataOut_payload_0_9020 ? _zz_dataOut_payload_0_8998 : _zz_dataOut_payload_0_9004);
  assign _zz_dataOut_payload_0_9022 = (_zz_dataOut_payload_0_9020 ? _zz_dataOut_payload_0_9004 : _zz_dataOut_payload_0_8998);
  assign _zz_dataOut_payload_0_9023 = (_zz_dataOut_payload_0_9001 < _zz_dataOut_payload_0_9007);
  assign _zz_dataOut_payload_0_9024 = (_zz_dataOut_payload_0_9023 ? _zz_dataOut_payload_0_9001 : _zz_dataOut_payload_0_9007);
  assign _zz_dataOut_payload_0_9025 = (_zz_dataOut_payload_0_9023 ? _zz_dataOut_payload_0_9007 : _zz_dataOut_payload_0_9001);
  assign _zz_dataOut_payload_0_9026 = (_zz_dataOut_payload_0_9021 < _zz_dataOut_payload_0_9024);
  assign _zz_dataOut_payload_0_9027 = (_zz_dataOut_payload_0_9022 < _zz_dataOut_payload_0_9025);
  assign _zz_dataOut_payload_0_9152 = (_zz_dataOut_payload_0_8128 < _zz_dataOut_payload_0_8191);
  assign _zz_dataOut_payload_0_9153 = (_zz_dataOut_payload_0_9152 ? _zz_dataOut_payload_0_8128 : _zz_dataOut_payload_0_8191);
  assign _zz_dataOut_payload_0_9154 = (_zz_dataOut_payload_0_9152 ? _zz_dataOut_payload_0_8191 : _zz_dataOut_payload_0_8128);
  assign _zz_dataOut_payload_0_9155 = (_zz_dataOut_payload_0_8129 < _zz_dataOut_payload_0_8190);
  assign _zz_dataOut_payload_0_9156 = (_zz_dataOut_payload_0_9155 ? _zz_dataOut_payload_0_8129 : _zz_dataOut_payload_0_8190);
  assign _zz_dataOut_payload_0_9157 = (_zz_dataOut_payload_0_9155 ? _zz_dataOut_payload_0_8190 : _zz_dataOut_payload_0_8129);
  assign _zz_dataOut_payload_0_9158 = (_zz_dataOut_payload_0_8130 < _zz_dataOut_payload_0_8189);
  assign _zz_dataOut_payload_0_9159 = (_zz_dataOut_payload_0_9158 ? _zz_dataOut_payload_0_8130 : _zz_dataOut_payload_0_8189);
  assign _zz_dataOut_payload_0_9160 = (_zz_dataOut_payload_0_9158 ? _zz_dataOut_payload_0_8189 : _zz_dataOut_payload_0_8130);
  assign _zz_dataOut_payload_0_9161 = (_zz_dataOut_payload_0_8131 < _zz_dataOut_payload_0_8188);
  assign _zz_dataOut_payload_0_9162 = (_zz_dataOut_payload_0_9161 ? _zz_dataOut_payload_0_8131 : _zz_dataOut_payload_0_8188);
  assign _zz_dataOut_payload_0_9163 = (_zz_dataOut_payload_0_9161 ? _zz_dataOut_payload_0_8188 : _zz_dataOut_payload_0_8131);
  assign _zz_dataOut_payload_0_9164 = (_zz_dataOut_payload_0_8132 < _zz_dataOut_payload_0_8187);
  assign _zz_dataOut_payload_0_9165 = (_zz_dataOut_payload_0_9164 ? _zz_dataOut_payload_0_8132 : _zz_dataOut_payload_0_8187);
  assign _zz_dataOut_payload_0_9166 = (_zz_dataOut_payload_0_9164 ? _zz_dataOut_payload_0_8187 : _zz_dataOut_payload_0_8132);
  assign _zz_dataOut_payload_0_9167 = (_zz_dataOut_payload_0_8133 < _zz_dataOut_payload_0_8186);
  assign _zz_dataOut_payload_0_9168 = (_zz_dataOut_payload_0_9167 ? _zz_dataOut_payload_0_8133 : _zz_dataOut_payload_0_8186);
  assign _zz_dataOut_payload_0_9169 = (_zz_dataOut_payload_0_9167 ? _zz_dataOut_payload_0_8186 : _zz_dataOut_payload_0_8133);
  assign _zz_dataOut_payload_0_9170 = (_zz_dataOut_payload_0_8134 < _zz_dataOut_payload_0_8185);
  assign _zz_dataOut_payload_0_9171 = (_zz_dataOut_payload_0_9170 ? _zz_dataOut_payload_0_8134 : _zz_dataOut_payload_0_8185);
  assign _zz_dataOut_payload_0_9172 = (_zz_dataOut_payload_0_9170 ? _zz_dataOut_payload_0_8185 : _zz_dataOut_payload_0_8134);
  assign _zz_dataOut_payload_0_9173 = (_zz_dataOut_payload_0_8135 < _zz_dataOut_payload_0_8184);
  assign _zz_dataOut_payload_0_9174 = (_zz_dataOut_payload_0_9173 ? _zz_dataOut_payload_0_8135 : _zz_dataOut_payload_0_8184);
  assign _zz_dataOut_payload_0_9175 = (_zz_dataOut_payload_0_9173 ? _zz_dataOut_payload_0_8184 : _zz_dataOut_payload_0_8135);
  assign _zz_dataOut_payload_0_9176 = (_zz_dataOut_payload_0_8136 < _zz_dataOut_payload_0_8183);
  assign _zz_dataOut_payload_0_9177 = (_zz_dataOut_payload_0_9176 ? _zz_dataOut_payload_0_8136 : _zz_dataOut_payload_0_8183);
  assign _zz_dataOut_payload_0_9178 = (_zz_dataOut_payload_0_9176 ? _zz_dataOut_payload_0_8183 : _zz_dataOut_payload_0_8136);
  assign _zz_dataOut_payload_0_9179 = (_zz_dataOut_payload_0_8137 < _zz_dataOut_payload_0_8182);
  assign _zz_dataOut_payload_0_9180 = (_zz_dataOut_payload_0_9179 ? _zz_dataOut_payload_0_8137 : _zz_dataOut_payload_0_8182);
  assign _zz_dataOut_payload_0_9181 = (_zz_dataOut_payload_0_9179 ? _zz_dataOut_payload_0_8182 : _zz_dataOut_payload_0_8137);
  assign _zz_dataOut_payload_0_9182 = (_zz_dataOut_payload_0_8138 < _zz_dataOut_payload_0_8181);
  assign _zz_dataOut_payload_0_9183 = (_zz_dataOut_payload_0_9182 ? _zz_dataOut_payload_0_8138 : _zz_dataOut_payload_0_8181);
  assign _zz_dataOut_payload_0_9184 = (_zz_dataOut_payload_0_9182 ? _zz_dataOut_payload_0_8181 : _zz_dataOut_payload_0_8138);
  assign _zz_dataOut_payload_0_9185 = (_zz_dataOut_payload_0_8139 < _zz_dataOut_payload_0_8180);
  assign _zz_dataOut_payload_0_9186 = (_zz_dataOut_payload_0_9185 ? _zz_dataOut_payload_0_8139 : _zz_dataOut_payload_0_8180);
  assign _zz_dataOut_payload_0_9187 = (_zz_dataOut_payload_0_9185 ? _zz_dataOut_payload_0_8180 : _zz_dataOut_payload_0_8139);
  assign _zz_dataOut_payload_0_9188 = (_zz_dataOut_payload_0_8140 < _zz_dataOut_payload_0_8179);
  assign _zz_dataOut_payload_0_9189 = (_zz_dataOut_payload_0_9188 ? _zz_dataOut_payload_0_8140 : _zz_dataOut_payload_0_8179);
  assign _zz_dataOut_payload_0_9190 = (_zz_dataOut_payload_0_9188 ? _zz_dataOut_payload_0_8179 : _zz_dataOut_payload_0_8140);
  assign _zz_dataOut_payload_0_9191 = (_zz_dataOut_payload_0_8141 < _zz_dataOut_payload_0_8178);
  assign _zz_dataOut_payload_0_9192 = (_zz_dataOut_payload_0_9191 ? _zz_dataOut_payload_0_8141 : _zz_dataOut_payload_0_8178);
  assign _zz_dataOut_payload_0_9193 = (_zz_dataOut_payload_0_9191 ? _zz_dataOut_payload_0_8178 : _zz_dataOut_payload_0_8141);
  assign _zz_dataOut_payload_0_9194 = (_zz_dataOut_payload_0_8142 < _zz_dataOut_payload_0_8177);
  assign _zz_dataOut_payload_0_9195 = (_zz_dataOut_payload_0_9194 ? _zz_dataOut_payload_0_8142 : _zz_dataOut_payload_0_8177);
  assign _zz_dataOut_payload_0_9196 = (_zz_dataOut_payload_0_9194 ? _zz_dataOut_payload_0_8177 : _zz_dataOut_payload_0_8142);
  assign _zz_dataOut_payload_0_9197 = (_zz_dataOut_payload_0_8143 < _zz_dataOut_payload_0_8176);
  assign _zz_dataOut_payload_0_9198 = (_zz_dataOut_payload_0_9197 ? _zz_dataOut_payload_0_8143 : _zz_dataOut_payload_0_8176);
  assign _zz_dataOut_payload_0_9199 = (_zz_dataOut_payload_0_9197 ? _zz_dataOut_payload_0_8176 : _zz_dataOut_payload_0_8143);
  assign _zz_dataOut_payload_0_9200 = (_zz_dataOut_payload_0_8144 < _zz_dataOut_payload_0_8175);
  assign _zz_dataOut_payload_0_9201 = (_zz_dataOut_payload_0_9200 ? _zz_dataOut_payload_0_8144 : _zz_dataOut_payload_0_8175);
  assign _zz_dataOut_payload_0_9202 = (_zz_dataOut_payload_0_9200 ? _zz_dataOut_payload_0_8175 : _zz_dataOut_payload_0_8144);
  assign _zz_dataOut_payload_0_9203 = (_zz_dataOut_payload_0_8145 < _zz_dataOut_payload_0_8174);
  assign _zz_dataOut_payload_0_9204 = (_zz_dataOut_payload_0_9203 ? _zz_dataOut_payload_0_8145 : _zz_dataOut_payload_0_8174);
  assign _zz_dataOut_payload_0_9205 = (_zz_dataOut_payload_0_9203 ? _zz_dataOut_payload_0_8174 : _zz_dataOut_payload_0_8145);
  assign _zz_dataOut_payload_0_9206 = (_zz_dataOut_payload_0_8146 < _zz_dataOut_payload_0_8173);
  assign _zz_dataOut_payload_0_9207 = (_zz_dataOut_payload_0_9206 ? _zz_dataOut_payload_0_8146 : _zz_dataOut_payload_0_8173);
  assign _zz_dataOut_payload_0_9208 = (_zz_dataOut_payload_0_9206 ? _zz_dataOut_payload_0_8173 : _zz_dataOut_payload_0_8146);
  assign _zz_dataOut_payload_0_9209 = (_zz_dataOut_payload_0_8147 < _zz_dataOut_payload_0_8172);
  assign _zz_dataOut_payload_0_9210 = (_zz_dataOut_payload_0_9209 ? _zz_dataOut_payload_0_8147 : _zz_dataOut_payload_0_8172);
  assign _zz_dataOut_payload_0_9211 = (_zz_dataOut_payload_0_9209 ? _zz_dataOut_payload_0_8172 : _zz_dataOut_payload_0_8147);
  assign _zz_dataOut_payload_0_9212 = (_zz_dataOut_payload_0_8148 < _zz_dataOut_payload_0_8171);
  assign _zz_dataOut_payload_0_9213 = (_zz_dataOut_payload_0_9212 ? _zz_dataOut_payload_0_8148 : _zz_dataOut_payload_0_8171);
  assign _zz_dataOut_payload_0_9214 = (_zz_dataOut_payload_0_9212 ? _zz_dataOut_payload_0_8171 : _zz_dataOut_payload_0_8148);
  assign _zz_dataOut_payload_0_9215 = (_zz_dataOut_payload_0_8149 < _zz_dataOut_payload_0_8170);
  assign _zz_dataOut_payload_0_9216 = (_zz_dataOut_payload_0_9215 ? _zz_dataOut_payload_0_8149 : _zz_dataOut_payload_0_8170);
  assign _zz_dataOut_payload_0_9217 = (_zz_dataOut_payload_0_9215 ? _zz_dataOut_payload_0_8170 : _zz_dataOut_payload_0_8149);
  assign _zz_dataOut_payload_0_9218 = (_zz_dataOut_payload_0_8150 < _zz_dataOut_payload_0_8169);
  assign _zz_dataOut_payload_0_9219 = (_zz_dataOut_payload_0_9218 ? _zz_dataOut_payload_0_8150 : _zz_dataOut_payload_0_8169);
  assign _zz_dataOut_payload_0_9220 = (_zz_dataOut_payload_0_9218 ? _zz_dataOut_payload_0_8169 : _zz_dataOut_payload_0_8150);
  assign _zz_dataOut_payload_0_9221 = (_zz_dataOut_payload_0_8151 < _zz_dataOut_payload_0_8168);
  assign _zz_dataOut_payload_0_9222 = (_zz_dataOut_payload_0_9221 ? _zz_dataOut_payload_0_8151 : _zz_dataOut_payload_0_8168);
  assign _zz_dataOut_payload_0_9223 = (_zz_dataOut_payload_0_9221 ? _zz_dataOut_payload_0_8168 : _zz_dataOut_payload_0_8151);
  assign _zz_dataOut_payload_0_9224 = (_zz_dataOut_payload_0_8152 < _zz_dataOut_payload_0_8167);
  assign _zz_dataOut_payload_0_9225 = (_zz_dataOut_payload_0_9224 ? _zz_dataOut_payload_0_8152 : _zz_dataOut_payload_0_8167);
  assign _zz_dataOut_payload_0_9226 = (_zz_dataOut_payload_0_9224 ? _zz_dataOut_payload_0_8167 : _zz_dataOut_payload_0_8152);
  assign _zz_dataOut_payload_0_9227 = (_zz_dataOut_payload_0_8153 < _zz_dataOut_payload_0_8166);
  assign _zz_dataOut_payload_0_9228 = (_zz_dataOut_payload_0_9227 ? _zz_dataOut_payload_0_8153 : _zz_dataOut_payload_0_8166);
  assign _zz_dataOut_payload_0_9229 = (_zz_dataOut_payload_0_9227 ? _zz_dataOut_payload_0_8166 : _zz_dataOut_payload_0_8153);
  assign _zz_dataOut_payload_0_9230 = (_zz_dataOut_payload_0_8154 < _zz_dataOut_payload_0_8165);
  assign _zz_dataOut_payload_0_9231 = (_zz_dataOut_payload_0_9230 ? _zz_dataOut_payload_0_8154 : _zz_dataOut_payload_0_8165);
  assign _zz_dataOut_payload_0_9232 = (_zz_dataOut_payload_0_9230 ? _zz_dataOut_payload_0_8165 : _zz_dataOut_payload_0_8154);
  assign _zz_dataOut_payload_0_9233 = (_zz_dataOut_payload_0_8155 < _zz_dataOut_payload_0_8164);
  assign _zz_dataOut_payload_0_9234 = (_zz_dataOut_payload_0_9233 ? _zz_dataOut_payload_0_8155 : _zz_dataOut_payload_0_8164);
  assign _zz_dataOut_payload_0_9235 = (_zz_dataOut_payload_0_9233 ? _zz_dataOut_payload_0_8164 : _zz_dataOut_payload_0_8155);
  assign _zz_dataOut_payload_0_9236 = (_zz_dataOut_payload_0_8156 < _zz_dataOut_payload_0_8163);
  assign _zz_dataOut_payload_0_9237 = (_zz_dataOut_payload_0_9236 ? _zz_dataOut_payload_0_8156 : _zz_dataOut_payload_0_8163);
  assign _zz_dataOut_payload_0_9238 = (_zz_dataOut_payload_0_9236 ? _zz_dataOut_payload_0_8163 : _zz_dataOut_payload_0_8156);
  assign _zz_dataOut_payload_0_9239 = (_zz_dataOut_payload_0_8157 < _zz_dataOut_payload_0_8162);
  assign _zz_dataOut_payload_0_9240 = (_zz_dataOut_payload_0_9239 ? _zz_dataOut_payload_0_8157 : _zz_dataOut_payload_0_8162);
  assign _zz_dataOut_payload_0_9241 = (_zz_dataOut_payload_0_9239 ? _zz_dataOut_payload_0_8162 : _zz_dataOut_payload_0_8157);
  assign _zz_dataOut_payload_0_9242 = (_zz_dataOut_payload_0_8158 < _zz_dataOut_payload_0_8161);
  assign _zz_dataOut_payload_0_9243 = (_zz_dataOut_payload_0_9242 ? _zz_dataOut_payload_0_8158 : _zz_dataOut_payload_0_8161);
  assign _zz_dataOut_payload_0_9244 = (_zz_dataOut_payload_0_9242 ? _zz_dataOut_payload_0_8161 : _zz_dataOut_payload_0_8158);
  assign _zz_dataOut_payload_0_9245 = (_zz_dataOut_payload_0_8159 < _zz_dataOut_payload_0_8160);
  assign _zz_dataOut_payload_0_9246 = (_zz_dataOut_payload_0_9245 ? _zz_dataOut_payload_0_8159 : _zz_dataOut_payload_0_8160);
  assign _zz_dataOut_payload_0_9247 = (_zz_dataOut_payload_0_9245 ? _zz_dataOut_payload_0_8160 : _zz_dataOut_payload_0_8159);
  assign _zz_dataOut_payload_0_9248 = (_zz_dataOut_payload_0_9153 < _zz_dataOut_payload_0_9201);
  assign _zz_dataOut_payload_0_9249 = (_zz_dataOut_payload_0_9248 ? _zz_dataOut_payload_0_9153 : _zz_dataOut_payload_0_9201);
  assign _zz_dataOut_payload_0_9250 = (_zz_dataOut_payload_0_9248 ? _zz_dataOut_payload_0_9201 : _zz_dataOut_payload_0_9153);
  assign _zz_dataOut_payload_0_9251 = (_zz_dataOut_payload_0_9156 < _zz_dataOut_payload_0_9204);
  assign _zz_dataOut_payload_0_9252 = (_zz_dataOut_payload_0_9251 ? _zz_dataOut_payload_0_9156 : _zz_dataOut_payload_0_9204);
  assign _zz_dataOut_payload_0_9253 = (_zz_dataOut_payload_0_9251 ? _zz_dataOut_payload_0_9204 : _zz_dataOut_payload_0_9156);
  assign _zz_dataOut_payload_0_9254 = (_zz_dataOut_payload_0_9159 < _zz_dataOut_payload_0_9207);
  assign _zz_dataOut_payload_0_9255 = (_zz_dataOut_payload_0_9254 ? _zz_dataOut_payload_0_9159 : _zz_dataOut_payload_0_9207);
  assign _zz_dataOut_payload_0_9256 = (_zz_dataOut_payload_0_9254 ? _zz_dataOut_payload_0_9207 : _zz_dataOut_payload_0_9159);
  assign _zz_dataOut_payload_0_9257 = (_zz_dataOut_payload_0_9162 < _zz_dataOut_payload_0_9210);
  assign _zz_dataOut_payload_0_9258 = (_zz_dataOut_payload_0_9257 ? _zz_dataOut_payload_0_9162 : _zz_dataOut_payload_0_9210);
  assign _zz_dataOut_payload_0_9259 = (_zz_dataOut_payload_0_9257 ? _zz_dataOut_payload_0_9210 : _zz_dataOut_payload_0_9162);
  assign _zz_dataOut_payload_0_9260 = (_zz_dataOut_payload_0_9165 < _zz_dataOut_payload_0_9213);
  assign _zz_dataOut_payload_0_9261 = (_zz_dataOut_payload_0_9260 ? _zz_dataOut_payload_0_9165 : _zz_dataOut_payload_0_9213);
  assign _zz_dataOut_payload_0_9262 = (_zz_dataOut_payload_0_9260 ? _zz_dataOut_payload_0_9213 : _zz_dataOut_payload_0_9165);
  assign _zz_dataOut_payload_0_9263 = (_zz_dataOut_payload_0_9168 < _zz_dataOut_payload_0_9216);
  assign _zz_dataOut_payload_0_9264 = (_zz_dataOut_payload_0_9263 ? _zz_dataOut_payload_0_9168 : _zz_dataOut_payload_0_9216);
  assign _zz_dataOut_payload_0_9265 = (_zz_dataOut_payload_0_9263 ? _zz_dataOut_payload_0_9216 : _zz_dataOut_payload_0_9168);
  assign _zz_dataOut_payload_0_9266 = (_zz_dataOut_payload_0_9171 < _zz_dataOut_payload_0_9219);
  assign _zz_dataOut_payload_0_9267 = (_zz_dataOut_payload_0_9266 ? _zz_dataOut_payload_0_9171 : _zz_dataOut_payload_0_9219);
  assign _zz_dataOut_payload_0_9268 = (_zz_dataOut_payload_0_9266 ? _zz_dataOut_payload_0_9219 : _zz_dataOut_payload_0_9171);
  assign _zz_dataOut_payload_0_9269 = (_zz_dataOut_payload_0_9174 < _zz_dataOut_payload_0_9222);
  assign _zz_dataOut_payload_0_9270 = (_zz_dataOut_payload_0_9269 ? _zz_dataOut_payload_0_9174 : _zz_dataOut_payload_0_9222);
  assign _zz_dataOut_payload_0_9271 = (_zz_dataOut_payload_0_9269 ? _zz_dataOut_payload_0_9222 : _zz_dataOut_payload_0_9174);
  assign _zz_dataOut_payload_0_9272 = (_zz_dataOut_payload_0_9177 < _zz_dataOut_payload_0_9225);
  assign _zz_dataOut_payload_0_9273 = (_zz_dataOut_payload_0_9272 ? _zz_dataOut_payload_0_9177 : _zz_dataOut_payload_0_9225);
  assign _zz_dataOut_payload_0_9274 = (_zz_dataOut_payload_0_9272 ? _zz_dataOut_payload_0_9225 : _zz_dataOut_payload_0_9177);
  assign _zz_dataOut_payload_0_9275 = (_zz_dataOut_payload_0_9180 < _zz_dataOut_payload_0_9228);
  assign _zz_dataOut_payload_0_9276 = (_zz_dataOut_payload_0_9275 ? _zz_dataOut_payload_0_9180 : _zz_dataOut_payload_0_9228);
  assign _zz_dataOut_payload_0_9277 = (_zz_dataOut_payload_0_9275 ? _zz_dataOut_payload_0_9228 : _zz_dataOut_payload_0_9180);
  assign _zz_dataOut_payload_0_9278 = (_zz_dataOut_payload_0_9183 < _zz_dataOut_payload_0_9231);
  assign _zz_dataOut_payload_0_9279 = (_zz_dataOut_payload_0_9278 ? _zz_dataOut_payload_0_9183 : _zz_dataOut_payload_0_9231);
  assign _zz_dataOut_payload_0_9280 = (_zz_dataOut_payload_0_9278 ? _zz_dataOut_payload_0_9231 : _zz_dataOut_payload_0_9183);
  assign _zz_dataOut_payload_0_9281 = (_zz_dataOut_payload_0_9186 < _zz_dataOut_payload_0_9234);
  assign _zz_dataOut_payload_0_9282 = (_zz_dataOut_payload_0_9281 ? _zz_dataOut_payload_0_9186 : _zz_dataOut_payload_0_9234);
  assign _zz_dataOut_payload_0_9283 = (_zz_dataOut_payload_0_9281 ? _zz_dataOut_payload_0_9234 : _zz_dataOut_payload_0_9186);
  assign _zz_dataOut_payload_0_9284 = (_zz_dataOut_payload_0_9189 < _zz_dataOut_payload_0_9237);
  assign _zz_dataOut_payload_0_9285 = (_zz_dataOut_payload_0_9284 ? _zz_dataOut_payload_0_9189 : _zz_dataOut_payload_0_9237);
  assign _zz_dataOut_payload_0_9286 = (_zz_dataOut_payload_0_9284 ? _zz_dataOut_payload_0_9237 : _zz_dataOut_payload_0_9189);
  assign _zz_dataOut_payload_0_9287 = (_zz_dataOut_payload_0_9192 < _zz_dataOut_payload_0_9240);
  assign _zz_dataOut_payload_0_9288 = (_zz_dataOut_payload_0_9287 ? _zz_dataOut_payload_0_9192 : _zz_dataOut_payload_0_9240);
  assign _zz_dataOut_payload_0_9289 = (_zz_dataOut_payload_0_9287 ? _zz_dataOut_payload_0_9240 : _zz_dataOut_payload_0_9192);
  assign _zz_dataOut_payload_0_9290 = (_zz_dataOut_payload_0_9195 < _zz_dataOut_payload_0_9243);
  assign _zz_dataOut_payload_0_9291 = (_zz_dataOut_payload_0_9290 ? _zz_dataOut_payload_0_9195 : _zz_dataOut_payload_0_9243);
  assign _zz_dataOut_payload_0_9292 = (_zz_dataOut_payload_0_9290 ? _zz_dataOut_payload_0_9243 : _zz_dataOut_payload_0_9195);
  assign _zz_dataOut_payload_0_9293 = (_zz_dataOut_payload_0_9198 < _zz_dataOut_payload_0_9246);
  assign _zz_dataOut_payload_0_9294 = (_zz_dataOut_payload_0_9293 ? _zz_dataOut_payload_0_9198 : _zz_dataOut_payload_0_9246);
  assign _zz_dataOut_payload_0_9295 = (_zz_dataOut_payload_0_9293 ? _zz_dataOut_payload_0_9246 : _zz_dataOut_payload_0_9198);
  assign _zz_dataOut_payload_0_9296 = (_zz_dataOut_payload_0_9249 < _zz_dataOut_payload_0_9273);
  assign _zz_dataOut_payload_0_9297 = (_zz_dataOut_payload_0_9296 ? _zz_dataOut_payload_0_9249 : _zz_dataOut_payload_0_9273);
  assign _zz_dataOut_payload_0_9298 = (_zz_dataOut_payload_0_9296 ? _zz_dataOut_payload_0_9273 : _zz_dataOut_payload_0_9249);
  assign _zz_dataOut_payload_0_9299 = (_zz_dataOut_payload_0_9252 < _zz_dataOut_payload_0_9276);
  assign _zz_dataOut_payload_0_9300 = (_zz_dataOut_payload_0_9299 ? _zz_dataOut_payload_0_9252 : _zz_dataOut_payload_0_9276);
  assign _zz_dataOut_payload_0_9301 = (_zz_dataOut_payload_0_9299 ? _zz_dataOut_payload_0_9276 : _zz_dataOut_payload_0_9252);
  assign _zz_dataOut_payload_0_9302 = (_zz_dataOut_payload_0_9255 < _zz_dataOut_payload_0_9279);
  assign _zz_dataOut_payload_0_9303 = (_zz_dataOut_payload_0_9302 ? _zz_dataOut_payload_0_9255 : _zz_dataOut_payload_0_9279);
  assign _zz_dataOut_payload_0_9304 = (_zz_dataOut_payload_0_9302 ? _zz_dataOut_payload_0_9279 : _zz_dataOut_payload_0_9255);
  assign _zz_dataOut_payload_0_9305 = (_zz_dataOut_payload_0_9258 < _zz_dataOut_payload_0_9282);
  assign _zz_dataOut_payload_0_9306 = (_zz_dataOut_payload_0_9305 ? _zz_dataOut_payload_0_9258 : _zz_dataOut_payload_0_9282);
  assign _zz_dataOut_payload_0_9307 = (_zz_dataOut_payload_0_9305 ? _zz_dataOut_payload_0_9282 : _zz_dataOut_payload_0_9258);
  assign _zz_dataOut_payload_0_9308 = (_zz_dataOut_payload_0_9261 < _zz_dataOut_payload_0_9285);
  assign _zz_dataOut_payload_0_9309 = (_zz_dataOut_payload_0_9308 ? _zz_dataOut_payload_0_9261 : _zz_dataOut_payload_0_9285);
  assign _zz_dataOut_payload_0_9310 = (_zz_dataOut_payload_0_9308 ? _zz_dataOut_payload_0_9285 : _zz_dataOut_payload_0_9261);
  assign _zz_dataOut_payload_0_9311 = (_zz_dataOut_payload_0_9264 < _zz_dataOut_payload_0_9288);
  assign _zz_dataOut_payload_0_9312 = (_zz_dataOut_payload_0_9311 ? _zz_dataOut_payload_0_9264 : _zz_dataOut_payload_0_9288);
  assign _zz_dataOut_payload_0_9313 = (_zz_dataOut_payload_0_9311 ? _zz_dataOut_payload_0_9288 : _zz_dataOut_payload_0_9264);
  assign _zz_dataOut_payload_0_9314 = (_zz_dataOut_payload_0_9267 < _zz_dataOut_payload_0_9291);
  assign _zz_dataOut_payload_0_9315 = (_zz_dataOut_payload_0_9314 ? _zz_dataOut_payload_0_9267 : _zz_dataOut_payload_0_9291);
  assign _zz_dataOut_payload_0_9316 = (_zz_dataOut_payload_0_9314 ? _zz_dataOut_payload_0_9291 : _zz_dataOut_payload_0_9267);
  assign _zz_dataOut_payload_0_9317 = (_zz_dataOut_payload_0_9270 < _zz_dataOut_payload_0_9294);
  assign _zz_dataOut_payload_0_9318 = (_zz_dataOut_payload_0_9317 ? _zz_dataOut_payload_0_9270 : _zz_dataOut_payload_0_9294);
  assign _zz_dataOut_payload_0_9319 = (_zz_dataOut_payload_0_9317 ? _zz_dataOut_payload_0_9294 : _zz_dataOut_payload_0_9270);
  assign _zz_dataOut_payload_0_9320 = (_zz_dataOut_payload_0_9297 < _zz_dataOut_payload_0_9309);
  assign _zz_dataOut_payload_0_9321 = (_zz_dataOut_payload_0_9320 ? _zz_dataOut_payload_0_9297 : _zz_dataOut_payload_0_9309);
  assign _zz_dataOut_payload_0_9322 = (_zz_dataOut_payload_0_9320 ? _zz_dataOut_payload_0_9309 : _zz_dataOut_payload_0_9297);
  assign _zz_dataOut_payload_0_9323 = (_zz_dataOut_payload_0_9300 < _zz_dataOut_payload_0_9312);
  assign _zz_dataOut_payload_0_9324 = (_zz_dataOut_payload_0_9323 ? _zz_dataOut_payload_0_9300 : _zz_dataOut_payload_0_9312);
  assign _zz_dataOut_payload_0_9325 = (_zz_dataOut_payload_0_9323 ? _zz_dataOut_payload_0_9312 : _zz_dataOut_payload_0_9300);
  assign _zz_dataOut_payload_0_9326 = (_zz_dataOut_payload_0_9303 < _zz_dataOut_payload_0_9315);
  assign _zz_dataOut_payload_0_9327 = (_zz_dataOut_payload_0_9326 ? _zz_dataOut_payload_0_9303 : _zz_dataOut_payload_0_9315);
  assign _zz_dataOut_payload_0_9328 = (_zz_dataOut_payload_0_9326 ? _zz_dataOut_payload_0_9315 : _zz_dataOut_payload_0_9303);
  assign _zz_dataOut_payload_0_9329 = (_zz_dataOut_payload_0_9306 < _zz_dataOut_payload_0_9318);
  assign _zz_dataOut_payload_0_9330 = (_zz_dataOut_payload_0_9329 ? _zz_dataOut_payload_0_9306 : _zz_dataOut_payload_0_9318);
  assign _zz_dataOut_payload_0_9331 = (_zz_dataOut_payload_0_9329 ? _zz_dataOut_payload_0_9318 : _zz_dataOut_payload_0_9306);
  assign _zz_dataOut_payload_0_9332 = (_zz_dataOut_payload_0_9321 < _zz_dataOut_payload_0_9327);
  assign _zz_dataOut_payload_0_9333 = (_zz_dataOut_payload_0_9332 ? _zz_dataOut_payload_0_9321 : _zz_dataOut_payload_0_9327);
  assign _zz_dataOut_payload_0_9334 = (_zz_dataOut_payload_0_9332 ? _zz_dataOut_payload_0_9327 : _zz_dataOut_payload_0_9321);
  assign _zz_dataOut_payload_0_9335 = (_zz_dataOut_payload_0_9324 < _zz_dataOut_payload_0_9330);
  assign _zz_dataOut_payload_0_9336 = (_zz_dataOut_payload_0_9335 ? _zz_dataOut_payload_0_9324 : _zz_dataOut_payload_0_9330);
  assign _zz_dataOut_payload_0_9337 = (_zz_dataOut_payload_0_9335 ? _zz_dataOut_payload_0_9330 : _zz_dataOut_payload_0_9324);
  assign _zz_dataOut_payload_0_9338 = (_zz_dataOut_payload_0_9333 < _zz_dataOut_payload_0_9336);
  assign _zz_dataOut_payload_0_9339 = (_zz_dataOut_payload_0_9334 < _zz_dataOut_payload_0_9337);
  assign _zz_dataOut_payload_0_9344 = (_zz_dataOut_payload_0_9322 < _zz_dataOut_payload_0_9328);
  assign _zz_dataOut_payload_0_9345 = (_zz_dataOut_payload_0_9344 ? _zz_dataOut_payload_0_9322 : _zz_dataOut_payload_0_9328);
  assign _zz_dataOut_payload_0_9346 = (_zz_dataOut_payload_0_9344 ? _zz_dataOut_payload_0_9328 : _zz_dataOut_payload_0_9322);
  assign _zz_dataOut_payload_0_9347 = (_zz_dataOut_payload_0_9325 < _zz_dataOut_payload_0_9331);
  assign _zz_dataOut_payload_0_9348 = (_zz_dataOut_payload_0_9347 ? _zz_dataOut_payload_0_9325 : _zz_dataOut_payload_0_9331);
  assign _zz_dataOut_payload_0_9349 = (_zz_dataOut_payload_0_9347 ? _zz_dataOut_payload_0_9331 : _zz_dataOut_payload_0_9325);
  assign _zz_dataOut_payload_0_9350 = (_zz_dataOut_payload_0_9345 < _zz_dataOut_payload_0_9348);
  assign _zz_dataOut_payload_0_9351 = (_zz_dataOut_payload_0_9346 < _zz_dataOut_payload_0_9349);
  assign _zz_dataOut_payload_0_9364 = (_zz_dataOut_payload_0_9298 < _zz_dataOut_payload_0_9310);
  assign _zz_dataOut_payload_0_9365 = (_zz_dataOut_payload_0_9364 ? _zz_dataOut_payload_0_9298 : _zz_dataOut_payload_0_9310);
  assign _zz_dataOut_payload_0_9366 = (_zz_dataOut_payload_0_9364 ? _zz_dataOut_payload_0_9310 : _zz_dataOut_payload_0_9298);
  assign _zz_dataOut_payload_0_9367 = (_zz_dataOut_payload_0_9301 < _zz_dataOut_payload_0_9313);
  assign _zz_dataOut_payload_0_9368 = (_zz_dataOut_payload_0_9367 ? _zz_dataOut_payload_0_9301 : _zz_dataOut_payload_0_9313);
  assign _zz_dataOut_payload_0_9369 = (_zz_dataOut_payload_0_9367 ? _zz_dataOut_payload_0_9313 : _zz_dataOut_payload_0_9301);
  assign _zz_dataOut_payload_0_9370 = (_zz_dataOut_payload_0_9304 < _zz_dataOut_payload_0_9316);
  assign _zz_dataOut_payload_0_9371 = (_zz_dataOut_payload_0_9370 ? _zz_dataOut_payload_0_9304 : _zz_dataOut_payload_0_9316);
  assign _zz_dataOut_payload_0_9372 = (_zz_dataOut_payload_0_9370 ? _zz_dataOut_payload_0_9316 : _zz_dataOut_payload_0_9304);
  assign _zz_dataOut_payload_0_9373 = (_zz_dataOut_payload_0_9307 < _zz_dataOut_payload_0_9319);
  assign _zz_dataOut_payload_0_9374 = (_zz_dataOut_payload_0_9373 ? _zz_dataOut_payload_0_9307 : _zz_dataOut_payload_0_9319);
  assign _zz_dataOut_payload_0_9375 = (_zz_dataOut_payload_0_9373 ? _zz_dataOut_payload_0_9319 : _zz_dataOut_payload_0_9307);
  assign _zz_dataOut_payload_0_9376 = (_zz_dataOut_payload_0_9365 < _zz_dataOut_payload_0_9371);
  assign _zz_dataOut_payload_0_9377 = (_zz_dataOut_payload_0_9376 ? _zz_dataOut_payload_0_9365 : _zz_dataOut_payload_0_9371);
  assign _zz_dataOut_payload_0_9378 = (_zz_dataOut_payload_0_9376 ? _zz_dataOut_payload_0_9371 : _zz_dataOut_payload_0_9365);
  assign _zz_dataOut_payload_0_9379 = (_zz_dataOut_payload_0_9368 < _zz_dataOut_payload_0_9374);
  assign _zz_dataOut_payload_0_9380 = (_zz_dataOut_payload_0_9379 ? _zz_dataOut_payload_0_9368 : _zz_dataOut_payload_0_9374);
  assign _zz_dataOut_payload_0_9381 = (_zz_dataOut_payload_0_9379 ? _zz_dataOut_payload_0_9374 : _zz_dataOut_payload_0_9368);
  assign _zz_dataOut_payload_0_9382 = (_zz_dataOut_payload_0_9377 < _zz_dataOut_payload_0_9380);
  assign _zz_dataOut_payload_0_9383 = (_zz_dataOut_payload_0_9378 < _zz_dataOut_payload_0_9381);
  assign _zz_dataOut_payload_0_9388 = (_zz_dataOut_payload_0_9366 < _zz_dataOut_payload_0_9372);
  assign _zz_dataOut_payload_0_9389 = (_zz_dataOut_payload_0_9388 ? _zz_dataOut_payload_0_9366 : _zz_dataOut_payload_0_9372);
  assign _zz_dataOut_payload_0_9390 = (_zz_dataOut_payload_0_9388 ? _zz_dataOut_payload_0_9372 : _zz_dataOut_payload_0_9366);
  assign _zz_dataOut_payload_0_9391 = (_zz_dataOut_payload_0_9369 < _zz_dataOut_payload_0_9375);
  assign _zz_dataOut_payload_0_9392 = (_zz_dataOut_payload_0_9391 ? _zz_dataOut_payload_0_9369 : _zz_dataOut_payload_0_9375);
  assign _zz_dataOut_payload_0_9393 = (_zz_dataOut_payload_0_9391 ? _zz_dataOut_payload_0_9375 : _zz_dataOut_payload_0_9369);
  assign _zz_dataOut_payload_0_9394 = (_zz_dataOut_payload_0_9389 < _zz_dataOut_payload_0_9392);
  assign _zz_dataOut_payload_0_9395 = (_zz_dataOut_payload_0_9390 < _zz_dataOut_payload_0_9393);
  assign _zz_dataOut_payload_0_9424 = (_zz_dataOut_payload_0_9250 < _zz_dataOut_payload_0_9274);
  assign _zz_dataOut_payload_0_9425 = (_zz_dataOut_payload_0_9424 ? _zz_dataOut_payload_0_9250 : _zz_dataOut_payload_0_9274);
  assign _zz_dataOut_payload_0_9426 = (_zz_dataOut_payload_0_9424 ? _zz_dataOut_payload_0_9274 : _zz_dataOut_payload_0_9250);
  assign _zz_dataOut_payload_0_9427 = (_zz_dataOut_payload_0_9253 < _zz_dataOut_payload_0_9277);
  assign _zz_dataOut_payload_0_9428 = (_zz_dataOut_payload_0_9427 ? _zz_dataOut_payload_0_9253 : _zz_dataOut_payload_0_9277);
  assign _zz_dataOut_payload_0_9429 = (_zz_dataOut_payload_0_9427 ? _zz_dataOut_payload_0_9277 : _zz_dataOut_payload_0_9253);
  assign _zz_dataOut_payload_0_9430 = (_zz_dataOut_payload_0_9256 < _zz_dataOut_payload_0_9280);
  assign _zz_dataOut_payload_0_9431 = (_zz_dataOut_payload_0_9430 ? _zz_dataOut_payload_0_9256 : _zz_dataOut_payload_0_9280);
  assign _zz_dataOut_payload_0_9432 = (_zz_dataOut_payload_0_9430 ? _zz_dataOut_payload_0_9280 : _zz_dataOut_payload_0_9256);
  assign _zz_dataOut_payload_0_9433 = (_zz_dataOut_payload_0_9259 < _zz_dataOut_payload_0_9283);
  assign _zz_dataOut_payload_0_9434 = (_zz_dataOut_payload_0_9433 ? _zz_dataOut_payload_0_9259 : _zz_dataOut_payload_0_9283);
  assign _zz_dataOut_payload_0_9435 = (_zz_dataOut_payload_0_9433 ? _zz_dataOut_payload_0_9283 : _zz_dataOut_payload_0_9259);
  assign _zz_dataOut_payload_0_9436 = (_zz_dataOut_payload_0_9262 < _zz_dataOut_payload_0_9286);
  assign _zz_dataOut_payload_0_9437 = (_zz_dataOut_payload_0_9436 ? _zz_dataOut_payload_0_9262 : _zz_dataOut_payload_0_9286);
  assign _zz_dataOut_payload_0_9438 = (_zz_dataOut_payload_0_9436 ? _zz_dataOut_payload_0_9286 : _zz_dataOut_payload_0_9262);
  assign _zz_dataOut_payload_0_9439 = (_zz_dataOut_payload_0_9265 < _zz_dataOut_payload_0_9289);
  assign _zz_dataOut_payload_0_9440 = (_zz_dataOut_payload_0_9439 ? _zz_dataOut_payload_0_9265 : _zz_dataOut_payload_0_9289);
  assign _zz_dataOut_payload_0_9441 = (_zz_dataOut_payload_0_9439 ? _zz_dataOut_payload_0_9289 : _zz_dataOut_payload_0_9265);
  assign _zz_dataOut_payload_0_9442 = (_zz_dataOut_payload_0_9268 < _zz_dataOut_payload_0_9292);
  assign _zz_dataOut_payload_0_9443 = (_zz_dataOut_payload_0_9442 ? _zz_dataOut_payload_0_9268 : _zz_dataOut_payload_0_9292);
  assign _zz_dataOut_payload_0_9444 = (_zz_dataOut_payload_0_9442 ? _zz_dataOut_payload_0_9292 : _zz_dataOut_payload_0_9268);
  assign _zz_dataOut_payload_0_9445 = (_zz_dataOut_payload_0_9271 < _zz_dataOut_payload_0_9295);
  assign _zz_dataOut_payload_0_9446 = (_zz_dataOut_payload_0_9445 ? _zz_dataOut_payload_0_9271 : _zz_dataOut_payload_0_9295);
  assign _zz_dataOut_payload_0_9447 = (_zz_dataOut_payload_0_9445 ? _zz_dataOut_payload_0_9295 : _zz_dataOut_payload_0_9271);
  assign _zz_dataOut_payload_0_9448 = (_zz_dataOut_payload_0_9425 < _zz_dataOut_payload_0_9437);
  assign _zz_dataOut_payload_0_9449 = (_zz_dataOut_payload_0_9448 ? _zz_dataOut_payload_0_9425 : _zz_dataOut_payload_0_9437);
  assign _zz_dataOut_payload_0_9450 = (_zz_dataOut_payload_0_9448 ? _zz_dataOut_payload_0_9437 : _zz_dataOut_payload_0_9425);
  assign _zz_dataOut_payload_0_9451 = (_zz_dataOut_payload_0_9428 < _zz_dataOut_payload_0_9440);
  assign _zz_dataOut_payload_0_9452 = (_zz_dataOut_payload_0_9451 ? _zz_dataOut_payload_0_9428 : _zz_dataOut_payload_0_9440);
  assign _zz_dataOut_payload_0_9453 = (_zz_dataOut_payload_0_9451 ? _zz_dataOut_payload_0_9440 : _zz_dataOut_payload_0_9428);
  assign _zz_dataOut_payload_0_9454 = (_zz_dataOut_payload_0_9431 < _zz_dataOut_payload_0_9443);
  assign _zz_dataOut_payload_0_9455 = (_zz_dataOut_payload_0_9454 ? _zz_dataOut_payload_0_9431 : _zz_dataOut_payload_0_9443);
  assign _zz_dataOut_payload_0_9456 = (_zz_dataOut_payload_0_9454 ? _zz_dataOut_payload_0_9443 : _zz_dataOut_payload_0_9431);
  assign _zz_dataOut_payload_0_9457 = (_zz_dataOut_payload_0_9434 < _zz_dataOut_payload_0_9446);
  assign _zz_dataOut_payload_0_9458 = (_zz_dataOut_payload_0_9457 ? _zz_dataOut_payload_0_9434 : _zz_dataOut_payload_0_9446);
  assign _zz_dataOut_payload_0_9459 = (_zz_dataOut_payload_0_9457 ? _zz_dataOut_payload_0_9446 : _zz_dataOut_payload_0_9434);
  assign _zz_dataOut_payload_0_9460 = (_zz_dataOut_payload_0_9449 < _zz_dataOut_payload_0_9455);
  assign _zz_dataOut_payload_0_9461 = (_zz_dataOut_payload_0_9460 ? _zz_dataOut_payload_0_9449 : _zz_dataOut_payload_0_9455);
  assign _zz_dataOut_payload_0_9462 = (_zz_dataOut_payload_0_9460 ? _zz_dataOut_payload_0_9455 : _zz_dataOut_payload_0_9449);
  assign _zz_dataOut_payload_0_9463 = (_zz_dataOut_payload_0_9452 < _zz_dataOut_payload_0_9458);
  assign _zz_dataOut_payload_0_9464 = (_zz_dataOut_payload_0_9463 ? _zz_dataOut_payload_0_9452 : _zz_dataOut_payload_0_9458);
  assign _zz_dataOut_payload_0_9465 = (_zz_dataOut_payload_0_9463 ? _zz_dataOut_payload_0_9458 : _zz_dataOut_payload_0_9452);
  assign _zz_dataOut_payload_0_9466 = (_zz_dataOut_payload_0_9461 < _zz_dataOut_payload_0_9464);
  assign _zz_dataOut_payload_0_9467 = (_zz_dataOut_payload_0_9462 < _zz_dataOut_payload_0_9465);
  assign _zz_dataOut_payload_0_9472 = (_zz_dataOut_payload_0_9450 < _zz_dataOut_payload_0_9456);
  assign _zz_dataOut_payload_0_9473 = (_zz_dataOut_payload_0_9472 ? _zz_dataOut_payload_0_9450 : _zz_dataOut_payload_0_9456);
  assign _zz_dataOut_payload_0_9474 = (_zz_dataOut_payload_0_9472 ? _zz_dataOut_payload_0_9456 : _zz_dataOut_payload_0_9450);
  assign _zz_dataOut_payload_0_9475 = (_zz_dataOut_payload_0_9453 < _zz_dataOut_payload_0_9459);
  assign _zz_dataOut_payload_0_9476 = (_zz_dataOut_payload_0_9475 ? _zz_dataOut_payload_0_9453 : _zz_dataOut_payload_0_9459);
  assign _zz_dataOut_payload_0_9477 = (_zz_dataOut_payload_0_9475 ? _zz_dataOut_payload_0_9459 : _zz_dataOut_payload_0_9453);
  assign _zz_dataOut_payload_0_9478 = (_zz_dataOut_payload_0_9473 < _zz_dataOut_payload_0_9476);
  assign _zz_dataOut_payload_0_9479 = (_zz_dataOut_payload_0_9474 < _zz_dataOut_payload_0_9477);
  assign _zz_dataOut_payload_0_9492 = (_zz_dataOut_payload_0_9426 < _zz_dataOut_payload_0_9438);
  assign _zz_dataOut_payload_0_9493 = (_zz_dataOut_payload_0_9492 ? _zz_dataOut_payload_0_9426 : _zz_dataOut_payload_0_9438);
  assign _zz_dataOut_payload_0_9494 = (_zz_dataOut_payload_0_9492 ? _zz_dataOut_payload_0_9438 : _zz_dataOut_payload_0_9426);
  assign _zz_dataOut_payload_0_9495 = (_zz_dataOut_payload_0_9429 < _zz_dataOut_payload_0_9441);
  assign _zz_dataOut_payload_0_9496 = (_zz_dataOut_payload_0_9495 ? _zz_dataOut_payload_0_9429 : _zz_dataOut_payload_0_9441);
  assign _zz_dataOut_payload_0_9497 = (_zz_dataOut_payload_0_9495 ? _zz_dataOut_payload_0_9441 : _zz_dataOut_payload_0_9429);
  assign _zz_dataOut_payload_0_9498 = (_zz_dataOut_payload_0_9432 < _zz_dataOut_payload_0_9444);
  assign _zz_dataOut_payload_0_9499 = (_zz_dataOut_payload_0_9498 ? _zz_dataOut_payload_0_9432 : _zz_dataOut_payload_0_9444);
  assign _zz_dataOut_payload_0_9500 = (_zz_dataOut_payload_0_9498 ? _zz_dataOut_payload_0_9444 : _zz_dataOut_payload_0_9432);
  assign _zz_dataOut_payload_0_9501 = (_zz_dataOut_payload_0_9435 < _zz_dataOut_payload_0_9447);
  assign _zz_dataOut_payload_0_9502 = (_zz_dataOut_payload_0_9501 ? _zz_dataOut_payload_0_9435 : _zz_dataOut_payload_0_9447);
  assign _zz_dataOut_payload_0_9503 = (_zz_dataOut_payload_0_9501 ? _zz_dataOut_payload_0_9447 : _zz_dataOut_payload_0_9435);
  assign _zz_dataOut_payload_0_9504 = (_zz_dataOut_payload_0_9493 < _zz_dataOut_payload_0_9499);
  assign _zz_dataOut_payload_0_9505 = (_zz_dataOut_payload_0_9504 ? _zz_dataOut_payload_0_9493 : _zz_dataOut_payload_0_9499);
  assign _zz_dataOut_payload_0_9506 = (_zz_dataOut_payload_0_9504 ? _zz_dataOut_payload_0_9499 : _zz_dataOut_payload_0_9493);
  assign _zz_dataOut_payload_0_9507 = (_zz_dataOut_payload_0_9496 < _zz_dataOut_payload_0_9502);
  assign _zz_dataOut_payload_0_9508 = (_zz_dataOut_payload_0_9507 ? _zz_dataOut_payload_0_9496 : _zz_dataOut_payload_0_9502);
  assign _zz_dataOut_payload_0_9509 = (_zz_dataOut_payload_0_9507 ? _zz_dataOut_payload_0_9502 : _zz_dataOut_payload_0_9496);
  assign _zz_dataOut_payload_0_9510 = (_zz_dataOut_payload_0_9505 < _zz_dataOut_payload_0_9508);
  assign _zz_dataOut_payload_0_9511 = (_zz_dataOut_payload_0_9506 < _zz_dataOut_payload_0_9509);
  assign _zz_dataOut_payload_0_9516 = (_zz_dataOut_payload_0_9494 < _zz_dataOut_payload_0_9500);
  assign _zz_dataOut_payload_0_9517 = (_zz_dataOut_payload_0_9516 ? _zz_dataOut_payload_0_9494 : _zz_dataOut_payload_0_9500);
  assign _zz_dataOut_payload_0_9518 = (_zz_dataOut_payload_0_9516 ? _zz_dataOut_payload_0_9500 : _zz_dataOut_payload_0_9494);
  assign _zz_dataOut_payload_0_9519 = (_zz_dataOut_payload_0_9497 < _zz_dataOut_payload_0_9503);
  assign _zz_dataOut_payload_0_9520 = (_zz_dataOut_payload_0_9519 ? _zz_dataOut_payload_0_9497 : _zz_dataOut_payload_0_9503);
  assign _zz_dataOut_payload_0_9521 = (_zz_dataOut_payload_0_9519 ? _zz_dataOut_payload_0_9503 : _zz_dataOut_payload_0_9497);
  assign _zz_dataOut_payload_0_9522 = (_zz_dataOut_payload_0_9517 < _zz_dataOut_payload_0_9520);
  assign _zz_dataOut_payload_0_9523 = (_zz_dataOut_payload_0_9518 < _zz_dataOut_payload_0_9521);
  assign _zz_dataOut_payload_0_9584 = (_zz_dataOut_payload_0_9247 < _zz_dataOut_payload_0_9199);
  assign _zz_dataOut_payload_0_9585 = (_zz_dataOut_payload_0_9584 ? _zz_dataOut_payload_0_9247 : _zz_dataOut_payload_0_9199);
  assign _zz_dataOut_payload_0_9586 = (_zz_dataOut_payload_0_9584 ? _zz_dataOut_payload_0_9199 : _zz_dataOut_payload_0_9247);
  assign _zz_dataOut_payload_0_9587 = (_zz_dataOut_payload_0_9244 < _zz_dataOut_payload_0_9196);
  assign _zz_dataOut_payload_0_9588 = (_zz_dataOut_payload_0_9587 ? _zz_dataOut_payload_0_9244 : _zz_dataOut_payload_0_9196);
  assign _zz_dataOut_payload_0_9589 = (_zz_dataOut_payload_0_9587 ? _zz_dataOut_payload_0_9196 : _zz_dataOut_payload_0_9244);
  assign _zz_dataOut_payload_0_9590 = (_zz_dataOut_payload_0_9241 < _zz_dataOut_payload_0_9193);
  assign _zz_dataOut_payload_0_9591 = (_zz_dataOut_payload_0_9590 ? _zz_dataOut_payload_0_9241 : _zz_dataOut_payload_0_9193);
  assign _zz_dataOut_payload_0_9592 = (_zz_dataOut_payload_0_9590 ? _zz_dataOut_payload_0_9193 : _zz_dataOut_payload_0_9241);
  assign _zz_dataOut_payload_0_9593 = (_zz_dataOut_payload_0_9238 < _zz_dataOut_payload_0_9190);
  assign _zz_dataOut_payload_0_9594 = (_zz_dataOut_payload_0_9593 ? _zz_dataOut_payload_0_9238 : _zz_dataOut_payload_0_9190);
  assign _zz_dataOut_payload_0_9595 = (_zz_dataOut_payload_0_9593 ? _zz_dataOut_payload_0_9190 : _zz_dataOut_payload_0_9238);
  assign _zz_dataOut_payload_0_9596 = (_zz_dataOut_payload_0_9235 < _zz_dataOut_payload_0_9187);
  assign _zz_dataOut_payload_0_9597 = (_zz_dataOut_payload_0_9596 ? _zz_dataOut_payload_0_9235 : _zz_dataOut_payload_0_9187);
  assign _zz_dataOut_payload_0_9598 = (_zz_dataOut_payload_0_9596 ? _zz_dataOut_payload_0_9187 : _zz_dataOut_payload_0_9235);
  assign _zz_dataOut_payload_0_9599 = (_zz_dataOut_payload_0_9232 < _zz_dataOut_payload_0_9184);
  assign _zz_dataOut_payload_0_9600 = (_zz_dataOut_payload_0_9599 ? _zz_dataOut_payload_0_9232 : _zz_dataOut_payload_0_9184);
  assign _zz_dataOut_payload_0_9601 = (_zz_dataOut_payload_0_9599 ? _zz_dataOut_payload_0_9184 : _zz_dataOut_payload_0_9232);
  assign _zz_dataOut_payload_0_9602 = (_zz_dataOut_payload_0_9229 < _zz_dataOut_payload_0_9181);
  assign _zz_dataOut_payload_0_9603 = (_zz_dataOut_payload_0_9602 ? _zz_dataOut_payload_0_9229 : _zz_dataOut_payload_0_9181);
  assign _zz_dataOut_payload_0_9604 = (_zz_dataOut_payload_0_9602 ? _zz_dataOut_payload_0_9181 : _zz_dataOut_payload_0_9229);
  assign _zz_dataOut_payload_0_9605 = (_zz_dataOut_payload_0_9226 < _zz_dataOut_payload_0_9178);
  assign _zz_dataOut_payload_0_9606 = (_zz_dataOut_payload_0_9605 ? _zz_dataOut_payload_0_9226 : _zz_dataOut_payload_0_9178);
  assign _zz_dataOut_payload_0_9607 = (_zz_dataOut_payload_0_9605 ? _zz_dataOut_payload_0_9178 : _zz_dataOut_payload_0_9226);
  assign _zz_dataOut_payload_0_9608 = (_zz_dataOut_payload_0_9223 < _zz_dataOut_payload_0_9175);
  assign _zz_dataOut_payload_0_9609 = (_zz_dataOut_payload_0_9608 ? _zz_dataOut_payload_0_9223 : _zz_dataOut_payload_0_9175);
  assign _zz_dataOut_payload_0_9610 = (_zz_dataOut_payload_0_9608 ? _zz_dataOut_payload_0_9175 : _zz_dataOut_payload_0_9223);
  assign _zz_dataOut_payload_0_9611 = (_zz_dataOut_payload_0_9220 < _zz_dataOut_payload_0_9172);
  assign _zz_dataOut_payload_0_9612 = (_zz_dataOut_payload_0_9611 ? _zz_dataOut_payload_0_9220 : _zz_dataOut_payload_0_9172);
  assign _zz_dataOut_payload_0_9613 = (_zz_dataOut_payload_0_9611 ? _zz_dataOut_payload_0_9172 : _zz_dataOut_payload_0_9220);
  assign _zz_dataOut_payload_0_9614 = (_zz_dataOut_payload_0_9217 < _zz_dataOut_payload_0_9169);
  assign _zz_dataOut_payload_0_9615 = (_zz_dataOut_payload_0_9614 ? _zz_dataOut_payload_0_9217 : _zz_dataOut_payload_0_9169);
  assign _zz_dataOut_payload_0_9616 = (_zz_dataOut_payload_0_9614 ? _zz_dataOut_payload_0_9169 : _zz_dataOut_payload_0_9217);
  assign _zz_dataOut_payload_0_9617 = (_zz_dataOut_payload_0_9214 < _zz_dataOut_payload_0_9166);
  assign _zz_dataOut_payload_0_9618 = (_zz_dataOut_payload_0_9617 ? _zz_dataOut_payload_0_9214 : _zz_dataOut_payload_0_9166);
  assign _zz_dataOut_payload_0_9619 = (_zz_dataOut_payload_0_9617 ? _zz_dataOut_payload_0_9166 : _zz_dataOut_payload_0_9214);
  assign _zz_dataOut_payload_0_9620 = (_zz_dataOut_payload_0_9211 < _zz_dataOut_payload_0_9163);
  assign _zz_dataOut_payload_0_9621 = (_zz_dataOut_payload_0_9620 ? _zz_dataOut_payload_0_9211 : _zz_dataOut_payload_0_9163);
  assign _zz_dataOut_payload_0_9622 = (_zz_dataOut_payload_0_9620 ? _zz_dataOut_payload_0_9163 : _zz_dataOut_payload_0_9211);
  assign _zz_dataOut_payload_0_9623 = (_zz_dataOut_payload_0_9208 < _zz_dataOut_payload_0_9160);
  assign _zz_dataOut_payload_0_9624 = (_zz_dataOut_payload_0_9623 ? _zz_dataOut_payload_0_9208 : _zz_dataOut_payload_0_9160);
  assign _zz_dataOut_payload_0_9625 = (_zz_dataOut_payload_0_9623 ? _zz_dataOut_payload_0_9160 : _zz_dataOut_payload_0_9208);
  assign _zz_dataOut_payload_0_9626 = (_zz_dataOut_payload_0_9205 < _zz_dataOut_payload_0_9157);
  assign _zz_dataOut_payload_0_9627 = (_zz_dataOut_payload_0_9626 ? _zz_dataOut_payload_0_9205 : _zz_dataOut_payload_0_9157);
  assign _zz_dataOut_payload_0_9628 = (_zz_dataOut_payload_0_9626 ? _zz_dataOut_payload_0_9157 : _zz_dataOut_payload_0_9205);
  assign _zz_dataOut_payload_0_9629 = (_zz_dataOut_payload_0_9202 < _zz_dataOut_payload_0_9154);
  assign _zz_dataOut_payload_0_9630 = (_zz_dataOut_payload_0_9629 ? _zz_dataOut_payload_0_9202 : _zz_dataOut_payload_0_9154);
  assign _zz_dataOut_payload_0_9631 = (_zz_dataOut_payload_0_9629 ? _zz_dataOut_payload_0_9154 : _zz_dataOut_payload_0_9202);
  assign _zz_dataOut_payload_0_9632 = (_zz_dataOut_payload_0_9585 < _zz_dataOut_payload_0_9609);
  assign _zz_dataOut_payload_0_9633 = (_zz_dataOut_payload_0_9632 ? _zz_dataOut_payload_0_9585 : _zz_dataOut_payload_0_9609);
  assign _zz_dataOut_payload_0_9634 = (_zz_dataOut_payload_0_9632 ? _zz_dataOut_payload_0_9609 : _zz_dataOut_payload_0_9585);
  assign _zz_dataOut_payload_0_9635 = (_zz_dataOut_payload_0_9588 < _zz_dataOut_payload_0_9612);
  assign _zz_dataOut_payload_0_9636 = (_zz_dataOut_payload_0_9635 ? _zz_dataOut_payload_0_9588 : _zz_dataOut_payload_0_9612);
  assign _zz_dataOut_payload_0_9637 = (_zz_dataOut_payload_0_9635 ? _zz_dataOut_payload_0_9612 : _zz_dataOut_payload_0_9588);
  assign _zz_dataOut_payload_0_9638 = (_zz_dataOut_payload_0_9591 < _zz_dataOut_payload_0_9615);
  assign _zz_dataOut_payload_0_9639 = (_zz_dataOut_payload_0_9638 ? _zz_dataOut_payload_0_9591 : _zz_dataOut_payload_0_9615);
  assign _zz_dataOut_payload_0_9640 = (_zz_dataOut_payload_0_9638 ? _zz_dataOut_payload_0_9615 : _zz_dataOut_payload_0_9591);
  assign _zz_dataOut_payload_0_9641 = (_zz_dataOut_payload_0_9594 < _zz_dataOut_payload_0_9618);
  assign _zz_dataOut_payload_0_9642 = (_zz_dataOut_payload_0_9641 ? _zz_dataOut_payload_0_9594 : _zz_dataOut_payload_0_9618);
  assign _zz_dataOut_payload_0_9643 = (_zz_dataOut_payload_0_9641 ? _zz_dataOut_payload_0_9618 : _zz_dataOut_payload_0_9594);
  assign _zz_dataOut_payload_0_9644 = (_zz_dataOut_payload_0_9597 < _zz_dataOut_payload_0_9621);
  assign _zz_dataOut_payload_0_9645 = (_zz_dataOut_payload_0_9644 ? _zz_dataOut_payload_0_9597 : _zz_dataOut_payload_0_9621);
  assign _zz_dataOut_payload_0_9646 = (_zz_dataOut_payload_0_9644 ? _zz_dataOut_payload_0_9621 : _zz_dataOut_payload_0_9597);
  assign _zz_dataOut_payload_0_9647 = (_zz_dataOut_payload_0_9600 < _zz_dataOut_payload_0_9624);
  assign _zz_dataOut_payload_0_9648 = (_zz_dataOut_payload_0_9647 ? _zz_dataOut_payload_0_9600 : _zz_dataOut_payload_0_9624);
  assign _zz_dataOut_payload_0_9649 = (_zz_dataOut_payload_0_9647 ? _zz_dataOut_payload_0_9624 : _zz_dataOut_payload_0_9600);
  assign _zz_dataOut_payload_0_9650 = (_zz_dataOut_payload_0_9603 < _zz_dataOut_payload_0_9627);
  assign _zz_dataOut_payload_0_9651 = (_zz_dataOut_payload_0_9650 ? _zz_dataOut_payload_0_9603 : _zz_dataOut_payload_0_9627);
  assign _zz_dataOut_payload_0_9652 = (_zz_dataOut_payload_0_9650 ? _zz_dataOut_payload_0_9627 : _zz_dataOut_payload_0_9603);
  assign _zz_dataOut_payload_0_9653 = (_zz_dataOut_payload_0_9606 < _zz_dataOut_payload_0_9630);
  assign _zz_dataOut_payload_0_9654 = (_zz_dataOut_payload_0_9653 ? _zz_dataOut_payload_0_9606 : _zz_dataOut_payload_0_9630);
  assign _zz_dataOut_payload_0_9655 = (_zz_dataOut_payload_0_9653 ? _zz_dataOut_payload_0_9630 : _zz_dataOut_payload_0_9606);
  assign _zz_dataOut_payload_0_9656 = (_zz_dataOut_payload_0_9633 < _zz_dataOut_payload_0_9645);
  assign _zz_dataOut_payload_0_9657 = (_zz_dataOut_payload_0_9656 ? _zz_dataOut_payload_0_9633 : _zz_dataOut_payload_0_9645);
  assign _zz_dataOut_payload_0_9658 = (_zz_dataOut_payload_0_9656 ? _zz_dataOut_payload_0_9645 : _zz_dataOut_payload_0_9633);
  assign _zz_dataOut_payload_0_9659 = (_zz_dataOut_payload_0_9636 < _zz_dataOut_payload_0_9648);
  assign _zz_dataOut_payload_0_9660 = (_zz_dataOut_payload_0_9659 ? _zz_dataOut_payload_0_9636 : _zz_dataOut_payload_0_9648);
  assign _zz_dataOut_payload_0_9661 = (_zz_dataOut_payload_0_9659 ? _zz_dataOut_payload_0_9648 : _zz_dataOut_payload_0_9636);
  assign _zz_dataOut_payload_0_9662 = (_zz_dataOut_payload_0_9639 < _zz_dataOut_payload_0_9651);
  assign _zz_dataOut_payload_0_9663 = (_zz_dataOut_payload_0_9662 ? _zz_dataOut_payload_0_9639 : _zz_dataOut_payload_0_9651);
  assign _zz_dataOut_payload_0_9664 = (_zz_dataOut_payload_0_9662 ? _zz_dataOut_payload_0_9651 : _zz_dataOut_payload_0_9639);
  assign _zz_dataOut_payload_0_9665 = (_zz_dataOut_payload_0_9642 < _zz_dataOut_payload_0_9654);
  assign _zz_dataOut_payload_0_9666 = (_zz_dataOut_payload_0_9665 ? _zz_dataOut_payload_0_9642 : _zz_dataOut_payload_0_9654);
  assign _zz_dataOut_payload_0_9667 = (_zz_dataOut_payload_0_9665 ? _zz_dataOut_payload_0_9654 : _zz_dataOut_payload_0_9642);
  assign _zz_dataOut_payload_0_9668 = (_zz_dataOut_payload_0_9657 < _zz_dataOut_payload_0_9663);
  assign _zz_dataOut_payload_0_9669 = (_zz_dataOut_payload_0_9668 ? _zz_dataOut_payload_0_9657 : _zz_dataOut_payload_0_9663);
  assign _zz_dataOut_payload_0_9670 = (_zz_dataOut_payload_0_9668 ? _zz_dataOut_payload_0_9663 : _zz_dataOut_payload_0_9657);
  assign _zz_dataOut_payload_0_9671 = (_zz_dataOut_payload_0_9660 < _zz_dataOut_payload_0_9666);
  assign _zz_dataOut_payload_0_9672 = (_zz_dataOut_payload_0_9671 ? _zz_dataOut_payload_0_9660 : _zz_dataOut_payload_0_9666);
  assign _zz_dataOut_payload_0_9673 = (_zz_dataOut_payload_0_9671 ? _zz_dataOut_payload_0_9666 : _zz_dataOut_payload_0_9660);
  assign _zz_dataOut_payload_0_9674 = (_zz_dataOut_payload_0_9669 < _zz_dataOut_payload_0_9672);
  assign _zz_dataOut_payload_0_9675 = (_zz_dataOut_payload_0_9670 < _zz_dataOut_payload_0_9673);
  assign _zz_dataOut_payload_0_9680 = (_zz_dataOut_payload_0_9658 < _zz_dataOut_payload_0_9664);
  assign _zz_dataOut_payload_0_9681 = (_zz_dataOut_payload_0_9680 ? _zz_dataOut_payload_0_9658 : _zz_dataOut_payload_0_9664);
  assign _zz_dataOut_payload_0_9682 = (_zz_dataOut_payload_0_9680 ? _zz_dataOut_payload_0_9664 : _zz_dataOut_payload_0_9658);
  assign _zz_dataOut_payload_0_9683 = (_zz_dataOut_payload_0_9661 < _zz_dataOut_payload_0_9667);
  assign _zz_dataOut_payload_0_9684 = (_zz_dataOut_payload_0_9683 ? _zz_dataOut_payload_0_9661 : _zz_dataOut_payload_0_9667);
  assign _zz_dataOut_payload_0_9685 = (_zz_dataOut_payload_0_9683 ? _zz_dataOut_payload_0_9667 : _zz_dataOut_payload_0_9661);
  assign _zz_dataOut_payload_0_9686 = (_zz_dataOut_payload_0_9681 < _zz_dataOut_payload_0_9684);
  assign _zz_dataOut_payload_0_9687 = (_zz_dataOut_payload_0_9682 < _zz_dataOut_payload_0_9685);
  assign _zz_dataOut_payload_0_9700 = (_zz_dataOut_payload_0_9634 < _zz_dataOut_payload_0_9646);
  assign _zz_dataOut_payload_0_9701 = (_zz_dataOut_payload_0_9700 ? _zz_dataOut_payload_0_9634 : _zz_dataOut_payload_0_9646);
  assign _zz_dataOut_payload_0_9702 = (_zz_dataOut_payload_0_9700 ? _zz_dataOut_payload_0_9646 : _zz_dataOut_payload_0_9634);
  assign _zz_dataOut_payload_0_9703 = (_zz_dataOut_payload_0_9637 < _zz_dataOut_payload_0_9649);
  assign _zz_dataOut_payload_0_9704 = (_zz_dataOut_payload_0_9703 ? _zz_dataOut_payload_0_9637 : _zz_dataOut_payload_0_9649);
  assign _zz_dataOut_payload_0_9705 = (_zz_dataOut_payload_0_9703 ? _zz_dataOut_payload_0_9649 : _zz_dataOut_payload_0_9637);
  assign _zz_dataOut_payload_0_9706 = (_zz_dataOut_payload_0_9640 < _zz_dataOut_payload_0_9652);
  assign _zz_dataOut_payload_0_9707 = (_zz_dataOut_payload_0_9706 ? _zz_dataOut_payload_0_9640 : _zz_dataOut_payload_0_9652);
  assign _zz_dataOut_payload_0_9708 = (_zz_dataOut_payload_0_9706 ? _zz_dataOut_payload_0_9652 : _zz_dataOut_payload_0_9640);
  assign _zz_dataOut_payload_0_9709 = (_zz_dataOut_payload_0_9643 < _zz_dataOut_payload_0_9655);
  assign _zz_dataOut_payload_0_9710 = (_zz_dataOut_payload_0_9709 ? _zz_dataOut_payload_0_9643 : _zz_dataOut_payload_0_9655);
  assign _zz_dataOut_payload_0_9711 = (_zz_dataOut_payload_0_9709 ? _zz_dataOut_payload_0_9655 : _zz_dataOut_payload_0_9643);
  assign _zz_dataOut_payload_0_9712 = (_zz_dataOut_payload_0_9701 < _zz_dataOut_payload_0_9707);
  assign _zz_dataOut_payload_0_9713 = (_zz_dataOut_payload_0_9712 ? _zz_dataOut_payload_0_9701 : _zz_dataOut_payload_0_9707);
  assign _zz_dataOut_payload_0_9714 = (_zz_dataOut_payload_0_9712 ? _zz_dataOut_payload_0_9707 : _zz_dataOut_payload_0_9701);
  assign _zz_dataOut_payload_0_9715 = (_zz_dataOut_payload_0_9704 < _zz_dataOut_payload_0_9710);
  assign _zz_dataOut_payload_0_9716 = (_zz_dataOut_payload_0_9715 ? _zz_dataOut_payload_0_9704 : _zz_dataOut_payload_0_9710);
  assign _zz_dataOut_payload_0_9717 = (_zz_dataOut_payload_0_9715 ? _zz_dataOut_payload_0_9710 : _zz_dataOut_payload_0_9704);
  assign _zz_dataOut_payload_0_9718 = (_zz_dataOut_payload_0_9713 < _zz_dataOut_payload_0_9716);
  assign _zz_dataOut_payload_0_9719 = (_zz_dataOut_payload_0_9714 < _zz_dataOut_payload_0_9717);
  assign _zz_dataOut_payload_0_9724 = (_zz_dataOut_payload_0_9702 < _zz_dataOut_payload_0_9708);
  assign _zz_dataOut_payload_0_9725 = (_zz_dataOut_payload_0_9724 ? _zz_dataOut_payload_0_9702 : _zz_dataOut_payload_0_9708);
  assign _zz_dataOut_payload_0_9726 = (_zz_dataOut_payload_0_9724 ? _zz_dataOut_payload_0_9708 : _zz_dataOut_payload_0_9702);
  assign _zz_dataOut_payload_0_9727 = (_zz_dataOut_payload_0_9705 < _zz_dataOut_payload_0_9711);
  assign _zz_dataOut_payload_0_9728 = (_zz_dataOut_payload_0_9727 ? _zz_dataOut_payload_0_9705 : _zz_dataOut_payload_0_9711);
  assign _zz_dataOut_payload_0_9729 = (_zz_dataOut_payload_0_9727 ? _zz_dataOut_payload_0_9711 : _zz_dataOut_payload_0_9705);
  assign _zz_dataOut_payload_0_9730 = (_zz_dataOut_payload_0_9725 < _zz_dataOut_payload_0_9728);
  assign _zz_dataOut_payload_0_9731 = (_zz_dataOut_payload_0_9726 < _zz_dataOut_payload_0_9729);
  assign _zz_dataOut_payload_0_9760 = (_zz_dataOut_payload_0_9586 < _zz_dataOut_payload_0_9610);
  assign _zz_dataOut_payload_0_9761 = (_zz_dataOut_payload_0_9760 ? _zz_dataOut_payload_0_9586 : _zz_dataOut_payload_0_9610);
  assign _zz_dataOut_payload_0_9762 = (_zz_dataOut_payload_0_9760 ? _zz_dataOut_payload_0_9610 : _zz_dataOut_payload_0_9586);
  assign _zz_dataOut_payload_0_9763 = (_zz_dataOut_payload_0_9589 < _zz_dataOut_payload_0_9613);
  assign _zz_dataOut_payload_0_9764 = (_zz_dataOut_payload_0_9763 ? _zz_dataOut_payload_0_9589 : _zz_dataOut_payload_0_9613);
  assign _zz_dataOut_payload_0_9765 = (_zz_dataOut_payload_0_9763 ? _zz_dataOut_payload_0_9613 : _zz_dataOut_payload_0_9589);
  assign _zz_dataOut_payload_0_9766 = (_zz_dataOut_payload_0_9592 < _zz_dataOut_payload_0_9616);
  assign _zz_dataOut_payload_0_9767 = (_zz_dataOut_payload_0_9766 ? _zz_dataOut_payload_0_9592 : _zz_dataOut_payload_0_9616);
  assign _zz_dataOut_payload_0_9768 = (_zz_dataOut_payload_0_9766 ? _zz_dataOut_payload_0_9616 : _zz_dataOut_payload_0_9592);
  assign _zz_dataOut_payload_0_9769 = (_zz_dataOut_payload_0_9595 < _zz_dataOut_payload_0_9619);
  assign _zz_dataOut_payload_0_9770 = (_zz_dataOut_payload_0_9769 ? _zz_dataOut_payload_0_9595 : _zz_dataOut_payload_0_9619);
  assign _zz_dataOut_payload_0_9771 = (_zz_dataOut_payload_0_9769 ? _zz_dataOut_payload_0_9619 : _zz_dataOut_payload_0_9595);
  assign _zz_dataOut_payload_0_9772 = (_zz_dataOut_payload_0_9598 < _zz_dataOut_payload_0_9622);
  assign _zz_dataOut_payload_0_9773 = (_zz_dataOut_payload_0_9772 ? _zz_dataOut_payload_0_9598 : _zz_dataOut_payload_0_9622);
  assign _zz_dataOut_payload_0_9774 = (_zz_dataOut_payload_0_9772 ? _zz_dataOut_payload_0_9622 : _zz_dataOut_payload_0_9598);
  assign _zz_dataOut_payload_0_9775 = (_zz_dataOut_payload_0_9601 < _zz_dataOut_payload_0_9625);
  assign _zz_dataOut_payload_0_9776 = (_zz_dataOut_payload_0_9775 ? _zz_dataOut_payload_0_9601 : _zz_dataOut_payload_0_9625);
  assign _zz_dataOut_payload_0_9777 = (_zz_dataOut_payload_0_9775 ? _zz_dataOut_payload_0_9625 : _zz_dataOut_payload_0_9601);
  assign _zz_dataOut_payload_0_9778 = (_zz_dataOut_payload_0_9604 < _zz_dataOut_payload_0_9628);
  assign _zz_dataOut_payload_0_9779 = (_zz_dataOut_payload_0_9778 ? _zz_dataOut_payload_0_9604 : _zz_dataOut_payload_0_9628);
  assign _zz_dataOut_payload_0_9780 = (_zz_dataOut_payload_0_9778 ? _zz_dataOut_payload_0_9628 : _zz_dataOut_payload_0_9604);
  assign _zz_dataOut_payload_0_9781 = (_zz_dataOut_payload_0_9607 < _zz_dataOut_payload_0_9631);
  assign _zz_dataOut_payload_0_9782 = (_zz_dataOut_payload_0_9781 ? _zz_dataOut_payload_0_9607 : _zz_dataOut_payload_0_9631);
  assign _zz_dataOut_payload_0_9783 = (_zz_dataOut_payload_0_9781 ? _zz_dataOut_payload_0_9631 : _zz_dataOut_payload_0_9607);
  assign _zz_dataOut_payload_0_9784 = (_zz_dataOut_payload_0_9761 < _zz_dataOut_payload_0_9773);
  assign _zz_dataOut_payload_0_9785 = (_zz_dataOut_payload_0_9784 ? _zz_dataOut_payload_0_9761 : _zz_dataOut_payload_0_9773);
  assign _zz_dataOut_payload_0_9786 = (_zz_dataOut_payload_0_9784 ? _zz_dataOut_payload_0_9773 : _zz_dataOut_payload_0_9761);
  assign _zz_dataOut_payload_0_9787 = (_zz_dataOut_payload_0_9764 < _zz_dataOut_payload_0_9776);
  assign _zz_dataOut_payload_0_9788 = (_zz_dataOut_payload_0_9787 ? _zz_dataOut_payload_0_9764 : _zz_dataOut_payload_0_9776);
  assign _zz_dataOut_payload_0_9789 = (_zz_dataOut_payload_0_9787 ? _zz_dataOut_payload_0_9776 : _zz_dataOut_payload_0_9764);
  assign _zz_dataOut_payload_0_9790 = (_zz_dataOut_payload_0_9767 < _zz_dataOut_payload_0_9779);
  assign _zz_dataOut_payload_0_9791 = (_zz_dataOut_payload_0_9790 ? _zz_dataOut_payload_0_9767 : _zz_dataOut_payload_0_9779);
  assign _zz_dataOut_payload_0_9792 = (_zz_dataOut_payload_0_9790 ? _zz_dataOut_payload_0_9779 : _zz_dataOut_payload_0_9767);
  assign _zz_dataOut_payload_0_9793 = (_zz_dataOut_payload_0_9770 < _zz_dataOut_payload_0_9782);
  assign _zz_dataOut_payload_0_9794 = (_zz_dataOut_payload_0_9793 ? _zz_dataOut_payload_0_9770 : _zz_dataOut_payload_0_9782);
  assign _zz_dataOut_payload_0_9795 = (_zz_dataOut_payload_0_9793 ? _zz_dataOut_payload_0_9782 : _zz_dataOut_payload_0_9770);
  assign _zz_dataOut_payload_0_9796 = (_zz_dataOut_payload_0_9785 < _zz_dataOut_payload_0_9791);
  assign _zz_dataOut_payload_0_9797 = (_zz_dataOut_payload_0_9796 ? _zz_dataOut_payload_0_9785 : _zz_dataOut_payload_0_9791);
  assign _zz_dataOut_payload_0_9798 = (_zz_dataOut_payload_0_9796 ? _zz_dataOut_payload_0_9791 : _zz_dataOut_payload_0_9785);
  assign _zz_dataOut_payload_0_9799 = (_zz_dataOut_payload_0_9788 < _zz_dataOut_payload_0_9794);
  assign _zz_dataOut_payload_0_9800 = (_zz_dataOut_payload_0_9799 ? _zz_dataOut_payload_0_9788 : _zz_dataOut_payload_0_9794);
  assign _zz_dataOut_payload_0_9801 = (_zz_dataOut_payload_0_9799 ? _zz_dataOut_payload_0_9794 : _zz_dataOut_payload_0_9788);
  assign _zz_dataOut_payload_0_9802 = (_zz_dataOut_payload_0_9797 < _zz_dataOut_payload_0_9800);
  assign _zz_dataOut_payload_0_9803 = (_zz_dataOut_payload_0_9798 < _zz_dataOut_payload_0_9801);
  assign _zz_dataOut_payload_0_9808 = (_zz_dataOut_payload_0_9786 < _zz_dataOut_payload_0_9792);
  assign _zz_dataOut_payload_0_9809 = (_zz_dataOut_payload_0_9808 ? _zz_dataOut_payload_0_9786 : _zz_dataOut_payload_0_9792);
  assign _zz_dataOut_payload_0_9810 = (_zz_dataOut_payload_0_9808 ? _zz_dataOut_payload_0_9792 : _zz_dataOut_payload_0_9786);
  assign _zz_dataOut_payload_0_9811 = (_zz_dataOut_payload_0_9789 < _zz_dataOut_payload_0_9795);
  assign _zz_dataOut_payload_0_9812 = (_zz_dataOut_payload_0_9811 ? _zz_dataOut_payload_0_9789 : _zz_dataOut_payload_0_9795);
  assign _zz_dataOut_payload_0_9813 = (_zz_dataOut_payload_0_9811 ? _zz_dataOut_payload_0_9795 : _zz_dataOut_payload_0_9789);
  assign _zz_dataOut_payload_0_9814 = (_zz_dataOut_payload_0_9809 < _zz_dataOut_payload_0_9812);
  assign _zz_dataOut_payload_0_9815 = (_zz_dataOut_payload_0_9810 < _zz_dataOut_payload_0_9813);
  assign _zz_dataOut_payload_0_9828 = (_zz_dataOut_payload_0_9762 < _zz_dataOut_payload_0_9774);
  assign _zz_dataOut_payload_0_9829 = (_zz_dataOut_payload_0_9828 ? _zz_dataOut_payload_0_9762 : _zz_dataOut_payload_0_9774);
  assign _zz_dataOut_payload_0_9830 = (_zz_dataOut_payload_0_9828 ? _zz_dataOut_payload_0_9774 : _zz_dataOut_payload_0_9762);
  assign _zz_dataOut_payload_0_9831 = (_zz_dataOut_payload_0_9765 < _zz_dataOut_payload_0_9777);
  assign _zz_dataOut_payload_0_9832 = (_zz_dataOut_payload_0_9831 ? _zz_dataOut_payload_0_9765 : _zz_dataOut_payload_0_9777);
  assign _zz_dataOut_payload_0_9833 = (_zz_dataOut_payload_0_9831 ? _zz_dataOut_payload_0_9777 : _zz_dataOut_payload_0_9765);
  assign _zz_dataOut_payload_0_9834 = (_zz_dataOut_payload_0_9768 < _zz_dataOut_payload_0_9780);
  assign _zz_dataOut_payload_0_9835 = (_zz_dataOut_payload_0_9834 ? _zz_dataOut_payload_0_9768 : _zz_dataOut_payload_0_9780);
  assign _zz_dataOut_payload_0_9836 = (_zz_dataOut_payload_0_9834 ? _zz_dataOut_payload_0_9780 : _zz_dataOut_payload_0_9768);
  assign _zz_dataOut_payload_0_9837 = (_zz_dataOut_payload_0_9771 < _zz_dataOut_payload_0_9783);
  assign _zz_dataOut_payload_0_9838 = (_zz_dataOut_payload_0_9837 ? _zz_dataOut_payload_0_9771 : _zz_dataOut_payload_0_9783);
  assign _zz_dataOut_payload_0_9839 = (_zz_dataOut_payload_0_9837 ? _zz_dataOut_payload_0_9783 : _zz_dataOut_payload_0_9771);
  assign _zz_dataOut_payload_0_9840 = (_zz_dataOut_payload_0_9829 < _zz_dataOut_payload_0_9835);
  assign _zz_dataOut_payload_0_9841 = (_zz_dataOut_payload_0_9840 ? _zz_dataOut_payload_0_9829 : _zz_dataOut_payload_0_9835);
  assign _zz_dataOut_payload_0_9842 = (_zz_dataOut_payload_0_9840 ? _zz_dataOut_payload_0_9835 : _zz_dataOut_payload_0_9829);
  assign _zz_dataOut_payload_0_9843 = (_zz_dataOut_payload_0_9832 < _zz_dataOut_payload_0_9838);
  assign _zz_dataOut_payload_0_9844 = (_zz_dataOut_payload_0_9843 ? _zz_dataOut_payload_0_9832 : _zz_dataOut_payload_0_9838);
  assign _zz_dataOut_payload_0_9845 = (_zz_dataOut_payload_0_9843 ? _zz_dataOut_payload_0_9838 : _zz_dataOut_payload_0_9832);
  assign _zz_dataOut_payload_0_9846 = (_zz_dataOut_payload_0_9841 < _zz_dataOut_payload_0_9844);
  assign _zz_dataOut_payload_0_9847 = (_zz_dataOut_payload_0_9842 < _zz_dataOut_payload_0_9845);
  assign _zz_dataOut_payload_0_9852 = (_zz_dataOut_payload_0_9830 < _zz_dataOut_payload_0_9836);
  assign _zz_dataOut_payload_0_9853 = (_zz_dataOut_payload_0_9852 ? _zz_dataOut_payload_0_9830 : _zz_dataOut_payload_0_9836);
  assign _zz_dataOut_payload_0_9854 = (_zz_dataOut_payload_0_9852 ? _zz_dataOut_payload_0_9836 : _zz_dataOut_payload_0_9830);
  assign _zz_dataOut_payload_0_9855 = (_zz_dataOut_payload_0_9833 < _zz_dataOut_payload_0_9839);
  assign _zz_dataOut_payload_0_9856 = (_zz_dataOut_payload_0_9855 ? _zz_dataOut_payload_0_9833 : _zz_dataOut_payload_0_9839);
  assign _zz_dataOut_payload_0_9857 = (_zz_dataOut_payload_0_9855 ? _zz_dataOut_payload_0_9839 : _zz_dataOut_payload_0_9833);
  assign _zz_dataOut_payload_0_9858 = (_zz_dataOut_payload_0_9853 < _zz_dataOut_payload_0_9856);
  assign _zz_dataOut_payload_0_9859 = (_zz_dataOut_payload_0_9854 < _zz_dataOut_payload_0_9857);
  assign _zz_dataOut_payload_0_9984 = (_zz_dataOut_payload_0_8192 < _zz_dataOut_payload_0_8255);
  assign _zz_dataOut_payload_0_9985 = (_zz_dataOut_payload_0_9984 ? _zz_dataOut_payload_0_8192 : _zz_dataOut_payload_0_8255);
  assign _zz_dataOut_payload_0_9986 = (_zz_dataOut_payload_0_9984 ? _zz_dataOut_payload_0_8255 : _zz_dataOut_payload_0_8192);
  assign _zz_dataOut_payload_0_9987 = (_zz_dataOut_payload_0_8193 < _zz_dataOut_payload_0_8254);
  assign _zz_dataOut_payload_0_9988 = (_zz_dataOut_payload_0_9987 ? _zz_dataOut_payload_0_8193 : _zz_dataOut_payload_0_8254);
  assign _zz_dataOut_payload_0_9989 = (_zz_dataOut_payload_0_9987 ? _zz_dataOut_payload_0_8254 : _zz_dataOut_payload_0_8193);
  assign _zz_dataOut_payload_0_9990 = (_zz_dataOut_payload_0_8194 < _zz_dataOut_payload_0_8253);
  assign _zz_dataOut_payload_0_9991 = (_zz_dataOut_payload_0_9990 ? _zz_dataOut_payload_0_8194 : _zz_dataOut_payload_0_8253);
  assign _zz_dataOut_payload_0_9992 = (_zz_dataOut_payload_0_9990 ? _zz_dataOut_payload_0_8253 : _zz_dataOut_payload_0_8194);
  assign _zz_dataOut_payload_0_9993 = (_zz_dataOut_payload_0_8195 < _zz_dataOut_payload_0_8252);
  assign _zz_dataOut_payload_0_9994 = (_zz_dataOut_payload_0_9993 ? _zz_dataOut_payload_0_8195 : _zz_dataOut_payload_0_8252);
  assign _zz_dataOut_payload_0_9995 = (_zz_dataOut_payload_0_9993 ? _zz_dataOut_payload_0_8252 : _zz_dataOut_payload_0_8195);
  assign _zz_dataOut_payload_0_9996 = (_zz_dataOut_payload_0_8196 < _zz_dataOut_payload_0_8251);
  assign _zz_dataOut_payload_0_9997 = (_zz_dataOut_payload_0_9996 ? _zz_dataOut_payload_0_8196 : _zz_dataOut_payload_0_8251);
  assign _zz_dataOut_payload_0_9998 = (_zz_dataOut_payload_0_9996 ? _zz_dataOut_payload_0_8251 : _zz_dataOut_payload_0_8196);
  assign _zz_dataOut_payload_0_9999 = (_zz_dataOut_payload_0_8197 < _zz_dataOut_payload_0_8250);
  assign _zz_dataOut_payload_0_10000 = (_zz_dataOut_payload_0_9999 ? _zz_dataOut_payload_0_8197 : _zz_dataOut_payload_0_8250);
  assign _zz_dataOut_payload_0_10001 = (_zz_dataOut_payload_0_9999 ? _zz_dataOut_payload_0_8250 : _zz_dataOut_payload_0_8197);
  assign _zz_dataOut_payload_0_10002 = (_zz_dataOut_payload_0_8198 < _zz_dataOut_payload_0_8249);
  assign _zz_dataOut_payload_0_10003 = (_zz_dataOut_payload_0_10002 ? _zz_dataOut_payload_0_8198 : _zz_dataOut_payload_0_8249);
  assign _zz_dataOut_payload_0_10004 = (_zz_dataOut_payload_0_10002 ? _zz_dataOut_payload_0_8249 : _zz_dataOut_payload_0_8198);
  assign _zz_dataOut_payload_0_10005 = (_zz_dataOut_payload_0_8199 < _zz_dataOut_payload_0_8248);
  assign _zz_dataOut_payload_0_10006 = (_zz_dataOut_payload_0_10005 ? _zz_dataOut_payload_0_8199 : _zz_dataOut_payload_0_8248);
  assign _zz_dataOut_payload_0_10007 = (_zz_dataOut_payload_0_10005 ? _zz_dataOut_payload_0_8248 : _zz_dataOut_payload_0_8199);
  assign _zz_dataOut_payload_0_10008 = (_zz_dataOut_payload_0_8200 < _zz_dataOut_payload_0_8247);
  assign _zz_dataOut_payload_0_10009 = (_zz_dataOut_payload_0_10008 ? _zz_dataOut_payload_0_8200 : _zz_dataOut_payload_0_8247);
  assign _zz_dataOut_payload_0_10010 = (_zz_dataOut_payload_0_10008 ? _zz_dataOut_payload_0_8247 : _zz_dataOut_payload_0_8200);
  assign _zz_dataOut_payload_0_10011 = (_zz_dataOut_payload_0_8201 < _zz_dataOut_payload_0_8246);
  assign _zz_dataOut_payload_0_10012 = (_zz_dataOut_payload_0_10011 ? _zz_dataOut_payload_0_8201 : _zz_dataOut_payload_0_8246);
  assign _zz_dataOut_payload_0_10013 = (_zz_dataOut_payload_0_10011 ? _zz_dataOut_payload_0_8246 : _zz_dataOut_payload_0_8201);
  assign _zz_dataOut_payload_0_10014 = (_zz_dataOut_payload_0_8202 < _zz_dataOut_payload_0_8245);
  assign _zz_dataOut_payload_0_10015 = (_zz_dataOut_payload_0_10014 ? _zz_dataOut_payload_0_8202 : _zz_dataOut_payload_0_8245);
  assign _zz_dataOut_payload_0_10016 = (_zz_dataOut_payload_0_10014 ? _zz_dataOut_payload_0_8245 : _zz_dataOut_payload_0_8202);
  assign _zz_dataOut_payload_0_10017 = (_zz_dataOut_payload_0_8203 < _zz_dataOut_payload_0_8244);
  assign _zz_dataOut_payload_0_10018 = (_zz_dataOut_payload_0_10017 ? _zz_dataOut_payload_0_8203 : _zz_dataOut_payload_0_8244);
  assign _zz_dataOut_payload_0_10019 = (_zz_dataOut_payload_0_10017 ? _zz_dataOut_payload_0_8244 : _zz_dataOut_payload_0_8203);
  assign _zz_dataOut_payload_0_10020 = (_zz_dataOut_payload_0_8204 < _zz_dataOut_payload_0_8243);
  assign _zz_dataOut_payload_0_10021 = (_zz_dataOut_payload_0_10020 ? _zz_dataOut_payload_0_8204 : _zz_dataOut_payload_0_8243);
  assign _zz_dataOut_payload_0_10022 = (_zz_dataOut_payload_0_10020 ? _zz_dataOut_payload_0_8243 : _zz_dataOut_payload_0_8204);
  assign _zz_dataOut_payload_0_10023 = (_zz_dataOut_payload_0_8205 < _zz_dataOut_payload_0_8242);
  assign _zz_dataOut_payload_0_10024 = (_zz_dataOut_payload_0_10023 ? _zz_dataOut_payload_0_8205 : _zz_dataOut_payload_0_8242);
  assign _zz_dataOut_payload_0_10025 = (_zz_dataOut_payload_0_10023 ? _zz_dataOut_payload_0_8242 : _zz_dataOut_payload_0_8205);
  assign _zz_dataOut_payload_0_10026 = (_zz_dataOut_payload_0_8206 < _zz_dataOut_payload_0_8241);
  assign _zz_dataOut_payload_0_10027 = (_zz_dataOut_payload_0_10026 ? _zz_dataOut_payload_0_8206 : _zz_dataOut_payload_0_8241);
  assign _zz_dataOut_payload_0_10028 = (_zz_dataOut_payload_0_10026 ? _zz_dataOut_payload_0_8241 : _zz_dataOut_payload_0_8206);
  assign _zz_dataOut_payload_0_10029 = (_zz_dataOut_payload_0_8207 < _zz_dataOut_payload_0_8240);
  assign _zz_dataOut_payload_0_10030 = (_zz_dataOut_payload_0_10029 ? _zz_dataOut_payload_0_8207 : _zz_dataOut_payload_0_8240);
  assign _zz_dataOut_payload_0_10031 = (_zz_dataOut_payload_0_10029 ? _zz_dataOut_payload_0_8240 : _zz_dataOut_payload_0_8207);
  assign _zz_dataOut_payload_0_10032 = (_zz_dataOut_payload_0_8208 < _zz_dataOut_payload_0_8239);
  assign _zz_dataOut_payload_0_10033 = (_zz_dataOut_payload_0_10032 ? _zz_dataOut_payload_0_8208 : _zz_dataOut_payload_0_8239);
  assign _zz_dataOut_payload_0_10034 = (_zz_dataOut_payload_0_10032 ? _zz_dataOut_payload_0_8239 : _zz_dataOut_payload_0_8208);
  assign _zz_dataOut_payload_0_10035 = (_zz_dataOut_payload_0_8209 < _zz_dataOut_payload_0_8238);
  assign _zz_dataOut_payload_0_10036 = (_zz_dataOut_payload_0_10035 ? _zz_dataOut_payload_0_8209 : _zz_dataOut_payload_0_8238);
  assign _zz_dataOut_payload_0_10037 = (_zz_dataOut_payload_0_10035 ? _zz_dataOut_payload_0_8238 : _zz_dataOut_payload_0_8209);
  assign _zz_dataOut_payload_0_10038 = (_zz_dataOut_payload_0_8210 < _zz_dataOut_payload_0_8237);
  assign _zz_dataOut_payload_0_10039 = (_zz_dataOut_payload_0_10038 ? _zz_dataOut_payload_0_8210 : _zz_dataOut_payload_0_8237);
  assign _zz_dataOut_payload_0_10040 = (_zz_dataOut_payload_0_10038 ? _zz_dataOut_payload_0_8237 : _zz_dataOut_payload_0_8210);
  assign _zz_dataOut_payload_0_10041 = (_zz_dataOut_payload_0_8211 < _zz_dataOut_payload_0_8236);
  assign _zz_dataOut_payload_0_10042 = (_zz_dataOut_payload_0_10041 ? _zz_dataOut_payload_0_8211 : _zz_dataOut_payload_0_8236);
  assign _zz_dataOut_payload_0_10043 = (_zz_dataOut_payload_0_10041 ? _zz_dataOut_payload_0_8236 : _zz_dataOut_payload_0_8211);
  assign _zz_dataOut_payload_0_10044 = (_zz_dataOut_payload_0_8212 < _zz_dataOut_payload_0_8235);
  assign _zz_dataOut_payload_0_10045 = (_zz_dataOut_payload_0_10044 ? _zz_dataOut_payload_0_8212 : _zz_dataOut_payload_0_8235);
  assign _zz_dataOut_payload_0_10046 = (_zz_dataOut_payload_0_10044 ? _zz_dataOut_payload_0_8235 : _zz_dataOut_payload_0_8212);
  assign _zz_dataOut_payload_0_10047 = (_zz_dataOut_payload_0_8213 < _zz_dataOut_payload_0_8234);
  assign _zz_dataOut_payload_0_10048 = (_zz_dataOut_payload_0_10047 ? _zz_dataOut_payload_0_8213 : _zz_dataOut_payload_0_8234);
  assign _zz_dataOut_payload_0_10049 = (_zz_dataOut_payload_0_10047 ? _zz_dataOut_payload_0_8234 : _zz_dataOut_payload_0_8213);
  assign _zz_dataOut_payload_0_10050 = (_zz_dataOut_payload_0_8214 < _zz_dataOut_payload_0_8233);
  assign _zz_dataOut_payload_0_10051 = (_zz_dataOut_payload_0_10050 ? _zz_dataOut_payload_0_8214 : _zz_dataOut_payload_0_8233);
  assign _zz_dataOut_payload_0_10052 = (_zz_dataOut_payload_0_10050 ? _zz_dataOut_payload_0_8233 : _zz_dataOut_payload_0_8214);
  assign _zz_dataOut_payload_0_10053 = (_zz_dataOut_payload_0_8215 < _zz_dataOut_payload_0_8232);
  assign _zz_dataOut_payload_0_10054 = (_zz_dataOut_payload_0_10053 ? _zz_dataOut_payload_0_8215 : _zz_dataOut_payload_0_8232);
  assign _zz_dataOut_payload_0_10055 = (_zz_dataOut_payload_0_10053 ? _zz_dataOut_payload_0_8232 : _zz_dataOut_payload_0_8215);
  assign _zz_dataOut_payload_0_10056 = (_zz_dataOut_payload_0_8216 < _zz_dataOut_payload_0_8231);
  assign _zz_dataOut_payload_0_10057 = (_zz_dataOut_payload_0_10056 ? _zz_dataOut_payload_0_8216 : _zz_dataOut_payload_0_8231);
  assign _zz_dataOut_payload_0_10058 = (_zz_dataOut_payload_0_10056 ? _zz_dataOut_payload_0_8231 : _zz_dataOut_payload_0_8216);
  assign _zz_dataOut_payload_0_10059 = (_zz_dataOut_payload_0_8217 < _zz_dataOut_payload_0_8230);
  assign _zz_dataOut_payload_0_10060 = (_zz_dataOut_payload_0_10059 ? _zz_dataOut_payload_0_8217 : _zz_dataOut_payload_0_8230);
  assign _zz_dataOut_payload_0_10061 = (_zz_dataOut_payload_0_10059 ? _zz_dataOut_payload_0_8230 : _zz_dataOut_payload_0_8217);
  assign _zz_dataOut_payload_0_10062 = (_zz_dataOut_payload_0_8218 < _zz_dataOut_payload_0_8229);
  assign _zz_dataOut_payload_0_10063 = (_zz_dataOut_payload_0_10062 ? _zz_dataOut_payload_0_8218 : _zz_dataOut_payload_0_8229);
  assign _zz_dataOut_payload_0_10064 = (_zz_dataOut_payload_0_10062 ? _zz_dataOut_payload_0_8229 : _zz_dataOut_payload_0_8218);
  assign _zz_dataOut_payload_0_10065 = (_zz_dataOut_payload_0_8219 < _zz_dataOut_payload_0_8228);
  assign _zz_dataOut_payload_0_10066 = (_zz_dataOut_payload_0_10065 ? _zz_dataOut_payload_0_8219 : _zz_dataOut_payload_0_8228);
  assign _zz_dataOut_payload_0_10067 = (_zz_dataOut_payload_0_10065 ? _zz_dataOut_payload_0_8228 : _zz_dataOut_payload_0_8219);
  assign _zz_dataOut_payload_0_10068 = (_zz_dataOut_payload_0_8220 < _zz_dataOut_payload_0_8227);
  assign _zz_dataOut_payload_0_10069 = (_zz_dataOut_payload_0_10068 ? _zz_dataOut_payload_0_8220 : _zz_dataOut_payload_0_8227);
  assign _zz_dataOut_payload_0_10070 = (_zz_dataOut_payload_0_10068 ? _zz_dataOut_payload_0_8227 : _zz_dataOut_payload_0_8220);
  assign _zz_dataOut_payload_0_10071 = (_zz_dataOut_payload_0_8221 < _zz_dataOut_payload_0_8226);
  assign _zz_dataOut_payload_0_10072 = (_zz_dataOut_payload_0_10071 ? _zz_dataOut_payload_0_8221 : _zz_dataOut_payload_0_8226);
  assign _zz_dataOut_payload_0_10073 = (_zz_dataOut_payload_0_10071 ? _zz_dataOut_payload_0_8226 : _zz_dataOut_payload_0_8221);
  assign _zz_dataOut_payload_0_10074 = (_zz_dataOut_payload_0_8222 < _zz_dataOut_payload_0_8225);
  assign _zz_dataOut_payload_0_10075 = (_zz_dataOut_payload_0_10074 ? _zz_dataOut_payload_0_8222 : _zz_dataOut_payload_0_8225);
  assign _zz_dataOut_payload_0_10076 = (_zz_dataOut_payload_0_10074 ? _zz_dataOut_payload_0_8225 : _zz_dataOut_payload_0_8222);
  assign _zz_dataOut_payload_0_10077 = (_zz_dataOut_payload_0_8223 < _zz_dataOut_payload_0_8224);
  assign _zz_dataOut_payload_0_10078 = (_zz_dataOut_payload_0_10077 ? _zz_dataOut_payload_0_8223 : _zz_dataOut_payload_0_8224);
  assign _zz_dataOut_payload_0_10079 = (_zz_dataOut_payload_0_10077 ? _zz_dataOut_payload_0_8224 : _zz_dataOut_payload_0_8223);
  assign _zz_dataOut_payload_0_10080 = (_zz_dataOut_payload_0_9985 < _zz_dataOut_payload_0_10033);
  assign _zz_dataOut_payload_0_10081 = (_zz_dataOut_payload_0_10080 ? _zz_dataOut_payload_0_9985 : _zz_dataOut_payload_0_10033);
  assign _zz_dataOut_payload_0_10082 = (_zz_dataOut_payload_0_10080 ? _zz_dataOut_payload_0_10033 : _zz_dataOut_payload_0_9985);
  assign _zz_dataOut_payload_0_10083 = (_zz_dataOut_payload_0_9988 < _zz_dataOut_payload_0_10036);
  assign _zz_dataOut_payload_0_10084 = (_zz_dataOut_payload_0_10083 ? _zz_dataOut_payload_0_9988 : _zz_dataOut_payload_0_10036);
  assign _zz_dataOut_payload_0_10085 = (_zz_dataOut_payload_0_10083 ? _zz_dataOut_payload_0_10036 : _zz_dataOut_payload_0_9988);
  assign _zz_dataOut_payload_0_10086 = (_zz_dataOut_payload_0_9991 < _zz_dataOut_payload_0_10039);
  assign _zz_dataOut_payload_0_10087 = (_zz_dataOut_payload_0_10086 ? _zz_dataOut_payload_0_9991 : _zz_dataOut_payload_0_10039);
  assign _zz_dataOut_payload_0_10088 = (_zz_dataOut_payload_0_10086 ? _zz_dataOut_payload_0_10039 : _zz_dataOut_payload_0_9991);
  assign _zz_dataOut_payload_0_10089 = (_zz_dataOut_payload_0_9994 < _zz_dataOut_payload_0_10042);
  assign _zz_dataOut_payload_0_10090 = (_zz_dataOut_payload_0_10089 ? _zz_dataOut_payload_0_9994 : _zz_dataOut_payload_0_10042);
  assign _zz_dataOut_payload_0_10091 = (_zz_dataOut_payload_0_10089 ? _zz_dataOut_payload_0_10042 : _zz_dataOut_payload_0_9994);
  assign _zz_dataOut_payload_0_10092 = (_zz_dataOut_payload_0_9997 < _zz_dataOut_payload_0_10045);
  assign _zz_dataOut_payload_0_10093 = (_zz_dataOut_payload_0_10092 ? _zz_dataOut_payload_0_9997 : _zz_dataOut_payload_0_10045);
  assign _zz_dataOut_payload_0_10094 = (_zz_dataOut_payload_0_10092 ? _zz_dataOut_payload_0_10045 : _zz_dataOut_payload_0_9997);
  assign _zz_dataOut_payload_0_10095 = (_zz_dataOut_payload_0_10000 < _zz_dataOut_payload_0_10048);
  assign _zz_dataOut_payload_0_10096 = (_zz_dataOut_payload_0_10095 ? _zz_dataOut_payload_0_10000 : _zz_dataOut_payload_0_10048);
  assign _zz_dataOut_payload_0_10097 = (_zz_dataOut_payload_0_10095 ? _zz_dataOut_payload_0_10048 : _zz_dataOut_payload_0_10000);
  assign _zz_dataOut_payload_0_10098 = (_zz_dataOut_payload_0_10003 < _zz_dataOut_payload_0_10051);
  assign _zz_dataOut_payload_0_10099 = (_zz_dataOut_payload_0_10098 ? _zz_dataOut_payload_0_10003 : _zz_dataOut_payload_0_10051);
  assign _zz_dataOut_payload_0_10100 = (_zz_dataOut_payload_0_10098 ? _zz_dataOut_payload_0_10051 : _zz_dataOut_payload_0_10003);
  assign _zz_dataOut_payload_0_10101 = (_zz_dataOut_payload_0_10006 < _zz_dataOut_payload_0_10054);
  assign _zz_dataOut_payload_0_10102 = (_zz_dataOut_payload_0_10101 ? _zz_dataOut_payload_0_10006 : _zz_dataOut_payload_0_10054);
  assign _zz_dataOut_payload_0_10103 = (_zz_dataOut_payload_0_10101 ? _zz_dataOut_payload_0_10054 : _zz_dataOut_payload_0_10006);
  assign _zz_dataOut_payload_0_10104 = (_zz_dataOut_payload_0_10009 < _zz_dataOut_payload_0_10057);
  assign _zz_dataOut_payload_0_10105 = (_zz_dataOut_payload_0_10104 ? _zz_dataOut_payload_0_10009 : _zz_dataOut_payload_0_10057);
  assign _zz_dataOut_payload_0_10106 = (_zz_dataOut_payload_0_10104 ? _zz_dataOut_payload_0_10057 : _zz_dataOut_payload_0_10009);
  assign _zz_dataOut_payload_0_10107 = (_zz_dataOut_payload_0_10012 < _zz_dataOut_payload_0_10060);
  assign _zz_dataOut_payload_0_10108 = (_zz_dataOut_payload_0_10107 ? _zz_dataOut_payload_0_10012 : _zz_dataOut_payload_0_10060);
  assign _zz_dataOut_payload_0_10109 = (_zz_dataOut_payload_0_10107 ? _zz_dataOut_payload_0_10060 : _zz_dataOut_payload_0_10012);
  assign _zz_dataOut_payload_0_10110 = (_zz_dataOut_payload_0_10015 < _zz_dataOut_payload_0_10063);
  assign _zz_dataOut_payload_0_10111 = (_zz_dataOut_payload_0_10110 ? _zz_dataOut_payload_0_10015 : _zz_dataOut_payload_0_10063);
  assign _zz_dataOut_payload_0_10112 = (_zz_dataOut_payload_0_10110 ? _zz_dataOut_payload_0_10063 : _zz_dataOut_payload_0_10015);
  assign _zz_dataOut_payload_0_10113 = (_zz_dataOut_payload_0_10018 < _zz_dataOut_payload_0_10066);
  assign _zz_dataOut_payload_0_10114 = (_zz_dataOut_payload_0_10113 ? _zz_dataOut_payload_0_10018 : _zz_dataOut_payload_0_10066);
  assign _zz_dataOut_payload_0_10115 = (_zz_dataOut_payload_0_10113 ? _zz_dataOut_payload_0_10066 : _zz_dataOut_payload_0_10018);
  assign _zz_dataOut_payload_0_10116 = (_zz_dataOut_payload_0_10021 < _zz_dataOut_payload_0_10069);
  assign _zz_dataOut_payload_0_10117 = (_zz_dataOut_payload_0_10116 ? _zz_dataOut_payload_0_10021 : _zz_dataOut_payload_0_10069);
  assign _zz_dataOut_payload_0_10118 = (_zz_dataOut_payload_0_10116 ? _zz_dataOut_payload_0_10069 : _zz_dataOut_payload_0_10021);
  assign _zz_dataOut_payload_0_10119 = (_zz_dataOut_payload_0_10024 < _zz_dataOut_payload_0_10072);
  assign _zz_dataOut_payload_0_10120 = (_zz_dataOut_payload_0_10119 ? _zz_dataOut_payload_0_10024 : _zz_dataOut_payload_0_10072);
  assign _zz_dataOut_payload_0_10121 = (_zz_dataOut_payload_0_10119 ? _zz_dataOut_payload_0_10072 : _zz_dataOut_payload_0_10024);
  assign _zz_dataOut_payload_0_10122 = (_zz_dataOut_payload_0_10027 < _zz_dataOut_payload_0_10075);
  assign _zz_dataOut_payload_0_10123 = (_zz_dataOut_payload_0_10122 ? _zz_dataOut_payload_0_10027 : _zz_dataOut_payload_0_10075);
  assign _zz_dataOut_payload_0_10124 = (_zz_dataOut_payload_0_10122 ? _zz_dataOut_payload_0_10075 : _zz_dataOut_payload_0_10027);
  assign _zz_dataOut_payload_0_10125 = (_zz_dataOut_payload_0_10030 < _zz_dataOut_payload_0_10078);
  assign _zz_dataOut_payload_0_10126 = (_zz_dataOut_payload_0_10125 ? _zz_dataOut_payload_0_10030 : _zz_dataOut_payload_0_10078);
  assign _zz_dataOut_payload_0_10127 = (_zz_dataOut_payload_0_10125 ? _zz_dataOut_payload_0_10078 : _zz_dataOut_payload_0_10030);
  assign _zz_dataOut_payload_0_10128 = (_zz_dataOut_payload_0_10081 < _zz_dataOut_payload_0_10105);
  assign _zz_dataOut_payload_0_10129 = (_zz_dataOut_payload_0_10128 ? _zz_dataOut_payload_0_10081 : _zz_dataOut_payload_0_10105);
  assign _zz_dataOut_payload_0_10130 = (_zz_dataOut_payload_0_10128 ? _zz_dataOut_payload_0_10105 : _zz_dataOut_payload_0_10081);
  assign _zz_dataOut_payload_0_10131 = (_zz_dataOut_payload_0_10084 < _zz_dataOut_payload_0_10108);
  assign _zz_dataOut_payload_0_10132 = (_zz_dataOut_payload_0_10131 ? _zz_dataOut_payload_0_10084 : _zz_dataOut_payload_0_10108);
  assign _zz_dataOut_payload_0_10133 = (_zz_dataOut_payload_0_10131 ? _zz_dataOut_payload_0_10108 : _zz_dataOut_payload_0_10084);
  assign _zz_dataOut_payload_0_10134 = (_zz_dataOut_payload_0_10087 < _zz_dataOut_payload_0_10111);
  assign _zz_dataOut_payload_0_10135 = (_zz_dataOut_payload_0_10134 ? _zz_dataOut_payload_0_10087 : _zz_dataOut_payload_0_10111);
  assign _zz_dataOut_payload_0_10136 = (_zz_dataOut_payload_0_10134 ? _zz_dataOut_payload_0_10111 : _zz_dataOut_payload_0_10087);
  assign _zz_dataOut_payload_0_10137 = (_zz_dataOut_payload_0_10090 < _zz_dataOut_payload_0_10114);
  assign _zz_dataOut_payload_0_10138 = (_zz_dataOut_payload_0_10137 ? _zz_dataOut_payload_0_10090 : _zz_dataOut_payload_0_10114);
  assign _zz_dataOut_payload_0_10139 = (_zz_dataOut_payload_0_10137 ? _zz_dataOut_payload_0_10114 : _zz_dataOut_payload_0_10090);
  assign _zz_dataOut_payload_0_10140 = (_zz_dataOut_payload_0_10093 < _zz_dataOut_payload_0_10117);
  assign _zz_dataOut_payload_0_10141 = (_zz_dataOut_payload_0_10140 ? _zz_dataOut_payload_0_10093 : _zz_dataOut_payload_0_10117);
  assign _zz_dataOut_payload_0_10142 = (_zz_dataOut_payload_0_10140 ? _zz_dataOut_payload_0_10117 : _zz_dataOut_payload_0_10093);
  assign _zz_dataOut_payload_0_10143 = (_zz_dataOut_payload_0_10096 < _zz_dataOut_payload_0_10120);
  assign _zz_dataOut_payload_0_10144 = (_zz_dataOut_payload_0_10143 ? _zz_dataOut_payload_0_10096 : _zz_dataOut_payload_0_10120);
  assign _zz_dataOut_payload_0_10145 = (_zz_dataOut_payload_0_10143 ? _zz_dataOut_payload_0_10120 : _zz_dataOut_payload_0_10096);
  assign _zz_dataOut_payload_0_10146 = (_zz_dataOut_payload_0_10099 < _zz_dataOut_payload_0_10123);
  assign _zz_dataOut_payload_0_10147 = (_zz_dataOut_payload_0_10146 ? _zz_dataOut_payload_0_10099 : _zz_dataOut_payload_0_10123);
  assign _zz_dataOut_payload_0_10148 = (_zz_dataOut_payload_0_10146 ? _zz_dataOut_payload_0_10123 : _zz_dataOut_payload_0_10099);
  assign _zz_dataOut_payload_0_10149 = (_zz_dataOut_payload_0_10102 < _zz_dataOut_payload_0_10126);
  assign _zz_dataOut_payload_0_10150 = (_zz_dataOut_payload_0_10149 ? _zz_dataOut_payload_0_10102 : _zz_dataOut_payload_0_10126);
  assign _zz_dataOut_payload_0_10151 = (_zz_dataOut_payload_0_10149 ? _zz_dataOut_payload_0_10126 : _zz_dataOut_payload_0_10102);
  assign _zz_dataOut_payload_0_10152 = (_zz_dataOut_payload_0_10129 < _zz_dataOut_payload_0_10141);
  assign _zz_dataOut_payload_0_10153 = (_zz_dataOut_payload_0_10152 ? _zz_dataOut_payload_0_10129 : _zz_dataOut_payload_0_10141);
  assign _zz_dataOut_payload_0_10154 = (_zz_dataOut_payload_0_10152 ? _zz_dataOut_payload_0_10141 : _zz_dataOut_payload_0_10129);
  assign _zz_dataOut_payload_0_10155 = (_zz_dataOut_payload_0_10132 < _zz_dataOut_payload_0_10144);
  assign _zz_dataOut_payload_0_10156 = (_zz_dataOut_payload_0_10155 ? _zz_dataOut_payload_0_10132 : _zz_dataOut_payload_0_10144);
  assign _zz_dataOut_payload_0_10157 = (_zz_dataOut_payload_0_10155 ? _zz_dataOut_payload_0_10144 : _zz_dataOut_payload_0_10132);
  assign _zz_dataOut_payload_0_10158 = (_zz_dataOut_payload_0_10135 < _zz_dataOut_payload_0_10147);
  assign _zz_dataOut_payload_0_10159 = (_zz_dataOut_payload_0_10158 ? _zz_dataOut_payload_0_10135 : _zz_dataOut_payload_0_10147);
  assign _zz_dataOut_payload_0_10160 = (_zz_dataOut_payload_0_10158 ? _zz_dataOut_payload_0_10147 : _zz_dataOut_payload_0_10135);
  assign _zz_dataOut_payload_0_10161 = (_zz_dataOut_payload_0_10138 < _zz_dataOut_payload_0_10150);
  assign _zz_dataOut_payload_0_10162 = (_zz_dataOut_payload_0_10161 ? _zz_dataOut_payload_0_10138 : _zz_dataOut_payload_0_10150);
  assign _zz_dataOut_payload_0_10163 = (_zz_dataOut_payload_0_10161 ? _zz_dataOut_payload_0_10150 : _zz_dataOut_payload_0_10138);
  assign _zz_dataOut_payload_0_10164 = (_zz_dataOut_payload_0_10153 < _zz_dataOut_payload_0_10159);
  assign _zz_dataOut_payload_0_10165 = (_zz_dataOut_payload_0_10164 ? _zz_dataOut_payload_0_10153 : _zz_dataOut_payload_0_10159);
  assign _zz_dataOut_payload_0_10166 = (_zz_dataOut_payload_0_10164 ? _zz_dataOut_payload_0_10159 : _zz_dataOut_payload_0_10153);
  assign _zz_dataOut_payload_0_10167 = (_zz_dataOut_payload_0_10156 < _zz_dataOut_payload_0_10162);
  assign _zz_dataOut_payload_0_10168 = (_zz_dataOut_payload_0_10167 ? _zz_dataOut_payload_0_10156 : _zz_dataOut_payload_0_10162);
  assign _zz_dataOut_payload_0_10169 = (_zz_dataOut_payload_0_10167 ? _zz_dataOut_payload_0_10162 : _zz_dataOut_payload_0_10156);
  assign _zz_dataOut_payload_0_10170 = (_zz_dataOut_payload_0_10165 < _zz_dataOut_payload_0_10168);
  assign _zz_dataOut_payload_0_10171 = (_zz_dataOut_payload_0_10166 < _zz_dataOut_payload_0_10169);
  assign _zz_dataOut_payload_0_10176 = (_zz_dataOut_payload_0_10154 < _zz_dataOut_payload_0_10160);
  assign _zz_dataOut_payload_0_10177 = (_zz_dataOut_payload_0_10176 ? _zz_dataOut_payload_0_10154 : _zz_dataOut_payload_0_10160);
  assign _zz_dataOut_payload_0_10178 = (_zz_dataOut_payload_0_10176 ? _zz_dataOut_payload_0_10160 : _zz_dataOut_payload_0_10154);
  assign _zz_dataOut_payload_0_10179 = (_zz_dataOut_payload_0_10157 < _zz_dataOut_payload_0_10163);
  assign _zz_dataOut_payload_0_10180 = (_zz_dataOut_payload_0_10179 ? _zz_dataOut_payload_0_10157 : _zz_dataOut_payload_0_10163);
  assign _zz_dataOut_payload_0_10181 = (_zz_dataOut_payload_0_10179 ? _zz_dataOut_payload_0_10163 : _zz_dataOut_payload_0_10157);
  assign _zz_dataOut_payload_0_10182 = (_zz_dataOut_payload_0_10177 < _zz_dataOut_payload_0_10180);
  assign _zz_dataOut_payload_0_10183 = (_zz_dataOut_payload_0_10178 < _zz_dataOut_payload_0_10181);
  assign _zz_dataOut_payload_0_10196 = (_zz_dataOut_payload_0_10130 < _zz_dataOut_payload_0_10142);
  assign _zz_dataOut_payload_0_10197 = (_zz_dataOut_payload_0_10196 ? _zz_dataOut_payload_0_10130 : _zz_dataOut_payload_0_10142);
  assign _zz_dataOut_payload_0_10198 = (_zz_dataOut_payload_0_10196 ? _zz_dataOut_payload_0_10142 : _zz_dataOut_payload_0_10130);
  assign _zz_dataOut_payload_0_10199 = (_zz_dataOut_payload_0_10133 < _zz_dataOut_payload_0_10145);
  assign _zz_dataOut_payload_0_10200 = (_zz_dataOut_payload_0_10199 ? _zz_dataOut_payload_0_10133 : _zz_dataOut_payload_0_10145);
  assign _zz_dataOut_payload_0_10201 = (_zz_dataOut_payload_0_10199 ? _zz_dataOut_payload_0_10145 : _zz_dataOut_payload_0_10133);
  assign _zz_dataOut_payload_0_10202 = (_zz_dataOut_payload_0_10136 < _zz_dataOut_payload_0_10148);
  assign _zz_dataOut_payload_0_10203 = (_zz_dataOut_payload_0_10202 ? _zz_dataOut_payload_0_10136 : _zz_dataOut_payload_0_10148);
  assign _zz_dataOut_payload_0_10204 = (_zz_dataOut_payload_0_10202 ? _zz_dataOut_payload_0_10148 : _zz_dataOut_payload_0_10136);
  assign _zz_dataOut_payload_0_10205 = (_zz_dataOut_payload_0_10139 < _zz_dataOut_payload_0_10151);
  assign _zz_dataOut_payload_0_10206 = (_zz_dataOut_payload_0_10205 ? _zz_dataOut_payload_0_10139 : _zz_dataOut_payload_0_10151);
  assign _zz_dataOut_payload_0_10207 = (_zz_dataOut_payload_0_10205 ? _zz_dataOut_payload_0_10151 : _zz_dataOut_payload_0_10139);
  assign _zz_dataOut_payload_0_10208 = (_zz_dataOut_payload_0_10197 < _zz_dataOut_payload_0_10203);
  assign _zz_dataOut_payload_0_10209 = (_zz_dataOut_payload_0_10208 ? _zz_dataOut_payload_0_10197 : _zz_dataOut_payload_0_10203);
  assign _zz_dataOut_payload_0_10210 = (_zz_dataOut_payload_0_10208 ? _zz_dataOut_payload_0_10203 : _zz_dataOut_payload_0_10197);
  assign _zz_dataOut_payload_0_10211 = (_zz_dataOut_payload_0_10200 < _zz_dataOut_payload_0_10206);
  assign _zz_dataOut_payload_0_10212 = (_zz_dataOut_payload_0_10211 ? _zz_dataOut_payload_0_10200 : _zz_dataOut_payload_0_10206);
  assign _zz_dataOut_payload_0_10213 = (_zz_dataOut_payload_0_10211 ? _zz_dataOut_payload_0_10206 : _zz_dataOut_payload_0_10200);
  assign _zz_dataOut_payload_0_10214 = (_zz_dataOut_payload_0_10209 < _zz_dataOut_payload_0_10212);
  assign _zz_dataOut_payload_0_10215 = (_zz_dataOut_payload_0_10210 < _zz_dataOut_payload_0_10213);
  assign _zz_dataOut_payload_0_10220 = (_zz_dataOut_payload_0_10198 < _zz_dataOut_payload_0_10204);
  assign _zz_dataOut_payload_0_10221 = (_zz_dataOut_payload_0_10220 ? _zz_dataOut_payload_0_10198 : _zz_dataOut_payload_0_10204);
  assign _zz_dataOut_payload_0_10222 = (_zz_dataOut_payload_0_10220 ? _zz_dataOut_payload_0_10204 : _zz_dataOut_payload_0_10198);
  assign _zz_dataOut_payload_0_10223 = (_zz_dataOut_payload_0_10201 < _zz_dataOut_payload_0_10207);
  assign _zz_dataOut_payload_0_10224 = (_zz_dataOut_payload_0_10223 ? _zz_dataOut_payload_0_10201 : _zz_dataOut_payload_0_10207);
  assign _zz_dataOut_payload_0_10225 = (_zz_dataOut_payload_0_10223 ? _zz_dataOut_payload_0_10207 : _zz_dataOut_payload_0_10201);
  assign _zz_dataOut_payload_0_10226 = (_zz_dataOut_payload_0_10221 < _zz_dataOut_payload_0_10224);
  assign _zz_dataOut_payload_0_10227 = (_zz_dataOut_payload_0_10222 < _zz_dataOut_payload_0_10225);
  assign _zz_dataOut_payload_0_10256 = (_zz_dataOut_payload_0_10082 < _zz_dataOut_payload_0_10106);
  assign _zz_dataOut_payload_0_10257 = (_zz_dataOut_payload_0_10256 ? _zz_dataOut_payload_0_10082 : _zz_dataOut_payload_0_10106);
  assign _zz_dataOut_payload_0_10258 = (_zz_dataOut_payload_0_10256 ? _zz_dataOut_payload_0_10106 : _zz_dataOut_payload_0_10082);
  assign _zz_dataOut_payload_0_10259 = (_zz_dataOut_payload_0_10085 < _zz_dataOut_payload_0_10109);
  assign _zz_dataOut_payload_0_10260 = (_zz_dataOut_payload_0_10259 ? _zz_dataOut_payload_0_10085 : _zz_dataOut_payload_0_10109);
  assign _zz_dataOut_payload_0_10261 = (_zz_dataOut_payload_0_10259 ? _zz_dataOut_payload_0_10109 : _zz_dataOut_payload_0_10085);
  assign _zz_dataOut_payload_0_10262 = (_zz_dataOut_payload_0_10088 < _zz_dataOut_payload_0_10112);
  assign _zz_dataOut_payload_0_10263 = (_zz_dataOut_payload_0_10262 ? _zz_dataOut_payload_0_10088 : _zz_dataOut_payload_0_10112);
  assign _zz_dataOut_payload_0_10264 = (_zz_dataOut_payload_0_10262 ? _zz_dataOut_payload_0_10112 : _zz_dataOut_payload_0_10088);
  assign _zz_dataOut_payload_0_10265 = (_zz_dataOut_payload_0_10091 < _zz_dataOut_payload_0_10115);
  assign _zz_dataOut_payload_0_10266 = (_zz_dataOut_payload_0_10265 ? _zz_dataOut_payload_0_10091 : _zz_dataOut_payload_0_10115);
  assign _zz_dataOut_payload_0_10267 = (_zz_dataOut_payload_0_10265 ? _zz_dataOut_payload_0_10115 : _zz_dataOut_payload_0_10091);
  assign _zz_dataOut_payload_0_10268 = (_zz_dataOut_payload_0_10094 < _zz_dataOut_payload_0_10118);
  assign _zz_dataOut_payload_0_10269 = (_zz_dataOut_payload_0_10268 ? _zz_dataOut_payload_0_10094 : _zz_dataOut_payload_0_10118);
  assign _zz_dataOut_payload_0_10270 = (_zz_dataOut_payload_0_10268 ? _zz_dataOut_payload_0_10118 : _zz_dataOut_payload_0_10094);
  assign _zz_dataOut_payload_0_10271 = (_zz_dataOut_payload_0_10097 < _zz_dataOut_payload_0_10121);
  assign _zz_dataOut_payload_0_10272 = (_zz_dataOut_payload_0_10271 ? _zz_dataOut_payload_0_10097 : _zz_dataOut_payload_0_10121);
  assign _zz_dataOut_payload_0_10273 = (_zz_dataOut_payload_0_10271 ? _zz_dataOut_payload_0_10121 : _zz_dataOut_payload_0_10097);
  assign _zz_dataOut_payload_0_10274 = (_zz_dataOut_payload_0_10100 < _zz_dataOut_payload_0_10124);
  assign _zz_dataOut_payload_0_10275 = (_zz_dataOut_payload_0_10274 ? _zz_dataOut_payload_0_10100 : _zz_dataOut_payload_0_10124);
  assign _zz_dataOut_payload_0_10276 = (_zz_dataOut_payload_0_10274 ? _zz_dataOut_payload_0_10124 : _zz_dataOut_payload_0_10100);
  assign _zz_dataOut_payload_0_10277 = (_zz_dataOut_payload_0_10103 < _zz_dataOut_payload_0_10127);
  assign _zz_dataOut_payload_0_10278 = (_zz_dataOut_payload_0_10277 ? _zz_dataOut_payload_0_10103 : _zz_dataOut_payload_0_10127);
  assign _zz_dataOut_payload_0_10279 = (_zz_dataOut_payload_0_10277 ? _zz_dataOut_payload_0_10127 : _zz_dataOut_payload_0_10103);
  assign _zz_dataOut_payload_0_10280 = (_zz_dataOut_payload_0_10257 < _zz_dataOut_payload_0_10269);
  assign _zz_dataOut_payload_0_10281 = (_zz_dataOut_payload_0_10280 ? _zz_dataOut_payload_0_10257 : _zz_dataOut_payload_0_10269);
  assign _zz_dataOut_payload_0_10282 = (_zz_dataOut_payload_0_10280 ? _zz_dataOut_payload_0_10269 : _zz_dataOut_payload_0_10257);
  assign _zz_dataOut_payload_0_10283 = (_zz_dataOut_payload_0_10260 < _zz_dataOut_payload_0_10272);
  assign _zz_dataOut_payload_0_10284 = (_zz_dataOut_payload_0_10283 ? _zz_dataOut_payload_0_10260 : _zz_dataOut_payload_0_10272);
  assign _zz_dataOut_payload_0_10285 = (_zz_dataOut_payload_0_10283 ? _zz_dataOut_payload_0_10272 : _zz_dataOut_payload_0_10260);
  assign _zz_dataOut_payload_0_10286 = (_zz_dataOut_payload_0_10263 < _zz_dataOut_payload_0_10275);
  assign _zz_dataOut_payload_0_10287 = (_zz_dataOut_payload_0_10286 ? _zz_dataOut_payload_0_10263 : _zz_dataOut_payload_0_10275);
  assign _zz_dataOut_payload_0_10288 = (_zz_dataOut_payload_0_10286 ? _zz_dataOut_payload_0_10275 : _zz_dataOut_payload_0_10263);
  assign _zz_dataOut_payload_0_10289 = (_zz_dataOut_payload_0_10266 < _zz_dataOut_payload_0_10278);
  assign _zz_dataOut_payload_0_10290 = (_zz_dataOut_payload_0_10289 ? _zz_dataOut_payload_0_10266 : _zz_dataOut_payload_0_10278);
  assign _zz_dataOut_payload_0_10291 = (_zz_dataOut_payload_0_10289 ? _zz_dataOut_payload_0_10278 : _zz_dataOut_payload_0_10266);
  assign _zz_dataOut_payload_0_10292 = (_zz_dataOut_payload_0_10281 < _zz_dataOut_payload_0_10287);
  assign _zz_dataOut_payload_0_10293 = (_zz_dataOut_payload_0_10292 ? _zz_dataOut_payload_0_10281 : _zz_dataOut_payload_0_10287);
  assign _zz_dataOut_payload_0_10294 = (_zz_dataOut_payload_0_10292 ? _zz_dataOut_payload_0_10287 : _zz_dataOut_payload_0_10281);
  assign _zz_dataOut_payload_0_10295 = (_zz_dataOut_payload_0_10284 < _zz_dataOut_payload_0_10290);
  assign _zz_dataOut_payload_0_10296 = (_zz_dataOut_payload_0_10295 ? _zz_dataOut_payload_0_10284 : _zz_dataOut_payload_0_10290);
  assign _zz_dataOut_payload_0_10297 = (_zz_dataOut_payload_0_10295 ? _zz_dataOut_payload_0_10290 : _zz_dataOut_payload_0_10284);
  assign _zz_dataOut_payload_0_10298 = (_zz_dataOut_payload_0_10293 < _zz_dataOut_payload_0_10296);
  assign _zz_dataOut_payload_0_10299 = (_zz_dataOut_payload_0_10294 < _zz_dataOut_payload_0_10297);
  assign _zz_dataOut_payload_0_10304 = (_zz_dataOut_payload_0_10282 < _zz_dataOut_payload_0_10288);
  assign _zz_dataOut_payload_0_10305 = (_zz_dataOut_payload_0_10304 ? _zz_dataOut_payload_0_10282 : _zz_dataOut_payload_0_10288);
  assign _zz_dataOut_payload_0_10306 = (_zz_dataOut_payload_0_10304 ? _zz_dataOut_payload_0_10288 : _zz_dataOut_payload_0_10282);
  assign _zz_dataOut_payload_0_10307 = (_zz_dataOut_payload_0_10285 < _zz_dataOut_payload_0_10291);
  assign _zz_dataOut_payload_0_10308 = (_zz_dataOut_payload_0_10307 ? _zz_dataOut_payload_0_10285 : _zz_dataOut_payload_0_10291);
  assign _zz_dataOut_payload_0_10309 = (_zz_dataOut_payload_0_10307 ? _zz_dataOut_payload_0_10291 : _zz_dataOut_payload_0_10285);
  assign _zz_dataOut_payload_0_10310 = (_zz_dataOut_payload_0_10305 < _zz_dataOut_payload_0_10308);
  assign _zz_dataOut_payload_0_10311 = (_zz_dataOut_payload_0_10306 < _zz_dataOut_payload_0_10309);
  assign _zz_dataOut_payload_0_10324 = (_zz_dataOut_payload_0_10258 < _zz_dataOut_payload_0_10270);
  assign _zz_dataOut_payload_0_10325 = (_zz_dataOut_payload_0_10324 ? _zz_dataOut_payload_0_10258 : _zz_dataOut_payload_0_10270);
  assign _zz_dataOut_payload_0_10326 = (_zz_dataOut_payload_0_10324 ? _zz_dataOut_payload_0_10270 : _zz_dataOut_payload_0_10258);
  assign _zz_dataOut_payload_0_10327 = (_zz_dataOut_payload_0_10261 < _zz_dataOut_payload_0_10273);
  assign _zz_dataOut_payload_0_10328 = (_zz_dataOut_payload_0_10327 ? _zz_dataOut_payload_0_10261 : _zz_dataOut_payload_0_10273);
  assign _zz_dataOut_payload_0_10329 = (_zz_dataOut_payload_0_10327 ? _zz_dataOut_payload_0_10273 : _zz_dataOut_payload_0_10261);
  assign _zz_dataOut_payload_0_10330 = (_zz_dataOut_payload_0_10264 < _zz_dataOut_payload_0_10276);
  assign _zz_dataOut_payload_0_10331 = (_zz_dataOut_payload_0_10330 ? _zz_dataOut_payload_0_10264 : _zz_dataOut_payload_0_10276);
  assign _zz_dataOut_payload_0_10332 = (_zz_dataOut_payload_0_10330 ? _zz_dataOut_payload_0_10276 : _zz_dataOut_payload_0_10264);
  assign _zz_dataOut_payload_0_10333 = (_zz_dataOut_payload_0_10267 < _zz_dataOut_payload_0_10279);
  assign _zz_dataOut_payload_0_10334 = (_zz_dataOut_payload_0_10333 ? _zz_dataOut_payload_0_10267 : _zz_dataOut_payload_0_10279);
  assign _zz_dataOut_payload_0_10335 = (_zz_dataOut_payload_0_10333 ? _zz_dataOut_payload_0_10279 : _zz_dataOut_payload_0_10267);
  assign _zz_dataOut_payload_0_10336 = (_zz_dataOut_payload_0_10325 < _zz_dataOut_payload_0_10331);
  assign _zz_dataOut_payload_0_10337 = (_zz_dataOut_payload_0_10336 ? _zz_dataOut_payload_0_10325 : _zz_dataOut_payload_0_10331);
  assign _zz_dataOut_payload_0_10338 = (_zz_dataOut_payload_0_10336 ? _zz_dataOut_payload_0_10331 : _zz_dataOut_payload_0_10325);
  assign _zz_dataOut_payload_0_10339 = (_zz_dataOut_payload_0_10328 < _zz_dataOut_payload_0_10334);
  assign _zz_dataOut_payload_0_10340 = (_zz_dataOut_payload_0_10339 ? _zz_dataOut_payload_0_10328 : _zz_dataOut_payload_0_10334);
  assign _zz_dataOut_payload_0_10341 = (_zz_dataOut_payload_0_10339 ? _zz_dataOut_payload_0_10334 : _zz_dataOut_payload_0_10328);
  assign _zz_dataOut_payload_0_10342 = (_zz_dataOut_payload_0_10337 < _zz_dataOut_payload_0_10340);
  assign _zz_dataOut_payload_0_10343 = (_zz_dataOut_payload_0_10338 < _zz_dataOut_payload_0_10341);
  assign _zz_dataOut_payload_0_10348 = (_zz_dataOut_payload_0_10326 < _zz_dataOut_payload_0_10332);
  assign _zz_dataOut_payload_0_10349 = (_zz_dataOut_payload_0_10348 ? _zz_dataOut_payload_0_10326 : _zz_dataOut_payload_0_10332);
  assign _zz_dataOut_payload_0_10350 = (_zz_dataOut_payload_0_10348 ? _zz_dataOut_payload_0_10332 : _zz_dataOut_payload_0_10326);
  assign _zz_dataOut_payload_0_10351 = (_zz_dataOut_payload_0_10329 < _zz_dataOut_payload_0_10335);
  assign _zz_dataOut_payload_0_10352 = (_zz_dataOut_payload_0_10351 ? _zz_dataOut_payload_0_10329 : _zz_dataOut_payload_0_10335);
  assign _zz_dataOut_payload_0_10353 = (_zz_dataOut_payload_0_10351 ? _zz_dataOut_payload_0_10335 : _zz_dataOut_payload_0_10329);
  assign _zz_dataOut_payload_0_10354 = (_zz_dataOut_payload_0_10349 < _zz_dataOut_payload_0_10352);
  assign _zz_dataOut_payload_0_10355 = (_zz_dataOut_payload_0_10350 < _zz_dataOut_payload_0_10353);
  assign _zz_dataOut_payload_0_10416 = (_zz_dataOut_payload_0_10079 < _zz_dataOut_payload_0_10031);
  assign _zz_dataOut_payload_0_10417 = (_zz_dataOut_payload_0_10416 ? _zz_dataOut_payload_0_10079 : _zz_dataOut_payload_0_10031);
  assign _zz_dataOut_payload_0_10418 = (_zz_dataOut_payload_0_10416 ? _zz_dataOut_payload_0_10031 : _zz_dataOut_payload_0_10079);
  assign _zz_dataOut_payload_0_10419 = (_zz_dataOut_payload_0_10076 < _zz_dataOut_payload_0_10028);
  assign _zz_dataOut_payload_0_10420 = (_zz_dataOut_payload_0_10419 ? _zz_dataOut_payload_0_10076 : _zz_dataOut_payload_0_10028);
  assign _zz_dataOut_payload_0_10421 = (_zz_dataOut_payload_0_10419 ? _zz_dataOut_payload_0_10028 : _zz_dataOut_payload_0_10076);
  assign _zz_dataOut_payload_0_10422 = (_zz_dataOut_payload_0_10073 < _zz_dataOut_payload_0_10025);
  assign _zz_dataOut_payload_0_10423 = (_zz_dataOut_payload_0_10422 ? _zz_dataOut_payload_0_10073 : _zz_dataOut_payload_0_10025);
  assign _zz_dataOut_payload_0_10424 = (_zz_dataOut_payload_0_10422 ? _zz_dataOut_payload_0_10025 : _zz_dataOut_payload_0_10073);
  assign _zz_dataOut_payload_0_10425 = (_zz_dataOut_payload_0_10070 < _zz_dataOut_payload_0_10022);
  assign _zz_dataOut_payload_0_10426 = (_zz_dataOut_payload_0_10425 ? _zz_dataOut_payload_0_10070 : _zz_dataOut_payload_0_10022);
  assign _zz_dataOut_payload_0_10427 = (_zz_dataOut_payload_0_10425 ? _zz_dataOut_payload_0_10022 : _zz_dataOut_payload_0_10070);
  assign _zz_dataOut_payload_0_10428 = (_zz_dataOut_payload_0_10067 < _zz_dataOut_payload_0_10019);
  assign _zz_dataOut_payload_0_10429 = (_zz_dataOut_payload_0_10428 ? _zz_dataOut_payload_0_10067 : _zz_dataOut_payload_0_10019);
  assign _zz_dataOut_payload_0_10430 = (_zz_dataOut_payload_0_10428 ? _zz_dataOut_payload_0_10019 : _zz_dataOut_payload_0_10067);
  assign _zz_dataOut_payload_0_10431 = (_zz_dataOut_payload_0_10064 < _zz_dataOut_payload_0_10016);
  assign _zz_dataOut_payload_0_10432 = (_zz_dataOut_payload_0_10431 ? _zz_dataOut_payload_0_10064 : _zz_dataOut_payload_0_10016);
  assign _zz_dataOut_payload_0_10433 = (_zz_dataOut_payload_0_10431 ? _zz_dataOut_payload_0_10016 : _zz_dataOut_payload_0_10064);
  assign _zz_dataOut_payload_0_10434 = (_zz_dataOut_payload_0_10061 < _zz_dataOut_payload_0_10013);
  assign _zz_dataOut_payload_0_10435 = (_zz_dataOut_payload_0_10434 ? _zz_dataOut_payload_0_10061 : _zz_dataOut_payload_0_10013);
  assign _zz_dataOut_payload_0_10436 = (_zz_dataOut_payload_0_10434 ? _zz_dataOut_payload_0_10013 : _zz_dataOut_payload_0_10061);
  assign _zz_dataOut_payload_0_10437 = (_zz_dataOut_payload_0_10058 < _zz_dataOut_payload_0_10010);
  assign _zz_dataOut_payload_0_10438 = (_zz_dataOut_payload_0_10437 ? _zz_dataOut_payload_0_10058 : _zz_dataOut_payload_0_10010);
  assign _zz_dataOut_payload_0_10439 = (_zz_dataOut_payload_0_10437 ? _zz_dataOut_payload_0_10010 : _zz_dataOut_payload_0_10058);
  assign _zz_dataOut_payload_0_10440 = (_zz_dataOut_payload_0_10055 < _zz_dataOut_payload_0_10007);
  assign _zz_dataOut_payload_0_10441 = (_zz_dataOut_payload_0_10440 ? _zz_dataOut_payload_0_10055 : _zz_dataOut_payload_0_10007);
  assign _zz_dataOut_payload_0_10442 = (_zz_dataOut_payload_0_10440 ? _zz_dataOut_payload_0_10007 : _zz_dataOut_payload_0_10055);
  assign _zz_dataOut_payload_0_10443 = (_zz_dataOut_payload_0_10052 < _zz_dataOut_payload_0_10004);
  assign _zz_dataOut_payload_0_10444 = (_zz_dataOut_payload_0_10443 ? _zz_dataOut_payload_0_10052 : _zz_dataOut_payload_0_10004);
  assign _zz_dataOut_payload_0_10445 = (_zz_dataOut_payload_0_10443 ? _zz_dataOut_payload_0_10004 : _zz_dataOut_payload_0_10052);
  assign _zz_dataOut_payload_0_10446 = (_zz_dataOut_payload_0_10049 < _zz_dataOut_payload_0_10001);
  assign _zz_dataOut_payload_0_10447 = (_zz_dataOut_payload_0_10446 ? _zz_dataOut_payload_0_10049 : _zz_dataOut_payload_0_10001);
  assign _zz_dataOut_payload_0_10448 = (_zz_dataOut_payload_0_10446 ? _zz_dataOut_payload_0_10001 : _zz_dataOut_payload_0_10049);
  assign _zz_dataOut_payload_0_10449 = (_zz_dataOut_payload_0_10046 < _zz_dataOut_payload_0_9998);
  assign _zz_dataOut_payload_0_10450 = (_zz_dataOut_payload_0_10449 ? _zz_dataOut_payload_0_10046 : _zz_dataOut_payload_0_9998);
  assign _zz_dataOut_payload_0_10451 = (_zz_dataOut_payload_0_10449 ? _zz_dataOut_payload_0_9998 : _zz_dataOut_payload_0_10046);
  assign _zz_dataOut_payload_0_10452 = (_zz_dataOut_payload_0_10043 < _zz_dataOut_payload_0_9995);
  assign _zz_dataOut_payload_0_10453 = (_zz_dataOut_payload_0_10452 ? _zz_dataOut_payload_0_10043 : _zz_dataOut_payload_0_9995);
  assign _zz_dataOut_payload_0_10454 = (_zz_dataOut_payload_0_10452 ? _zz_dataOut_payload_0_9995 : _zz_dataOut_payload_0_10043);
  assign _zz_dataOut_payload_0_10455 = (_zz_dataOut_payload_0_10040 < _zz_dataOut_payload_0_9992);
  assign _zz_dataOut_payload_0_10456 = (_zz_dataOut_payload_0_10455 ? _zz_dataOut_payload_0_10040 : _zz_dataOut_payload_0_9992);
  assign _zz_dataOut_payload_0_10457 = (_zz_dataOut_payload_0_10455 ? _zz_dataOut_payload_0_9992 : _zz_dataOut_payload_0_10040);
  assign _zz_dataOut_payload_0_10458 = (_zz_dataOut_payload_0_10037 < _zz_dataOut_payload_0_9989);
  assign _zz_dataOut_payload_0_10459 = (_zz_dataOut_payload_0_10458 ? _zz_dataOut_payload_0_10037 : _zz_dataOut_payload_0_9989);
  assign _zz_dataOut_payload_0_10460 = (_zz_dataOut_payload_0_10458 ? _zz_dataOut_payload_0_9989 : _zz_dataOut_payload_0_10037);
  assign _zz_dataOut_payload_0_10461 = (_zz_dataOut_payload_0_10034 < _zz_dataOut_payload_0_9986);
  assign _zz_dataOut_payload_0_10462 = (_zz_dataOut_payload_0_10461 ? _zz_dataOut_payload_0_10034 : _zz_dataOut_payload_0_9986);
  assign _zz_dataOut_payload_0_10463 = (_zz_dataOut_payload_0_10461 ? _zz_dataOut_payload_0_9986 : _zz_dataOut_payload_0_10034);
  assign _zz_dataOut_payload_0_10464 = (_zz_dataOut_payload_0_10417 < _zz_dataOut_payload_0_10441);
  assign _zz_dataOut_payload_0_10465 = (_zz_dataOut_payload_0_10464 ? _zz_dataOut_payload_0_10417 : _zz_dataOut_payload_0_10441);
  assign _zz_dataOut_payload_0_10466 = (_zz_dataOut_payload_0_10464 ? _zz_dataOut_payload_0_10441 : _zz_dataOut_payload_0_10417);
  assign _zz_dataOut_payload_0_10467 = (_zz_dataOut_payload_0_10420 < _zz_dataOut_payload_0_10444);
  assign _zz_dataOut_payload_0_10468 = (_zz_dataOut_payload_0_10467 ? _zz_dataOut_payload_0_10420 : _zz_dataOut_payload_0_10444);
  assign _zz_dataOut_payload_0_10469 = (_zz_dataOut_payload_0_10467 ? _zz_dataOut_payload_0_10444 : _zz_dataOut_payload_0_10420);
  assign _zz_dataOut_payload_0_10470 = (_zz_dataOut_payload_0_10423 < _zz_dataOut_payload_0_10447);
  assign _zz_dataOut_payload_0_10471 = (_zz_dataOut_payload_0_10470 ? _zz_dataOut_payload_0_10423 : _zz_dataOut_payload_0_10447);
  assign _zz_dataOut_payload_0_10472 = (_zz_dataOut_payload_0_10470 ? _zz_dataOut_payload_0_10447 : _zz_dataOut_payload_0_10423);
  assign _zz_dataOut_payload_0_10473 = (_zz_dataOut_payload_0_10426 < _zz_dataOut_payload_0_10450);
  assign _zz_dataOut_payload_0_10474 = (_zz_dataOut_payload_0_10473 ? _zz_dataOut_payload_0_10426 : _zz_dataOut_payload_0_10450);
  assign _zz_dataOut_payload_0_10475 = (_zz_dataOut_payload_0_10473 ? _zz_dataOut_payload_0_10450 : _zz_dataOut_payload_0_10426);
  assign _zz_dataOut_payload_0_10476 = (_zz_dataOut_payload_0_10429 < _zz_dataOut_payload_0_10453);
  assign _zz_dataOut_payload_0_10477 = (_zz_dataOut_payload_0_10476 ? _zz_dataOut_payload_0_10429 : _zz_dataOut_payload_0_10453);
  assign _zz_dataOut_payload_0_10478 = (_zz_dataOut_payload_0_10476 ? _zz_dataOut_payload_0_10453 : _zz_dataOut_payload_0_10429);
  assign _zz_dataOut_payload_0_10479 = (_zz_dataOut_payload_0_10432 < _zz_dataOut_payload_0_10456);
  assign _zz_dataOut_payload_0_10480 = (_zz_dataOut_payload_0_10479 ? _zz_dataOut_payload_0_10432 : _zz_dataOut_payload_0_10456);
  assign _zz_dataOut_payload_0_10481 = (_zz_dataOut_payload_0_10479 ? _zz_dataOut_payload_0_10456 : _zz_dataOut_payload_0_10432);
  assign _zz_dataOut_payload_0_10482 = (_zz_dataOut_payload_0_10435 < _zz_dataOut_payload_0_10459);
  assign _zz_dataOut_payload_0_10483 = (_zz_dataOut_payload_0_10482 ? _zz_dataOut_payload_0_10435 : _zz_dataOut_payload_0_10459);
  assign _zz_dataOut_payload_0_10484 = (_zz_dataOut_payload_0_10482 ? _zz_dataOut_payload_0_10459 : _zz_dataOut_payload_0_10435);
  assign _zz_dataOut_payload_0_10485 = (_zz_dataOut_payload_0_10438 < _zz_dataOut_payload_0_10462);
  assign _zz_dataOut_payload_0_10486 = (_zz_dataOut_payload_0_10485 ? _zz_dataOut_payload_0_10438 : _zz_dataOut_payload_0_10462);
  assign _zz_dataOut_payload_0_10487 = (_zz_dataOut_payload_0_10485 ? _zz_dataOut_payload_0_10462 : _zz_dataOut_payload_0_10438);
  assign _zz_dataOut_payload_0_10488 = (_zz_dataOut_payload_0_10465 < _zz_dataOut_payload_0_10477);
  assign _zz_dataOut_payload_0_10489 = (_zz_dataOut_payload_0_10488 ? _zz_dataOut_payload_0_10465 : _zz_dataOut_payload_0_10477);
  assign _zz_dataOut_payload_0_10490 = (_zz_dataOut_payload_0_10488 ? _zz_dataOut_payload_0_10477 : _zz_dataOut_payload_0_10465);
  assign _zz_dataOut_payload_0_10491 = (_zz_dataOut_payload_0_10468 < _zz_dataOut_payload_0_10480);
  assign _zz_dataOut_payload_0_10492 = (_zz_dataOut_payload_0_10491 ? _zz_dataOut_payload_0_10468 : _zz_dataOut_payload_0_10480);
  assign _zz_dataOut_payload_0_10493 = (_zz_dataOut_payload_0_10491 ? _zz_dataOut_payload_0_10480 : _zz_dataOut_payload_0_10468);
  assign _zz_dataOut_payload_0_10494 = (_zz_dataOut_payload_0_10471 < _zz_dataOut_payload_0_10483);
  assign _zz_dataOut_payload_0_10495 = (_zz_dataOut_payload_0_10494 ? _zz_dataOut_payload_0_10471 : _zz_dataOut_payload_0_10483);
  assign _zz_dataOut_payload_0_10496 = (_zz_dataOut_payload_0_10494 ? _zz_dataOut_payload_0_10483 : _zz_dataOut_payload_0_10471);
  assign _zz_dataOut_payload_0_10497 = (_zz_dataOut_payload_0_10474 < _zz_dataOut_payload_0_10486);
  assign _zz_dataOut_payload_0_10498 = (_zz_dataOut_payload_0_10497 ? _zz_dataOut_payload_0_10474 : _zz_dataOut_payload_0_10486);
  assign _zz_dataOut_payload_0_10499 = (_zz_dataOut_payload_0_10497 ? _zz_dataOut_payload_0_10486 : _zz_dataOut_payload_0_10474);
  assign _zz_dataOut_payload_0_10500 = (_zz_dataOut_payload_0_10489 < _zz_dataOut_payload_0_10495);
  assign _zz_dataOut_payload_0_10501 = (_zz_dataOut_payload_0_10500 ? _zz_dataOut_payload_0_10489 : _zz_dataOut_payload_0_10495);
  assign _zz_dataOut_payload_0_10502 = (_zz_dataOut_payload_0_10500 ? _zz_dataOut_payload_0_10495 : _zz_dataOut_payload_0_10489);
  assign _zz_dataOut_payload_0_10503 = (_zz_dataOut_payload_0_10492 < _zz_dataOut_payload_0_10498);
  assign _zz_dataOut_payload_0_10504 = (_zz_dataOut_payload_0_10503 ? _zz_dataOut_payload_0_10492 : _zz_dataOut_payload_0_10498);
  assign _zz_dataOut_payload_0_10505 = (_zz_dataOut_payload_0_10503 ? _zz_dataOut_payload_0_10498 : _zz_dataOut_payload_0_10492);
  assign _zz_dataOut_payload_0_10506 = (_zz_dataOut_payload_0_10501 < _zz_dataOut_payload_0_10504);
  assign _zz_dataOut_payload_0_10507 = (_zz_dataOut_payload_0_10502 < _zz_dataOut_payload_0_10505);
  assign _zz_dataOut_payload_0_10512 = (_zz_dataOut_payload_0_10490 < _zz_dataOut_payload_0_10496);
  assign _zz_dataOut_payload_0_10513 = (_zz_dataOut_payload_0_10512 ? _zz_dataOut_payload_0_10490 : _zz_dataOut_payload_0_10496);
  assign _zz_dataOut_payload_0_10514 = (_zz_dataOut_payload_0_10512 ? _zz_dataOut_payload_0_10496 : _zz_dataOut_payload_0_10490);
  assign _zz_dataOut_payload_0_10515 = (_zz_dataOut_payload_0_10493 < _zz_dataOut_payload_0_10499);
  assign _zz_dataOut_payload_0_10516 = (_zz_dataOut_payload_0_10515 ? _zz_dataOut_payload_0_10493 : _zz_dataOut_payload_0_10499);
  assign _zz_dataOut_payload_0_10517 = (_zz_dataOut_payload_0_10515 ? _zz_dataOut_payload_0_10499 : _zz_dataOut_payload_0_10493);
  assign _zz_dataOut_payload_0_10518 = (_zz_dataOut_payload_0_10513 < _zz_dataOut_payload_0_10516);
  assign _zz_dataOut_payload_0_10519 = (_zz_dataOut_payload_0_10514 < _zz_dataOut_payload_0_10517);
  assign _zz_dataOut_payload_0_10532 = (_zz_dataOut_payload_0_10466 < _zz_dataOut_payload_0_10478);
  assign _zz_dataOut_payload_0_10533 = (_zz_dataOut_payload_0_10532 ? _zz_dataOut_payload_0_10466 : _zz_dataOut_payload_0_10478);
  assign _zz_dataOut_payload_0_10534 = (_zz_dataOut_payload_0_10532 ? _zz_dataOut_payload_0_10478 : _zz_dataOut_payload_0_10466);
  assign _zz_dataOut_payload_0_10535 = (_zz_dataOut_payload_0_10469 < _zz_dataOut_payload_0_10481);
  assign _zz_dataOut_payload_0_10536 = (_zz_dataOut_payload_0_10535 ? _zz_dataOut_payload_0_10469 : _zz_dataOut_payload_0_10481);
  assign _zz_dataOut_payload_0_10537 = (_zz_dataOut_payload_0_10535 ? _zz_dataOut_payload_0_10481 : _zz_dataOut_payload_0_10469);
  assign _zz_dataOut_payload_0_10538 = (_zz_dataOut_payload_0_10472 < _zz_dataOut_payload_0_10484);
  assign _zz_dataOut_payload_0_10539 = (_zz_dataOut_payload_0_10538 ? _zz_dataOut_payload_0_10472 : _zz_dataOut_payload_0_10484);
  assign _zz_dataOut_payload_0_10540 = (_zz_dataOut_payload_0_10538 ? _zz_dataOut_payload_0_10484 : _zz_dataOut_payload_0_10472);
  assign _zz_dataOut_payload_0_10541 = (_zz_dataOut_payload_0_10475 < _zz_dataOut_payload_0_10487);
  assign _zz_dataOut_payload_0_10542 = (_zz_dataOut_payload_0_10541 ? _zz_dataOut_payload_0_10475 : _zz_dataOut_payload_0_10487);
  assign _zz_dataOut_payload_0_10543 = (_zz_dataOut_payload_0_10541 ? _zz_dataOut_payload_0_10487 : _zz_dataOut_payload_0_10475);
  assign _zz_dataOut_payload_0_10544 = (_zz_dataOut_payload_0_10533 < _zz_dataOut_payload_0_10539);
  assign _zz_dataOut_payload_0_10545 = (_zz_dataOut_payload_0_10544 ? _zz_dataOut_payload_0_10533 : _zz_dataOut_payload_0_10539);
  assign _zz_dataOut_payload_0_10546 = (_zz_dataOut_payload_0_10544 ? _zz_dataOut_payload_0_10539 : _zz_dataOut_payload_0_10533);
  assign _zz_dataOut_payload_0_10547 = (_zz_dataOut_payload_0_10536 < _zz_dataOut_payload_0_10542);
  assign _zz_dataOut_payload_0_10548 = (_zz_dataOut_payload_0_10547 ? _zz_dataOut_payload_0_10536 : _zz_dataOut_payload_0_10542);
  assign _zz_dataOut_payload_0_10549 = (_zz_dataOut_payload_0_10547 ? _zz_dataOut_payload_0_10542 : _zz_dataOut_payload_0_10536);
  assign _zz_dataOut_payload_0_10550 = (_zz_dataOut_payload_0_10545 < _zz_dataOut_payload_0_10548);
  assign _zz_dataOut_payload_0_10551 = (_zz_dataOut_payload_0_10546 < _zz_dataOut_payload_0_10549);
  assign _zz_dataOut_payload_0_10556 = (_zz_dataOut_payload_0_10534 < _zz_dataOut_payload_0_10540);
  assign _zz_dataOut_payload_0_10557 = (_zz_dataOut_payload_0_10556 ? _zz_dataOut_payload_0_10534 : _zz_dataOut_payload_0_10540);
  assign _zz_dataOut_payload_0_10558 = (_zz_dataOut_payload_0_10556 ? _zz_dataOut_payload_0_10540 : _zz_dataOut_payload_0_10534);
  assign _zz_dataOut_payload_0_10559 = (_zz_dataOut_payload_0_10537 < _zz_dataOut_payload_0_10543);
  assign _zz_dataOut_payload_0_10560 = (_zz_dataOut_payload_0_10559 ? _zz_dataOut_payload_0_10537 : _zz_dataOut_payload_0_10543);
  assign _zz_dataOut_payload_0_10561 = (_zz_dataOut_payload_0_10559 ? _zz_dataOut_payload_0_10543 : _zz_dataOut_payload_0_10537);
  assign _zz_dataOut_payload_0_10562 = (_zz_dataOut_payload_0_10557 < _zz_dataOut_payload_0_10560);
  assign _zz_dataOut_payload_0_10563 = (_zz_dataOut_payload_0_10558 < _zz_dataOut_payload_0_10561);
  assign _zz_dataOut_payload_0_10592 = (_zz_dataOut_payload_0_10418 < _zz_dataOut_payload_0_10442);
  assign _zz_dataOut_payload_0_10593 = (_zz_dataOut_payload_0_10592 ? _zz_dataOut_payload_0_10418 : _zz_dataOut_payload_0_10442);
  assign _zz_dataOut_payload_0_10594 = (_zz_dataOut_payload_0_10592 ? _zz_dataOut_payload_0_10442 : _zz_dataOut_payload_0_10418);
  assign _zz_dataOut_payload_0_10595 = (_zz_dataOut_payload_0_10421 < _zz_dataOut_payload_0_10445);
  assign _zz_dataOut_payload_0_10596 = (_zz_dataOut_payload_0_10595 ? _zz_dataOut_payload_0_10421 : _zz_dataOut_payload_0_10445);
  assign _zz_dataOut_payload_0_10597 = (_zz_dataOut_payload_0_10595 ? _zz_dataOut_payload_0_10445 : _zz_dataOut_payload_0_10421);
  assign _zz_dataOut_payload_0_10598 = (_zz_dataOut_payload_0_10424 < _zz_dataOut_payload_0_10448);
  assign _zz_dataOut_payload_0_10599 = (_zz_dataOut_payload_0_10598 ? _zz_dataOut_payload_0_10424 : _zz_dataOut_payload_0_10448);
  assign _zz_dataOut_payload_0_10600 = (_zz_dataOut_payload_0_10598 ? _zz_dataOut_payload_0_10448 : _zz_dataOut_payload_0_10424);
  assign _zz_dataOut_payload_0_10601 = (_zz_dataOut_payload_0_10427 < _zz_dataOut_payload_0_10451);
  assign _zz_dataOut_payload_0_10602 = (_zz_dataOut_payload_0_10601 ? _zz_dataOut_payload_0_10427 : _zz_dataOut_payload_0_10451);
  assign _zz_dataOut_payload_0_10603 = (_zz_dataOut_payload_0_10601 ? _zz_dataOut_payload_0_10451 : _zz_dataOut_payload_0_10427);
  assign _zz_dataOut_payload_0_10604 = (_zz_dataOut_payload_0_10430 < _zz_dataOut_payload_0_10454);
  assign _zz_dataOut_payload_0_10605 = (_zz_dataOut_payload_0_10604 ? _zz_dataOut_payload_0_10430 : _zz_dataOut_payload_0_10454);
  assign _zz_dataOut_payload_0_10606 = (_zz_dataOut_payload_0_10604 ? _zz_dataOut_payload_0_10454 : _zz_dataOut_payload_0_10430);
  assign _zz_dataOut_payload_0_10607 = (_zz_dataOut_payload_0_10433 < _zz_dataOut_payload_0_10457);
  assign _zz_dataOut_payload_0_10608 = (_zz_dataOut_payload_0_10607 ? _zz_dataOut_payload_0_10433 : _zz_dataOut_payload_0_10457);
  assign _zz_dataOut_payload_0_10609 = (_zz_dataOut_payload_0_10607 ? _zz_dataOut_payload_0_10457 : _zz_dataOut_payload_0_10433);
  assign _zz_dataOut_payload_0_10610 = (_zz_dataOut_payload_0_10436 < _zz_dataOut_payload_0_10460);
  assign _zz_dataOut_payload_0_10611 = (_zz_dataOut_payload_0_10610 ? _zz_dataOut_payload_0_10436 : _zz_dataOut_payload_0_10460);
  assign _zz_dataOut_payload_0_10612 = (_zz_dataOut_payload_0_10610 ? _zz_dataOut_payload_0_10460 : _zz_dataOut_payload_0_10436);
  assign _zz_dataOut_payload_0_10613 = (_zz_dataOut_payload_0_10439 < _zz_dataOut_payload_0_10463);
  assign _zz_dataOut_payload_0_10614 = (_zz_dataOut_payload_0_10613 ? _zz_dataOut_payload_0_10439 : _zz_dataOut_payload_0_10463);
  assign _zz_dataOut_payload_0_10615 = (_zz_dataOut_payload_0_10613 ? _zz_dataOut_payload_0_10463 : _zz_dataOut_payload_0_10439);
  assign _zz_dataOut_payload_0_10616 = (_zz_dataOut_payload_0_10593 < _zz_dataOut_payload_0_10605);
  assign _zz_dataOut_payload_0_10617 = (_zz_dataOut_payload_0_10616 ? _zz_dataOut_payload_0_10593 : _zz_dataOut_payload_0_10605);
  assign _zz_dataOut_payload_0_10618 = (_zz_dataOut_payload_0_10616 ? _zz_dataOut_payload_0_10605 : _zz_dataOut_payload_0_10593);
  assign _zz_dataOut_payload_0_10619 = (_zz_dataOut_payload_0_10596 < _zz_dataOut_payload_0_10608);
  assign _zz_dataOut_payload_0_10620 = (_zz_dataOut_payload_0_10619 ? _zz_dataOut_payload_0_10596 : _zz_dataOut_payload_0_10608);
  assign _zz_dataOut_payload_0_10621 = (_zz_dataOut_payload_0_10619 ? _zz_dataOut_payload_0_10608 : _zz_dataOut_payload_0_10596);
  assign _zz_dataOut_payload_0_10622 = (_zz_dataOut_payload_0_10599 < _zz_dataOut_payload_0_10611);
  assign _zz_dataOut_payload_0_10623 = (_zz_dataOut_payload_0_10622 ? _zz_dataOut_payload_0_10599 : _zz_dataOut_payload_0_10611);
  assign _zz_dataOut_payload_0_10624 = (_zz_dataOut_payload_0_10622 ? _zz_dataOut_payload_0_10611 : _zz_dataOut_payload_0_10599);
  assign _zz_dataOut_payload_0_10625 = (_zz_dataOut_payload_0_10602 < _zz_dataOut_payload_0_10614);
  assign _zz_dataOut_payload_0_10626 = (_zz_dataOut_payload_0_10625 ? _zz_dataOut_payload_0_10602 : _zz_dataOut_payload_0_10614);
  assign _zz_dataOut_payload_0_10627 = (_zz_dataOut_payload_0_10625 ? _zz_dataOut_payload_0_10614 : _zz_dataOut_payload_0_10602);
  assign _zz_dataOut_payload_0_10628 = (_zz_dataOut_payload_0_10617 < _zz_dataOut_payload_0_10623);
  assign _zz_dataOut_payload_0_10629 = (_zz_dataOut_payload_0_10628 ? _zz_dataOut_payload_0_10617 : _zz_dataOut_payload_0_10623);
  assign _zz_dataOut_payload_0_10630 = (_zz_dataOut_payload_0_10628 ? _zz_dataOut_payload_0_10623 : _zz_dataOut_payload_0_10617);
  assign _zz_dataOut_payload_0_10631 = (_zz_dataOut_payload_0_10620 < _zz_dataOut_payload_0_10626);
  assign _zz_dataOut_payload_0_10632 = (_zz_dataOut_payload_0_10631 ? _zz_dataOut_payload_0_10620 : _zz_dataOut_payload_0_10626);
  assign _zz_dataOut_payload_0_10633 = (_zz_dataOut_payload_0_10631 ? _zz_dataOut_payload_0_10626 : _zz_dataOut_payload_0_10620);
  assign _zz_dataOut_payload_0_10634 = (_zz_dataOut_payload_0_10629 < _zz_dataOut_payload_0_10632);
  assign _zz_dataOut_payload_0_10635 = (_zz_dataOut_payload_0_10630 < _zz_dataOut_payload_0_10633);
  assign _zz_dataOut_payload_0_10640 = (_zz_dataOut_payload_0_10618 < _zz_dataOut_payload_0_10624);
  assign _zz_dataOut_payload_0_10641 = (_zz_dataOut_payload_0_10640 ? _zz_dataOut_payload_0_10618 : _zz_dataOut_payload_0_10624);
  assign _zz_dataOut_payload_0_10642 = (_zz_dataOut_payload_0_10640 ? _zz_dataOut_payload_0_10624 : _zz_dataOut_payload_0_10618);
  assign _zz_dataOut_payload_0_10643 = (_zz_dataOut_payload_0_10621 < _zz_dataOut_payload_0_10627);
  assign _zz_dataOut_payload_0_10644 = (_zz_dataOut_payload_0_10643 ? _zz_dataOut_payload_0_10621 : _zz_dataOut_payload_0_10627);
  assign _zz_dataOut_payload_0_10645 = (_zz_dataOut_payload_0_10643 ? _zz_dataOut_payload_0_10627 : _zz_dataOut_payload_0_10621);
  assign _zz_dataOut_payload_0_10646 = (_zz_dataOut_payload_0_10641 < _zz_dataOut_payload_0_10644);
  assign _zz_dataOut_payload_0_10647 = (_zz_dataOut_payload_0_10642 < _zz_dataOut_payload_0_10645);
  assign _zz_dataOut_payload_0_10660 = (_zz_dataOut_payload_0_10594 < _zz_dataOut_payload_0_10606);
  assign _zz_dataOut_payload_0_10661 = (_zz_dataOut_payload_0_10660 ? _zz_dataOut_payload_0_10594 : _zz_dataOut_payload_0_10606);
  assign _zz_dataOut_payload_0_10662 = (_zz_dataOut_payload_0_10660 ? _zz_dataOut_payload_0_10606 : _zz_dataOut_payload_0_10594);
  assign _zz_dataOut_payload_0_10663 = (_zz_dataOut_payload_0_10597 < _zz_dataOut_payload_0_10609);
  assign _zz_dataOut_payload_0_10664 = (_zz_dataOut_payload_0_10663 ? _zz_dataOut_payload_0_10597 : _zz_dataOut_payload_0_10609);
  assign _zz_dataOut_payload_0_10665 = (_zz_dataOut_payload_0_10663 ? _zz_dataOut_payload_0_10609 : _zz_dataOut_payload_0_10597);
  assign _zz_dataOut_payload_0_10666 = (_zz_dataOut_payload_0_10600 < _zz_dataOut_payload_0_10612);
  assign _zz_dataOut_payload_0_10667 = (_zz_dataOut_payload_0_10666 ? _zz_dataOut_payload_0_10600 : _zz_dataOut_payload_0_10612);
  assign _zz_dataOut_payload_0_10668 = (_zz_dataOut_payload_0_10666 ? _zz_dataOut_payload_0_10612 : _zz_dataOut_payload_0_10600);
  assign _zz_dataOut_payload_0_10669 = (_zz_dataOut_payload_0_10603 < _zz_dataOut_payload_0_10615);
  assign _zz_dataOut_payload_0_10670 = (_zz_dataOut_payload_0_10669 ? _zz_dataOut_payload_0_10603 : _zz_dataOut_payload_0_10615);
  assign _zz_dataOut_payload_0_10671 = (_zz_dataOut_payload_0_10669 ? _zz_dataOut_payload_0_10615 : _zz_dataOut_payload_0_10603);
  assign _zz_dataOut_payload_0_10672 = (_zz_dataOut_payload_0_10661 < _zz_dataOut_payload_0_10667);
  assign _zz_dataOut_payload_0_10673 = (_zz_dataOut_payload_0_10672 ? _zz_dataOut_payload_0_10661 : _zz_dataOut_payload_0_10667);
  assign _zz_dataOut_payload_0_10674 = (_zz_dataOut_payload_0_10672 ? _zz_dataOut_payload_0_10667 : _zz_dataOut_payload_0_10661);
  assign _zz_dataOut_payload_0_10675 = (_zz_dataOut_payload_0_10664 < _zz_dataOut_payload_0_10670);
  assign _zz_dataOut_payload_0_10676 = (_zz_dataOut_payload_0_10675 ? _zz_dataOut_payload_0_10664 : _zz_dataOut_payload_0_10670);
  assign _zz_dataOut_payload_0_10677 = (_zz_dataOut_payload_0_10675 ? _zz_dataOut_payload_0_10670 : _zz_dataOut_payload_0_10664);
  assign _zz_dataOut_payload_0_10678 = (_zz_dataOut_payload_0_10673 < _zz_dataOut_payload_0_10676);
  assign _zz_dataOut_payload_0_10679 = (_zz_dataOut_payload_0_10674 < _zz_dataOut_payload_0_10677);
  assign _zz_dataOut_payload_0_10684 = (_zz_dataOut_payload_0_10662 < _zz_dataOut_payload_0_10668);
  assign _zz_dataOut_payload_0_10685 = (_zz_dataOut_payload_0_10684 ? _zz_dataOut_payload_0_10662 : _zz_dataOut_payload_0_10668);
  assign _zz_dataOut_payload_0_10686 = (_zz_dataOut_payload_0_10684 ? _zz_dataOut_payload_0_10668 : _zz_dataOut_payload_0_10662);
  assign _zz_dataOut_payload_0_10687 = (_zz_dataOut_payload_0_10665 < _zz_dataOut_payload_0_10671);
  assign _zz_dataOut_payload_0_10688 = (_zz_dataOut_payload_0_10687 ? _zz_dataOut_payload_0_10665 : _zz_dataOut_payload_0_10671);
  assign _zz_dataOut_payload_0_10689 = (_zz_dataOut_payload_0_10687 ? _zz_dataOut_payload_0_10671 : _zz_dataOut_payload_0_10665);
  assign _zz_dataOut_payload_0_10690 = (_zz_dataOut_payload_0_10685 < _zz_dataOut_payload_0_10688);
  assign _zz_dataOut_payload_0_10691 = (_zz_dataOut_payload_0_10686 < _zz_dataOut_payload_0_10689);
  assign _zz_dataOut_payload_0_10816 = (_zz_dataOut_payload_0_8256 < _zz_dataOut_payload_0_8319);
  assign _zz_dataOut_payload_0_10817 = (_zz_dataOut_payload_0_10816 ? _zz_dataOut_payload_0_8256 : _zz_dataOut_payload_0_8319);
  assign _zz_dataOut_payload_0_10818 = (_zz_dataOut_payload_0_10816 ? _zz_dataOut_payload_0_8319 : _zz_dataOut_payload_0_8256);
  assign _zz_dataOut_payload_0_10819 = (_zz_dataOut_payload_0_8257 < _zz_dataOut_payload_0_8318);
  assign _zz_dataOut_payload_0_10820 = (_zz_dataOut_payload_0_10819 ? _zz_dataOut_payload_0_8257 : _zz_dataOut_payload_0_8318);
  assign _zz_dataOut_payload_0_10821 = (_zz_dataOut_payload_0_10819 ? _zz_dataOut_payload_0_8318 : _zz_dataOut_payload_0_8257);
  assign _zz_dataOut_payload_0_10822 = (_zz_dataOut_payload_0_8258 < _zz_dataOut_payload_0_8317);
  assign _zz_dataOut_payload_0_10823 = (_zz_dataOut_payload_0_10822 ? _zz_dataOut_payload_0_8258 : _zz_dataOut_payload_0_8317);
  assign _zz_dataOut_payload_0_10824 = (_zz_dataOut_payload_0_10822 ? _zz_dataOut_payload_0_8317 : _zz_dataOut_payload_0_8258);
  assign _zz_dataOut_payload_0_10825 = (_zz_dataOut_payload_0_8259 < _zz_dataOut_payload_0_8316);
  assign _zz_dataOut_payload_0_10826 = (_zz_dataOut_payload_0_10825 ? _zz_dataOut_payload_0_8259 : _zz_dataOut_payload_0_8316);
  assign _zz_dataOut_payload_0_10827 = (_zz_dataOut_payload_0_10825 ? _zz_dataOut_payload_0_8316 : _zz_dataOut_payload_0_8259);
  assign _zz_dataOut_payload_0_10828 = (_zz_dataOut_payload_0_8260 < _zz_dataOut_payload_0_8315);
  assign _zz_dataOut_payload_0_10829 = (_zz_dataOut_payload_0_10828 ? _zz_dataOut_payload_0_8260 : _zz_dataOut_payload_0_8315);
  assign _zz_dataOut_payload_0_10830 = (_zz_dataOut_payload_0_10828 ? _zz_dataOut_payload_0_8315 : _zz_dataOut_payload_0_8260);
  assign _zz_dataOut_payload_0_10831 = (_zz_dataOut_payload_0_8261 < _zz_dataOut_payload_0_8314);
  assign _zz_dataOut_payload_0_10832 = (_zz_dataOut_payload_0_10831 ? _zz_dataOut_payload_0_8261 : _zz_dataOut_payload_0_8314);
  assign _zz_dataOut_payload_0_10833 = (_zz_dataOut_payload_0_10831 ? _zz_dataOut_payload_0_8314 : _zz_dataOut_payload_0_8261);
  assign _zz_dataOut_payload_0_10834 = (_zz_dataOut_payload_0_8262 < _zz_dataOut_payload_0_8313);
  assign _zz_dataOut_payload_0_10835 = (_zz_dataOut_payload_0_10834 ? _zz_dataOut_payload_0_8262 : _zz_dataOut_payload_0_8313);
  assign _zz_dataOut_payload_0_10836 = (_zz_dataOut_payload_0_10834 ? _zz_dataOut_payload_0_8313 : _zz_dataOut_payload_0_8262);
  assign _zz_dataOut_payload_0_10837 = (_zz_dataOut_payload_0_8263 < _zz_dataOut_payload_0_8312);
  assign _zz_dataOut_payload_0_10838 = (_zz_dataOut_payload_0_10837 ? _zz_dataOut_payload_0_8263 : _zz_dataOut_payload_0_8312);
  assign _zz_dataOut_payload_0_10839 = (_zz_dataOut_payload_0_10837 ? _zz_dataOut_payload_0_8312 : _zz_dataOut_payload_0_8263);
  assign _zz_dataOut_payload_0_10840 = (_zz_dataOut_payload_0_8264 < _zz_dataOut_payload_0_8311);
  assign _zz_dataOut_payload_0_10841 = (_zz_dataOut_payload_0_10840 ? _zz_dataOut_payload_0_8264 : _zz_dataOut_payload_0_8311);
  assign _zz_dataOut_payload_0_10842 = (_zz_dataOut_payload_0_10840 ? _zz_dataOut_payload_0_8311 : _zz_dataOut_payload_0_8264);
  assign _zz_dataOut_payload_0_10843 = (_zz_dataOut_payload_0_8265 < _zz_dataOut_payload_0_8310);
  assign _zz_dataOut_payload_0_10844 = (_zz_dataOut_payload_0_10843 ? _zz_dataOut_payload_0_8265 : _zz_dataOut_payload_0_8310);
  assign _zz_dataOut_payload_0_10845 = (_zz_dataOut_payload_0_10843 ? _zz_dataOut_payload_0_8310 : _zz_dataOut_payload_0_8265);
  assign _zz_dataOut_payload_0_10846 = (_zz_dataOut_payload_0_8266 < _zz_dataOut_payload_0_8309);
  assign _zz_dataOut_payload_0_10847 = (_zz_dataOut_payload_0_10846 ? _zz_dataOut_payload_0_8266 : _zz_dataOut_payload_0_8309);
  assign _zz_dataOut_payload_0_10848 = (_zz_dataOut_payload_0_10846 ? _zz_dataOut_payload_0_8309 : _zz_dataOut_payload_0_8266);
  assign _zz_dataOut_payload_0_10849 = (_zz_dataOut_payload_0_8267 < _zz_dataOut_payload_0_8308);
  assign _zz_dataOut_payload_0_10850 = (_zz_dataOut_payload_0_10849 ? _zz_dataOut_payload_0_8267 : _zz_dataOut_payload_0_8308);
  assign _zz_dataOut_payload_0_10851 = (_zz_dataOut_payload_0_10849 ? _zz_dataOut_payload_0_8308 : _zz_dataOut_payload_0_8267);
  assign _zz_dataOut_payload_0_10852 = (_zz_dataOut_payload_0_8268 < _zz_dataOut_payload_0_8307);
  assign _zz_dataOut_payload_0_10853 = (_zz_dataOut_payload_0_10852 ? _zz_dataOut_payload_0_8268 : _zz_dataOut_payload_0_8307);
  assign _zz_dataOut_payload_0_10854 = (_zz_dataOut_payload_0_10852 ? _zz_dataOut_payload_0_8307 : _zz_dataOut_payload_0_8268);
  assign _zz_dataOut_payload_0_10855 = (_zz_dataOut_payload_0_8269 < _zz_dataOut_payload_0_8306);
  assign _zz_dataOut_payload_0_10856 = (_zz_dataOut_payload_0_10855 ? _zz_dataOut_payload_0_8269 : _zz_dataOut_payload_0_8306);
  assign _zz_dataOut_payload_0_10857 = (_zz_dataOut_payload_0_10855 ? _zz_dataOut_payload_0_8306 : _zz_dataOut_payload_0_8269);
  assign _zz_dataOut_payload_0_10858 = (_zz_dataOut_payload_0_8270 < _zz_dataOut_payload_0_8305);
  assign _zz_dataOut_payload_0_10859 = (_zz_dataOut_payload_0_10858 ? _zz_dataOut_payload_0_8270 : _zz_dataOut_payload_0_8305);
  assign _zz_dataOut_payload_0_10860 = (_zz_dataOut_payload_0_10858 ? _zz_dataOut_payload_0_8305 : _zz_dataOut_payload_0_8270);
  assign _zz_dataOut_payload_0_10861 = (_zz_dataOut_payload_0_8271 < _zz_dataOut_payload_0_8304);
  assign _zz_dataOut_payload_0_10862 = (_zz_dataOut_payload_0_10861 ? _zz_dataOut_payload_0_8271 : _zz_dataOut_payload_0_8304);
  assign _zz_dataOut_payload_0_10863 = (_zz_dataOut_payload_0_10861 ? _zz_dataOut_payload_0_8304 : _zz_dataOut_payload_0_8271);
  assign _zz_dataOut_payload_0_10864 = (_zz_dataOut_payload_0_8272 < _zz_dataOut_payload_0_8303);
  assign _zz_dataOut_payload_0_10865 = (_zz_dataOut_payload_0_10864 ? _zz_dataOut_payload_0_8272 : _zz_dataOut_payload_0_8303);
  assign _zz_dataOut_payload_0_10866 = (_zz_dataOut_payload_0_10864 ? _zz_dataOut_payload_0_8303 : _zz_dataOut_payload_0_8272);
  assign _zz_dataOut_payload_0_10867 = (_zz_dataOut_payload_0_8273 < _zz_dataOut_payload_0_8302);
  assign _zz_dataOut_payload_0_10868 = (_zz_dataOut_payload_0_10867 ? _zz_dataOut_payload_0_8273 : _zz_dataOut_payload_0_8302);
  assign _zz_dataOut_payload_0_10869 = (_zz_dataOut_payload_0_10867 ? _zz_dataOut_payload_0_8302 : _zz_dataOut_payload_0_8273);
  assign _zz_dataOut_payload_0_10870 = (_zz_dataOut_payload_0_8274 < _zz_dataOut_payload_0_8301);
  assign _zz_dataOut_payload_0_10871 = (_zz_dataOut_payload_0_10870 ? _zz_dataOut_payload_0_8274 : _zz_dataOut_payload_0_8301);
  assign _zz_dataOut_payload_0_10872 = (_zz_dataOut_payload_0_10870 ? _zz_dataOut_payload_0_8301 : _zz_dataOut_payload_0_8274);
  assign _zz_dataOut_payload_0_10873 = (_zz_dataOut_payload_0_8275 < _zz_dataOut_payload_0_8300);
  assign _zz_dataOut_payload_0_10874 = (_zz_dataOut_payload_0_10873 ? _zz_dataOut_payload_0_8275 : _zz_dataOut_payload_0_8300);
  assign _zz_dataOut_payload_0_10875 = (_zz_dataOut_payload_0_10873 ? _zz_dataOut_payload_0_8300 : _zz_dataOut_payload_0_8275);
  assign _zz_dataOut_payload_0_10876 = (_zz_dataOut_payload_0_8276 < _zz_dataOut_payload_0_8299);
  assign _zz_dataOut_payload_0_10877 = (_zz_dataOut_payload_0_10876 ? _zz_dataOut_payload_0_8276 : _zz_dataOut_payload_0_8299);
  assign _zz_dataOut_payload_0_10878 = (_zz_dataOut_payload_0_10876 ? _zz_dataOut_payload_0_8299 : _zz_dataOut_payload_0_8276);
  assign _zz_dataOut_payload_0_10879 = (_zz_dataOut_payload_0_8277 < _zz_dataOut_payload_0_8298);
  assign _zz_dataOut_payload_0_10880 = (_zz_dataOut_payload_0_10879 ? _zz_dataOut_payload_0_8277 : _zz_dataOut_payload_0_8298);
  assign _zz_dataOut_payload_0_10881 = (_zz_dataOut_payload_0_10879 ? _zz_dataOut_payload_0_8298 : _zz_dataOut_payload_0_8277);
  assign _zz_dataOut_payload_0_10882 = (_zz_dataOut_payload_0_8278 < _zz_dataOut_payload_0_8297);
  assign _zz_dataOut_payload_0_10883 = (_zz_dataOut_payload_0_10882 ? _zz_dataOut_payload_0_8278 : _zz_dataOut_payload_0_8297);
  assign _zz_dataOut_payload_0_10884 = (_zz_dataOut_payload_0_10882 ? _zz_dataOut_payload_0_8297 : _zz_dataOut_payload_0_8278);
  assign _zz_dataOut_payload_0_10885 = (_zz_dataOut_payload_0_8279 < _zz_dataOut_payload_0_8296);
  assign _zz_dataOut_payload_0_10886 = (_zz_dataOut_payload_0_10885 ? _zz_dataOut_payload_0_8279 : _zz_dataOut_payload_0_8296);
  assign _zz_dataOut_payload_0_10887 = (_zz_dataOut_payload_0_10885 ? _zz_dataOut_payload_0_8296 : _zz_dataOut_payload_0_8279);
  assign _zz_dataOut_payload_0_10888 = (_zz_dataOut_payload_0_8280 < _zz_dataOut_payload_0_8295);
  assign _zz_dataOut_payload_0_10889 = (_zz_dataOut_payload_0_10888 ? _zz_dataOut_payload_0_8280 : _zz_dataOut_payload_0_8295);
  assign _zz_dataOut_payload_0_10890 = (_zz_dataOut_payload_0_10888 ? _zz_dataOut_payload_0_8295 : _zz_dataOut_payload_0_8280);
  assign _zz_dataOut_payload_0_10891 = (_zz_dataOut_payload_0_8281 < _zz_dataOut_payload_0_8294);
  assign _zz_dataOut_payload_0_10892 = (_zz_dataOut_payload_0_10891 ? _zz_dataOut_payload_0_8281 : _zz_dataOut_payload_0_8294);
  assign _zz_dataOut_payload_0_10893 = (_zz_dataOut_payload_0_10891 ? _zz_dataOut_payload_0_8294 : _zz_dataOut_payload_0_8281);
  assign _zz_dataOut_payload_0_10894 = (_zz_dataOut_payload_0_8282 < _zz_dataOut_payload_0_8293);
  assign _zz_dataOut_payload_0_10895 = (_zz_dataOut_payload_0_10894 ? _zz_dataOut_payload_0_8282 : _zz_dataOut_payload_0_8293);
  assign _zz_dataOut_payload_0_10896 = (_zz_dataOut_payload_0_10894 ? _zz_dataOut_payload_0_8293 : _zz_dataOut_payload_0_8282);
  assign _zz_dataOut_payload_0_10897 = (_zz_dataOut_payload_0_8283 < _zz_dataOut_payload_0_8292);
  assign _zz_dataOut_payload_0_10898 = (_zz_dataOut_payload_0_10897 ? _zz_dataOut_payload_0_8283 : _zz_dataOut_payload_0_8292);
  assign _zz_dataOut_payload_0_10899 = (_zz_dataOut_payload_0_10897 ? _zz_dataOut_payload_0_8292 : _zz_dataOut_payload_0_8283);
  assign _zz_dataOut_payload_0_10900 = (_zz_dataOut_payload_0_8284 < _zz_dataOut_payload_0_8291);
  assign _zz_dataOut_payload_0_10901 = (_zz_dataOut_payload_0_10900 ? _zz_dataOut_payload_0_8284 : _zz_dataOut_payload_0_8291);
  assign _zz_dataOut_payload_0_10902 = (_zz_dataOut_payload_0_10900 ? _zz_dataOut_payload_0_8291 : _zz_dataOut_payload_0_8284);
  assign _zz_dataOut_payload_0_10903 = (_zz_dataOut_payload_0_8285 < _zz_dataOut_payload_0_8290);
  assign _zz_dataOut_payload_0_10904 = (_zz_dataOut_payload_0_10903 ? _zz_dataOut_payload_0_8285 : _zz_dataOut_payload_0_8290);
  assign _zz_dataOut_payload_0_10905 = (_zz_dataOut_payload_0_10903 ? _zz_dataOut_payload_0_8290 : _zz_dataOut_payload_0_8285);
  assign _zz_dataOut_payload_0_10906 = (_zz_dataOut_payload_0_8286 < _zz_dataOut_payload_0_8289);
  assign _zz_dataOut_payload_0_10907 = (_zz_dataOut_payload_0_10906 ? _zz_dataOut_payload_0_8286 : _zz_dataOut_payload_0_8289);
  assign _zz_dataOut_payload_0_10908 = (_zz_dataOut_payload_0_10906 ? _zz_dataOut_payload_0_8289 : _zz_dataOut_payload_0_8286);
  assign _zz_dataOut_payload_0_10909 = (_zz_dataOut_payload_0_8287 < _zz_dataOut_payload_0_8288);
  assign _zz_dataOut_payload_0_10910 = (_zz_dataOut_payload_0_10909 ? _zz_dataOut_payload_0_8287 : _zz_dataOut_payload_0_8288);
  assign _zz_dataOut_payload_0_10911 = (_zz_dataOut_payload_0_10909 ? _zz_dataOut_payload_0_8288 : _zz_dataOut_payload_0_8287);
  assign _zz_dataOut_payload_0_10912 = (_zz_dataOut_payload_0_10817 < _zz_dataOut_payload_0_10865);
  assign _zz_dataOut_payload_0_10913 = (_zz_dataOut_payload_0_10912 ? _zz_dataOut_payload_0_10817 : _zz_dataOut_payload_0_10865);
  assign _zz_dataOut_payload_0_10914 = (_zz_dataOut_payload_0_10912 ? _zz_dataOut_payload_0_10865 : _zz_dataOut_payload_0_10817);
  assign _zz_dataOut_payload_0_10915 = (_zz_dataOut_payload_0_10820 < _zz_dataOut_payload_0_10868);
  assign _zz_dataOut_payload_0_10916 = (_zz_dataOut_payload_0_10915 ? _zz_dataOut_payload_0_10820 : _zz_dataOut_payload_0_10868);
  assign _zz_dataOut_payload_0_10917 = (_zz_dataOut_payload_0_10915 ? _zz_dataOut_payload_0_10868 : _zz_dataOut_payload_0_10820);
  assign _zz_dataOut_payload_0_10918 = (_zz_dataOut_payload_0_10823 < _zz_dataOut_payload_0_10871);
  assign _zz_dataOut_payload_0_10919 = (_zz_dataOut_payload_0_10918 ? _zz_dataOut_payload_0_10823 : _zz_dataOut_payload_0_10871);
  assign _zz_dataOut_payload_0_10920 = (_zz_dataOut_payload_0_10918 ? _zz_dataOut_payload_0_10871 : _zz_dataOut_payload_0_10823);
  assign _zz_dataOut_payload_0_10921 = (_zz_dataOut_payload_0_10826 < _zz_dataOut_payload_0_10874);
  assign _zz_dataOut_payload_0_10922 = (_zz_dataOut_payload_0_10921 ? _zz_dataOut_payload_0_10826 : _zz_dataOut_payload_0_10874);
  assign _zz_dataOut_payload_0_10923 = (_zz_dataOut_payload_0_10921 ? _zz_dataOut_payload_0_10874 : _zz_dataOut_payload_0_10826);
  assign _zz_dataOut_payload_0_10924 = (_zz_dataOut_payload_0_10829 < _zz_dataOut_payload_0_10877);
  assign _zz_dataOut_payload_0_10925 = (_zz_dataOut_payload_0_10924 ? _zz_dataOut_payload_0_10829 : _zz_dataOut_payload_0_10877);
  assign _zz_dataOut_payload_0_10926 = (_zz_dataOut_payload_0_10924 ? _zz_dataOut_payload_0_10877 : _zz_dataOut_payload_0_10829);
  assign _zz_dataOut_payload_0_10927 = (_zz_dataOut_payload_0_10832 < _zz_dataOut_payload_0_10880);
  assign _zz_dataOut_payload_0_10928 = (_zz_dataOut_payload_0_10927 ? _zz_dataOut_payload_0_10832 : _zz_dataOut_payload_0_10880);
  assign _zz_dataOut_payload_0_10929 = (_zz_dataOut_payload_0_10927 ? _zz_dataOut_payload_0_10880 : _zz_dataOut_payload_0_10832);
  assign _zz_dataOut_payload_0_10930 = (_zz_dataOut_payload_0_10835 < _zz_dataOut_payload_0_10883);
  assign _zz_dataOut_payload_0_10931 = (_zz_dataOut_payload_0_10930 ? _zz_dataOut_payload_0_10835 : _zz_dataOut_payload_0_10883);
  assign _zz_dataOut_payload_0_10932 = (_zz_dataOut_payload_0_10930 ? _zz_dataOut_payload_0_10883 : _zz_dataOut_payload_0_10835);
  assign _zz_dataOut_payload_0_10933 = (_zz_dataOut_payload_0_10838 < _zz_dataOut_payload_0_10886);
  assign _zz_dataOut_payload_0_10934 = (_zz_dataOut_payload_0_10933 ? _zz_dataOut_payload_0_10838 : _zz_dataOut_payload_0_10886);
  assign _zz_dataOut_payload_0_10935 = (_zz_dataOut_payload_0_10933 ? _zz_dataOut_payload_0_10886 : _zz_dataOut_payload_0_10838);
  assign _zz_dataOut_payload_0_10936 = (_zz_dataOut_payload_0_10841 < _zz_dataOut_payload_0_10889);
  assign _zz_dataOut_payload_0_10937 = (_zz_dataOut_payload_0_10936 ? _zz_dataOut_payload_0_10841 : _zz_dataOut_payload_0_10889);
  assign _zz_dataOut_payload_0_10938 = (_zz_dataOut_payload_0_10936 ? _zz_dataOut_payload_0_10889 : _zz_dataOut_payload_0_10841);
  assign _zz_dataOut_payload_0_10939 = (_zz_dataOut_payload_0_10844 < _zz_dataOut_payload_0_10892);
  assign _zz_dataOut_payload_0_10940 = (_zz_dataOut_payload_0_10939 ? _zz_dataOut_payload_0_10844 : _zz_dataOut_payload_0_10892);
  assign _zz_dataOut_payload_0_10941 = (_zz_dataOut_payload_0_10939 ? _zz_dataOut_payload_0_10892 : _zz_dataOut_payload_0_10844);
  assign _zz_dataOut_payload_0_10942 = (_zz_dataOut_payload_0_10847 < _zz_dataOut_payload_0_10895);
  assign _zz_dataOut_payload_0_10943 = (_zz_dataOut_payload_0_10942 ? _zz_dataOut_payload_0_10847 : _zz_dataOut_payload_0_10895);
  assign _zz_dataOut_payload_0_10944 = (_zz_dataOut_payload_0_10942 ? _zz_dataOut_payload_0_10895 : _zz_dataOut_payload_0_10847);
  assign _zz_dataOut_payload_0_10945 = (_zz_dataOut_payload_0_10850 < _zz_dataOut_payload_0_10898);
  assign _zz_dataOut_payload_0_10946 = (_zz_dataOut_payload_0_10945 ? _zz_dataOut_payload_0_10850 : _zz_dataOut_payload_0_10898);
  assign _zz_dataOut_payload_0_10947 = (_zz_dataOut_payload_0_10945 ? _zz_dataOut_payload_0_10898 : _zz_dataOut_payload_0_10850);
  assign _zz_dataOut_payload_0_10948 = (_zz_dataOut_payload_0_10853 < _zz_dataOut_payload_0_10901);
  assign _zz_dataOut_payload_0_10949 = (_zz_dataOut_payload_0_10948 ? _zz_dataOut_payload_0_10853 : _zz_dataOut_payload_0_10901);
  assign _zz_dataOut_payload_0_10950 = (_zz_dataOut_payload_0_10948 ? _zz_dataOut_payload_0_10901 : _zz_dataOut_payload_0_10853);
  assign _zz_dataOut_payload_0_10951 = (_zz_dataOut_payload_0_10856 < _zz_dataOut_payload_0_10904);
  assign _zz_dataOut_payload_0_10952 = (_zz_dataOut_payload_0_10951 ? _zz_dataOut_payload_0_10856 : _zz_dataOut_payload_0_10904);
  assign _zz_dataOut_payload_0_10953 = (_zz_dataOut_payload_0_10951 ? _zz_dataOut_payload_0_10904 : _zz_dataOut_payload_0_10856);
  assign _zz_dataOut_payload_0_10954 = (_zz_dataOut_payload_0_10859 < _zz_dataOut_payload_0_10907);
  assign _zz_dataOut_payload_0_10955 = (_zz_dataOut_payload_0_10954 ? _zz_dataOut_payload_0_10859 : _zz_dataOut_payload_0_10907);
  assign _zz_dataOut_payload_0_10956 = (_zz_dataOut_payload_0_10954 ? _zz_dataOut_payload_0_10907 : _zz_dataOut_payload_0_10859);
  assign _zz_dataOut_payload_0_10957 = (_zz_dataOut_payload_0_10862 < _zz_dataOut_payload_0_10910);
  assign _zz_dataOut_payload_0_10958 = (_zz_dataOut_payload_0_10957 ? _zz_dataOut_payload_0_10862 : _zz_dataOut_payload_0_10910);
  assign _zz_dataOut_payload_0_10959 = (_zz_dataOut_payload_0_10957 ? _zz_dataOut_payload_0_10910 : _zz_dataOut_payload_0_10862);
  assign _zz_dataOut_payload_0_10960 = (_zz_dataOut_payload_0_10913 < _zz_dataOut_payload_0_10937);
  assign _zz_dataOut_payload_0_10961 = (_zz_dataOut_payload_0_10960 ? _zz_dataOut_payload_0_10913 : _zz_dataOut_payload_0_10937);
  assign _zz_dataOut_payload_0_10962 = (_zz_dataOut_payload_0_10960 ? _zz_dataOut_payload_0_10937 : _zz_dataOut_payload_0_10913);
  assign _zz_dataOut_payload_0_10963 = (_zz_dataOut_payload_0_10916 < _zz_dataOut_payload_0_10940);
  assign _zz_dataOut_payload_0_10964 = (_zz_dataOut_payload_0_10963 ? _zz_dataOut_payload_0_10916 : _zz_dataOut_payload_0_10940);
  assign _zz_dataOut_payload_0_10965 = (_zz_dataOut_payload_0_10963 ? _zz_dataOut_payload_0_10940 : _zz_dataOut_payload_0_10916);
  assign _zz_dataOut_payload_0_10966 = (_zz_dataOut_payload_0_10919 < _zz_dataOut_payload_0_10943);
  assign _zz_dataOut_payload_0_10967 = (_zz_dataOut_payload_0_10966 ? _zz_dataOut_payload_0_10919 : _zz_dataOut_payload_0_10943);
  assign _zz_dataOut_payload_0_10968 = (_zz_dataOut_payload_0_10966 ? _zz_dataOut_payload_0_10943 : _zz_dataOut_payload_0_10919);
  assign _zz_dataOut_payload_0_10969 = (_zz_dataOut_payload_0_10922 < _zz_dataOut_payload_0_10946);
  assign _zz_dataOut_payload_0_10970 = (_zz_dataOut_payload_0_10969 ? _zz_dataOut_payload_0_10922 : _zz_dataOut_payload_0_10946);
  assign _zz_dataOut_payload_0_10971 = (_zz_dataOut_payload_0_10969 ? _zz_dataOut_payload_0_10946 : _zz_dataOut_payload_0_10922);
  assign _zz_dataOut_payload_0_10972 = (_zz_dataOut_payload_0_10925 < _zz_dataOut_payload_0_10949);
  assign _zz_dataOut_payload_0_10973 = (_zz_dataOut_payload_0_10972 ? _zz_dataOut_payload_0_10925 : _zz_dataOut_payload_0_10949);
  assign _zz_dataOut_payload_0_10974 = (_zz_dataOut_payload_0_10972 ? _zz_dataOut_payload_0_10949 : _zz_dataOut_payload_0_10925);
  assign _zz_dataOut_payload_0_10975 = (_zz_dataOut_payload_0_10928 < _zz_dataOut_payload_0_10952);
  assign _zz_dataOut_payload_0_10976 = (_zz_dataOut_payload_0_10975 ? _zz_dataOut_payload_0_10928 : _zz_dataOut_payload_0_10952);
  assign _zz_dataOut_payload_0_10977 = (_zz_dataOut_payload_0_10975 ? _zz_dataOut_payload_0_10952 : _zz_dataOut_payload_0_10928);
  assign _zz_dataOut_payload_0_10978 = (_zz_dataOut_payload_0_10931 < _zz_dataOut_payload_0_10955);
  assign _zz_dataOut_payload_0_10979 = (_zz_dataOut_payload_0_10978 ? _zz_dataOut_payload_0_10931 : _zz_dataOut_payload_0_10955);
  assign _zz_dataOut_payload_0_10980 = (_zz_dataOut_payload_0_10978 ? _zz_dataOut_payload_0_10955 : _zz_dataOut_payload_0_10931);
  assign _zz_dataOut_payload_0_10981 = (_zz_dataOut_payload_0_10934 < _zz_dataOut_payload_0_10958);
  assign _zz_dataOut_payload_0_10982 = (_zz_dataOut_payload_0_10981 ? _zz_dataOut_payload_0_10934 : _zz_dataOut_payload_0_10958);
  assign _zz_dataOut_payload_0_10983 = (_zz_dataOut_payload_0_10981 ? _zz_dataOut_payload_0_10958 : _zz_dataOut_payload_0_10934);
  assign _zz_dataOut_payload_0_10984 = (_zz_dataOut_payload_0_10961 < _zz_dataOut_payload_0_10973);
  assign _zz_dataOut_payload_0_10985 = (_zz_dataOut_payload_0_10984 ? _zz_dataOut_payload_0_10961 : _zz_dataOut_payload_0_10973);
  assign _zz_dataOut_payload_0_10986 = (_zz_dataOut_payload_0_10984 ? _zz_dataOut_payload_0_10973 : _zz_dataOut_payload_0_10961);
  assign _zz_dataOut_payload_0_10987 = (_zz_dataOut_payload_0_10964 < _zz_dataOut_payload_0_10976);
  assign _zz_dataOut_payload_0_10988 = (_zz_dataOut_payload_0_10987 ? _zz_dataOut_payload_0_10964 : _zz_dataOut_payload_0_10976);
  assign _zz_dataOut_payload_0_10989 = (_zz_dataOut_payload_0_10987 ? _zz_dataOut_payload_0_10976 : _zz_dataOut_payload_0_10964);
  assign _zz_dataOut_payload_0_10990 = (_zz_dataOut_payload_0_10967 < _zz_dataOut_payload_0_10979);
  assign _zz_dataOut_payload_0_10991 = (_zz_dataOut_payload_0_10990 ? _zz_dataOut_payload_0_10967 : _zz_dataOut_payload_0_10979);
  assign _zz_dataOut_payload_0_10992 = (_zz_dataOut_payload_0_10990 ? _zz_dataOut_payload_0_10979 : _zz_dataOut_payload_0_10967);
  assign _zz_dataOut_payload_0_10993 = (_zz_dataOut_payload_0_10970 < _zz_dataOut_payload_0_10982);
  assign _zz_dataOut_payload_0_10994 = (_zz_dataOut_payload_0_10993 ? _zz_dataOut_payload_0_10970 : _zz_dataOut_payload_0_10982);
  assign _zz_dataOut_payload_0_10995 = (_zz_dataOut_payload_0_10993 ? _zz_dataOut_payload_0_10982 : _zz_dataOut_payload_0_10970);
  assign _zz_dataOut_payload_0_10996 = (_zz_dataOut_payload_0_10985 < _zz_dataOut_payload_0_10991);
  assign _zz_dataOut_payload_0_10997 = (_zz_dataOut_payload_0_10996 ? _zz_dataOut_payload_0_10985 : _zz_dataOut_payload_0_10991);
  assign _zz_dataOut_payload_0_10998 = (_zz_dataOut_payload_0_10996 ? _zz_dataOut_payload_0_10991 : _zz_dataOut_payload_0_10985);
  assign _zz_dataOut_payload_0_10999 = (_zz_dataOut_payload_0_10988 < _zz_dataOut_payload_0_10994);
  assign _zz_dataOut_payload_0_11000 = (_zz_dataOut_payload_0_10999 ? _zz_dataOut_payload_0_10988 : _zz_dataOut_payload_0_10994);
  assign _zz_dataOut_payload_0_11001 = (_zz_dataOut_payload_0_10999 ? _zz_dataOut_payload_0_10994 : _zz_dataOut_payload_0_10988);
  assign _zz_dataOut_payload_0_11002 = (_zz_dataOut_payload_0_10997 < _zz_dataOut_payload_0_11000);
  assign _zz_dataOut_payload_0_11003 = (_zz_dataOut_payload_0_10998 < _zz_dataOut_payload_0_11001);
  assign _zz_dataOut_payload_0_11008 = (_zz_dataOut_payload_0_10986 < _zz_dataOut_payload_0_10992);
  assign _zz_dataOut_payload_0_11009 = (_zz_dataOut_payload_0_11008 ? _zz_dataOut_payload_0_10986 : _zz_dataOut_payload_0_10992);
  assign _zz_dataOut_payload_0_11010 = (_zz_dataOut_payload_0_11008 ? _zz_dataOut_payload_0_10992 : _zz_dataOut_payload_0_10986);
  assign _zz_dataOut_payload_0_11011 = (_zz_dataOut_payload_0_10989 < _zz_dataOut_payload_0_10995);
  assign _zz_dataOut_payload_0_11012 = (_zz_dataOut_payload_0_11011 ? _zz_dataOut_payload_0_10989 : _zz_dataOut_payload_0_10995);
  assign _zz_dataOut_payload_0_11013 = (_zz_dataOut_payload_0_11011 ? _zz_dataOut_payload_0_10995 : _zz_dataOut_payload_0_10989);
  assign _zz_dataOut_payload_0_11014 = (_zz_dataOut_payload_0_11009 < _zz_dataOut_payload_0_11012);
  assign _zz_dataOut_payload_0_11015 = (_zz_dataOut_payload_0_11010 < _zz_dataOut_payload_0_11013);
  assign _zz_dataOut_payload_0_11028 = (_zz_dataOut_payload_0_10962 < _zz_dataOut_payload_0_10974);
  assign _zz_dataOut_payload_0_11029 = (_zz_dataOut_payload_0_11028 ? _zz_dataOut_payload_0_10962 : _zz_dataOut_payload_0_10974);
  assign _zz_dataOut_payload_0_11030 = (_zz_dataOut_payload_0_11028 ? _zz_dataOut_payload_0_10974 : _zz_dataOut_payload_0_10962);
  assign _zz_dataOut_payload_0_11031 = (_zz_dataOut_payload_0_10965 < _zz_dataOut_payload_0_10977);
  assign _zz_dataOut_payload_0_11032 = (_zz_dataOut_payload_0_11031 ? _zz_dataOut_payload_0_10965 : _zz_dataOut_payload_0_10977);
  assign _zz_dataOut_payload_0_11033 = (_zz_dataOut_payload_0_11031 ? _zz_dataOut_payload_0_10977 : _zz_dataOut_payload_0_10965);
  assign _zz_dataOut_payload_0_11034 = (_zz_dataOut_payload_0_10968 < _zz_dataOut_payload_0_10980);
  assign _zz_dataOut_payload_0_11035 = (_zz_dataOut_payload_0_11034 ? _zz_dataOut_payload_0_10968 : _zz_dataOut_payload_0_10980);
  assign _zz_dataOut_payload_0_11036 = (_zz_dataOut_payload_0_11034 ? _zz_dataOut_payload_0_10980 : _zz_dataOut_payload_0_10968);
  assign _zz_dataOut_payload_0_11037 = (_zz_dataOut_payload_0_10971 < _zz_dataOut_payload_0_10983);
  assign _zz_dataOut_payload_0_11038 = (_zz_dataOut_payload_0_11037 ? _zz_dataOut_payload_0_10971 : _zz_dataOut_payload_0_10983);
  assign _zz_dataOut_payload_0_11039 = (_zz_dataOut_payload_0_11037 ? _zz_dataOut_payload_0_10983 : _zz_dataOut_payload_0_10971);
  assign _zz_dataOut_payload_0_11040 = (_zz_dataOut_payload_0_11029 < _zz_dataOut_payload_0_11035);
  assign _zz_dataOut_payload_0_11041 = (_zz_dataOut_payload_0_11040 ? _zz_dataOut_payload_0_11029 : _zz_dataOut_payload_0_11035);
  assign _zz_dataOut_payload_0_11042 = (_zz_dataOut_payload_0_11040 ? _zz_dataOut_payload_0_11035 : _zz_dataOut_payload_0_11029);
  assign _zz_dataOut_payload_0_11043 = (_zz_dataOut_payload_0_11032 < _zz_dataOut_payload_0_11038);
  assign _zz_dataOut_payload_0_11044 = (_zz_dataOut_payload_0_11043 ? _zz_dataOut_payload_0_11032 : _zz_dataOut_payload_0_11038);
  assign _zz_dataOut_payload_0_11045 = (_zz_dataOut_payload_0_11043 ? _zz_dataOut_payload_0_11038 : _zz_dataOut_payload_0_11032);
  assign _zz_dataOut_payload_0_11046 = (_zz_dataOut_payload_0_11041 < _zz_dataOut_payload_0_11044);
  assign _zz_dataOut_payload_0_11047 = (_zz_dataOut_payload_0_11042 < _zz_dataOut_payload_0_11045);
  assign _zz_dataOut_payload_0_11052 = (_zz_dataOut_payload_0_11030 < _zz_dataOut_payload_0_11036);
  assign _zz_dataOut_payload_0_11053 = (_zz_dataOut_payload_0_11052 ? _zz_dataOut_payload_0_11030 : _zz_dataOut_payload_0_11036);
  assign _zz_dataOut_payload_0_11054 = (_zz_dataOut_payload_0_11052 ? _zz_dataOut_payload_0_11036 : _zz_dataOut_payload_0_11030);
  assign _zz_dataOut_payload_0_11055 = (_zz_dataOut_payload_0_11033 < _zz_dataOut_payload_0_11039);
  assign _zz_dataOut_payload_0_11056 = (_zz_dataOut_payload_0_11055 ? _zz_dataOut_payload_0_11033 : _zz_dataOut_payload_0_11039);
  assign _zz_dataOut_payload_0_11057 = (_zz_dataOut_payload_0_11055 ? _zz_dataOut_payload_0_11039 : _zz_dataOut_payload_0_11033);
  assign _zz_dataOut_payload_0_11058 = (_zz_dataOut_payload_0_11053 < _zz_dataOut_payload_0_11056);
  assign _zz_dataOut_payload_0_11059 = (_zz_dataOut_payload_0_11054 < _zz_dataOut_payload_0_11057);
  assign _zz_dataOut_payload_0_11088 = (_zz_dataOut_payload_0_10914 < _zz_dataOut_payload_0_10938);
  assign _zz_dataOut_payload_0_11089 = (_zz_dataOut_payload_0_11088 ? _zz_dataOut_payload_0_10914 : _zz_dataOut_payload_0_10938);
  assign _zz_dataOut_payload_0_11090 = (_zz_dataOut_payload_0_11088 ? _zz_dataOut_payload_0_10938 : _zz_dataOut_payload_0_10914);
  assign _zz_dataOut_payload_0_11091 = (_zz_dataOut_payload_0_10917 < _zz_dataOut_payload_0_10941);
  assign _zz_dataOut_payload_0_11092 = (_zz_dataOut_payload_0_11091 ? _zz_dataOut_payload_0_10917 : _zz_dataOut_payload_0_10941);
  assign _zz_dataOut_payload_0_11093 = (_zz_dataOut_payload_0_11091 ? _zz_dataOut_payload_0_10941 : _zz_dataOut_payload_0_10917);
  assign _zz_dataOut_payload_0_11094 = (_zz_dataOut_payload_0_10920 < _zz_dataOut_payload_0_10944);
  assign _zz_dataOut_payload_0_11095 = (_zz_dataOut_payload_0_11094 ? _zz_dataOut_payload_0_10920 : _zz_dataOut_payload_0_10944);
  assign _zz_dataOut_payload_0_11096 = (_zz_dataOut_payload_0_11094 ? _zz_dataOut_payload_0_10944 : _zz_dataOut_payload_0_10920);
  assign _zz_dataOut_payload_0_11097 = (_zz_dataOut_payload_0_10923 < _zz_dataOut_payload_0_10947);
  assign _zz_dataOut_payload_0_11098 = (_zz_dataOut_payload_0_11097 ? _zz_dataOut_payload_0_10923 : _zz_dataOut_payload_0_10947);
  assign _zz_dataOut_payload_0_11099 = (_zz_dataOut_payload_0_11097 ? _zz_dataOut_payload_0_10947 : _zz_dataOut_payload_0_10923);
  assign _zz_dataOut_payload_0_11100 = (_zz_dataOut_payload_0_10926 < _zz_dataOut_payload_0_10950);
  assign _zz_dataOut_payload_0_11101 = (_zz_dataOut_payload_0_11100 ? _zz_dataOut_payload_0_10926 : _zz_dataOut_payload_0_10950);
  assign _zz_dataOut_payload_0_11102 = (_zz_dataOut_payload_0_11100 ? _zz_dataOut_payload_0_10950 : _zz_dataOut_payload_0_10926);
  assign _zz_dataOut_payload_0_11103 = (_zz_dataOut_payload_0_10929 < _zz_dataOut_payload_0_10953);
  assign _zz_dataOut_payload_0_11104 = (_zz_dataOut_payload_0_11103 ? _zz_dataOut_payload_0_10929 : _zz_dataOut_payload_0_10953);
  assign _zz_dataOut_payload_0_11105 = (_zz_dataOut_payload_0_11103 ? _zz_dataOut_payload_0_10953 : _zz_dataOut_payload_0_10929);
  assign _zz_dataOut_payload_0_11106 = (_zz_dataOut_payload_0_10932 < _zz_dataOut_payload_0_10956);
  assign _zz_dataOut_payload_0_11107 = (_zz_dataOut_payload_0_11106 ? _zz_dataOut_payload_0_10932 : _zz_dataOut_payload_0_10956);
  assign _zz_dataOut_payload_0_11108 = (_zz_dataOut_payload_0_11106 ? _zz_dataOut_payload_0_10956 : _zz_dataOut_payload_0_10932);
  assign _zz_dataOut_payload_0_11109 = (_zz_dataOut_payload_0_10935 < _zz_dataOut_payload_0_10959);
  assign _zz_dataOut_payload_0_11110 = (_zz_dataOut_payload_0_11109 ? _zz_dataOut_payload_0_10935 : _zz_dataOut_payload_0_10959);
  assign _zz_dataOut_payload_0_11111 = (_zz_dataOut_payload_0_11109 ? _zz_dataOut_payload_0_10959 : _zz_dataOut_payload_0_10935);
  assign _zz_dataOut_payload_0_11112 = (_zz_dataOut_payload_0_11089 < _zz_dataOut_payload_0_11101);
  assign _zz_dataOut_payload_0_11113 = (_zz_dataOut_payload_0_11112 ? _zz_dataOut_payload_0_11089 : _zz_dataOut_payload_0_11101);
  assign _zz_dataOut_payload_0_11114 = (_zz_dataOut_payload_0_11112 ? _zz_dataOut_payload_0_11101 : _zz_dataOut_payload_0_11089);
  assign _zz_dataOut_payload_0_11115 = (_zz_dataOut_payload_0_11092 < _zz_dataOut_payload_0_11104);
  assign _zz_dataOut_payload_0_11116 = (_zz_dataOut_payload_0_11115 ? _zz_dataOut_payload_0_11092 : _zz_dataOut_payload_0_11104);
  assign _zz_dataOut_payload_0_11117 = (_zz_dataOut_payload_0_11115 ? _zz_dataOut_payload_0_11104 : _zz_dataOut_payload_0_11092);
  assign _zz_dataOut_payload_0_11118 = (_zz_dataOut_payload_0_11095 < _zz_dataOut_payload_0_11107);
  assign _zz_dataOut_payload_0_11119 = (_zz_dataOut_payload_0_11118 ? _zz_dataOut_payload_0_11095 : _zz_dataOut_payload_0_11107);
  assign _zz_dataOut_payload_0_11120 = (_zz_dataOut_payload_0_11118 ? _zz_dataOut_payload_0_11107 : _zz_dataOut_payload_0_11095);
  assign _zz_dataOut_payload_0_11121 = (_zz_dataOut_payload_0_11098 < _zz_dataOut_payload_0_11110);
  assign _zz_dataOut_payload_0_11122 = (_zz_dataOut_payload_0_11121 ? _zz_dataOut_payload_0_11098 : _zz_dataOut_payload_0_11110);
  assign _zz_dataOut_payload_0_11123 = (_zz_dataOut_payload_0_11121 ? _zz_dataOut_payload_0_11110 : _zz_dataOut_payload_0_11098);
  assign _zz_dataOut_payload_0_11124 = (_zz_dataOut_payload_0_11113 < _zz_dataOut_payload_0_11119);
  assign _zz_dataOut_payload_0_11125 = (_zz_dataOut_payload_0_11124 ? _zz_dataOut_payload_0_11113 : _zz_dataOut_payload_0_11119);
  assign _zz_dataOut_payload_0_11126 = (_zz_dataOut_payload_0_11124 ? _zz_dataOut_payload_0_11119 : _zz_dataOut_payload_0_11113);
  assign _zz_dataOut_payload_0_11127 = (_zz_dataOut_payload_0_11116 < _zz_dataOut_payload_0_11122);
  assign _zz_dataOut_payload_0_11128 = (_zz_dataOut_payload_0_11127 ? _zz_dataOut_payload_0_11116 : _zz_dataOut_payload_0_11122);
  assign _zz_dataOut_payload_0_11129 = (_zz_dataOut_payload_0_11127 ? _zz_dataOut_payload_0_11122 : _zz_dataOut_payload_0_11116);
  assign _zz_dataOut_payload_0_11130 = (_zz_dataOut_payload_0_11125 < _zz_dataOut_payload_0_11128);
  assign _zz_dataOut_payload_0_11131 = (_zz_dataOut_payload_0_11126 < _zz_dataOut_payload_0_11129);
  assign _zz_dataOut_payload_0_11136 = (_zz_dataOut_payload_0_11114 < _zz_dataOut_payload_0_11120);
  assign _zz_dataOut_payload_0_11137 = (_zz_dataOut_payload_0_11136 ? _zz_dataOut_payload_0_11114 : _zz_dataOut_payload_0_11120);
  assign _zz_dataOut_payload_0_11138 = (_zz_dataOut_payload_0_11136 ? _zz_dataOut_payload_0_11120 : _zz_dataOut_payload_0_11114);
  assign _zz_dataOut_payload_0_11139 = (_zz_dataOut_payload_0_11117 < _zz_dataOut_payload_0_11123);
  assign _zz_dataOut_payload_0_11140 = (_zz_dataOut_payload_0_11139 ? _zz_dataOut_payload_0_11117 : _zz_dataOut_payload_0_11123);
  assign _zz_dataOut_payload_0_11141 = (_zz_dataOut_payload_0_11139 ? _zz_dataOut_payload_0_11123 : _zz_dataOut_payload_0_11117);
  assign _zz_dataOut_payload_0_11142 = (_zz_dataOut_payload_0_11137 < _zz_dataOut_payload_0_11140);
  assign _zz_dataOut_payload_0_11143 = (_zz_dataOut_payload_0_11138 < _zz_dataOut_payload_0_11141);
  assign _zz_dataOut_payload_0_11156 = (_zz_dataOut_payload_0_11090 < _zz_dataOut_payload_0_11102);
  assign _zz_dataOut_payload_0_11157 = (_zz_dataOut_payload_0_11156 ? _zz_dataOut_payload_0_11090 : _zz_dataOut_payload_0_11102);
  assign _zz_dataOut_payload_0_11158 = (_zz_dataOut_payload_0_11156 ? _zz_dataOut_payload_0_11102 : _zz_dataOut_payload_0_11090);
  assign _zz_dataOut_payload_0_11159 = (_zz_dataOut_payload_0_11093 < _zz_dataOut_payload_0_11105);
  assign _zz_dataOut_payload_0_11160 = (_zz_dataOut_payload_0_11159 ? _zz_dataOut_payload_0_11093 : _zz_dataOut_payload_0_11105);
  assign _zz_dataOut_payload_0_11161 = (_zz_dataOut_payload_0_11159 ? _zz_dataOut_payload_0_11105 : _zz_dataOut_payload_0_11093);
  assign _zz_dataOut_payload_0_11162 = (_zz_dataOut_payload_0_11096 < _zz_dataOut_payload_0_11108);
  assign _zz_dataOut_payload_0_11163 = (_zz_dataOut_payload_0_11162 ? _zz_dataOut_payload_0_11096 : _zz_dataOut_payload_0_11108);
  assign _zz_dataOut_payload_0_11164 = (_zz_dataOut_payload_0_11162 ? _zz_dataOut_payload_0_11108 : _zz_dataOut_payload_0_11096);
  assign _zz_dataOut_payload_0_11165 = (_zz_dataOut_payload_0_11099 < _zz_dataOut_payload_0_11111);
  assign _zz_dataOut_payload_0_11166 = (_zz_dataOut_payload_0_11165 ? _zz_dataOut_payload_0_11099 : _zz_dataOut_payload_0_11111);
  assign _zz_dataOut_payload_0_11167 = (_zz_dataOut_payload_0_11165 ? _zz_dataOut_payload_0_11111 : _zz_dataOut_payload_0_11099);
  assign _zz_dataOut_payload_0_11168 = (_zz_dataOut_payload_0_11157 < _zz_dataOut_payload_0_11163);
  assign _zz_dataOut_payload_0_11169 = (_zz_dataOut_payload_0_11168 ? _zz_dataOut_payload_0_11157 : _zz_dataOut_payload_0_11163);
  assign _zz_dataOut_payload_0_11170 = (_zz_dataOut_payload_0_11168 ? _zz_dataOut_payload_0_11163 : _zz_dataOut_payload_0_11157);
  assign _zz_dataOut_payload_0_11171 = (_zz_dataOut_payload_0_11160 < _zz_dataOut_payload_0_11166);
  assign _zz_dataOut_payload_0_11172 = (_zz_dataOut_payload_0_11171 ? _zz_dataOut_payload_0_11160 : _zz_dataOut_payload_0_11166);
  assign _zz_dataOut_payload_0_11173 = (_zz_dataOut_payload_0_11171 ? _zz_dataOut_payload_0_11166 : _zz_dataOut_payload_0_11160);
  assign _zz_dataOut_payload_0_11174 = (_zz_dataOut_payload_0_11169 < _zz_dataOut_payload_0_11172);
  assign _zz_dataOut_payload_0_11175 = (_zz_dataOut_payload_0_11170 < _zz_dataOut_payload_0_11173);
  assign _zz_dataOut_payload_0_11180 = (_zz_dataOut_payload_0_11158 < _zz_dataOut_payload_0_11164);
  assign _zz_dataOut_payload_0_11181 = (_zz_dataOut_payload_0_11180 ? _zz_dataOut_payload_0_11158 : _zz_dataOut_payload_0_11164);
  assign _zz_dataOut_payload_0_11182 = (_zz_dataOut_payload_0_11180 ? _zz_dataOut_payload_0_11164 : _zz_dataOut_payload_0_11158);
  assign _zz_dataOut_payload_0_11183 = (_zz_dataOut_payload_0_11161 < _zz_dataOut_payload_0_11167);
  assign _zz_dataOut_payload_0_11184 = (_zz_dataOut_payload_0_11183 ? _zz_dataOut_payload_0_11161 : _zz_dataOut_payload_0_11167);
  assign _zz_dataOut_payload_0_11185 = (_zz_dataOut_payload_0_11183 ? _zz_dataOut_payload_0_11167 : _zz_dataOut_payload_0_11161);
  assign _zz_dataOut_payload_0_11186 = (_zz_dataOut_payload_0_11181 < _zz_dataOut_payload_0_11184);
  assign _zz_dataOut_payload_0_11187 = (_zz_dataOut_payload_0_11182 < _zz_dataOut_payload_0_11185);
  assign _zz_dataOut_payload_0_11248 = (_zz_dataOut_payload_0_10911 < _zz_dataOut_payload_0_10863);
  assign _zz_dataOut_payload_0_11249 = (_zz_dataOut_payload_0_11248 ? _zz_dataOut_payload_0_10911 : _zz_dataOut_payload_0_10863);
  assign _zz_dataOut_payload_0_11250 = (_zz_dataOut_payload_0_11248 ? _zz_dataOut_payload_0_10863 : _zz_dataOut_payload_0_10911);
  assign _zz_dataOut_payload_0_11251 = (_zz_dataOut_payload_0_10908 < _zz_dataOut_payload_0_10860);
  assign _zz_dataOut_payload_0_11252 = (_zz_dataOut_payload_0_11251 ? _zz_dataOut_payload_0_10908 : _zz_dataOut_payload_0_10860);
  assign _zz_dataOut_payload_0_11253 = (_zz_dataOut_payload_0_11251 ? _zz_dataOut_payload_0_10860 : _zz_dataOut_payload_0_10908);
  assign _zz_dataOut_payload_0_11254 = (_zz_dataOut_payload_0_10905 < _zz_dataOut_payload_0_10857);
  assign _zz_dataOut_payload_0_11255 = (_zz_dataOut_payload_0_11254 ? _zz_dataOut_payload_0_10905 : _zz_dataOut_payload_0_10857);
  assign _zz_dataOut_payload_0_11256 = (_zz_dataOut_payload_0_11254 ? _zz_dataOut_payload_0_10857 : _zz_dataOut_payload_0_10905);
  assign _zz_dataOut_payload_0_11257 = (_zz_dataOut_payload_0_10902 < _zz_dataOut_payload_0_10854);
  assign _zz_dataOut_payload_0_11258 = (_zz_dataOut_payload_0_11257 ? _zz_dataOut_payload_0_10902 : _zz_dataOut_payload_0_10854);
  assign _zz_dataOut_payload_0_11259 = (_zz_dataOut_payload_0_11257 ? _zz_dataOut_payload_0_10854 : _zz_dataOut_payload_0_10902);
  assign _zz_dataOut_payload_0_11260 = (_zz_dataOut_payload_0_10899 < _zz_dataOut_payload_0_10851);
  assign _zz_dataOut_payload_0_11261 = (_zz_dataOut_payload_0_11260 ? _zz_dataOut_payload_0_10899 : _zz_dataOut_payload_0_10851);
  assign _zz_dataOut_payload_0_11262 = (_zz_dataOut_payload_0_11260 ? _zz_dataOut_payload_0_10851 : _zz_dataOut_payload_0_10899);
  assign _zz_dataOut_payload_0_11263 = (_zz_dataOut_payload_0_10896 < _zz_dataOut_payload_0_10848);
  assign _zz_dataOut_payload_0_11264 = (_zz_dataOut_payload_0_11263 ? _zz_dataOut_payload_0_10896 : _zz_dataOut_payload_0_10848);
  assign _zz_dataOut_payload_0_11265 = (_zz_dataOut_payload_0_11263 ? _zz_dataOut_payload_0_10848 : _zz_dataOut_payload_0_10896);
  assign _zz_dataOut_payload_0_11266 = (_zz_dataOut_payload_0_10893 < _zz_dataOut_payload_0_10845);
  assign _zz_dataOut_payload_0_11267 = (_zz_dataOut_payload_0_11266 ? _zz_dataOut_payload_0_10893 : _zz_dataOut_payload_0_10845);
  assign _zz_dataOut_payload_0_11268 = (_zz_dataOut_payload_0_11266 ? _zz_dataOut_payload_0_10845 : _zz_dataOut_payload_0_10893);
  assign _zz_dataOut_payload_0_11269 = (_zz_dataOut_payload_0_10890 < _zz_dataOut_payload_0_10842);
  assign _zz_dataOut_payload_0_11270 = (_zz_dataOut_payload_0_11269 ? _zz_dataOut_payload_0_10890 : _zz_dataOut_payload_0_10842);
  assign _zz_dataOut_payload_0_11271 = (_zz_dataOut_payload_0_11269 ? _zz_dataOut_payload_0_10842 : _zz_dataOut_payload_0_10890);
  assign _zz_dataOut_payload_0_11272 = (_zz_dataOut_payload_0_10887 < _zz_dataOut_payload_0_10839);
  assign _zz_dataOut_payload_0_11273 = (_zz_dataOut_payload_0_11272 ? _zz_dataOut_payload_0_10887 : _zz_dataOut_payload_0_10839);
  assign _zz_dataOut_payload_0_11274 = (_zz_dataOut_payload_0_11272 ? _zz_dataOut_payload_0_10839 : _zz_dataOut_payload_0_10887);
  assign _zz_dataOut_payload_0_11275 = (_zz_dataOut_payload_0_10884 < _zz_dataOut_payload_0_10836);
  assign _zz_dataOut_payload_0_11276 = (_zz_dataOut_payload_0_11275 ? _zz_dataOut_payload_0_10884 : _zz_dataOut_payload_0_10836);
  assign _zz_dataOut_payload_0_11277 = (_zz_dataOut_payload_0_11275 ? _zz_dataOut_payload_0_10836 : _zz_dataOut_payload_0_10884);
  assign _zz_dataOut_payload_0_11278 = (_zz_dataOut_payload_0_10881 < _zz_dataOut_payload_0_10833);
  assign _zz_dataOut_payload_0_11279 = (_zz_dataOut_payload_0_11278 ? _zz_dataOut_payload_0_10881 : _zz_dataOut_payload_0_10833);
  assign _zz_dataOut_payload_0_11280 = (_zz_dataOut_payload_0_11278 ? _zz_dataOut_payload_0_10833 : _zz_dataOut_payload_0_10881);
  assign _zz_dataOut_payload_0_11281 = (_zz_dataOut_payload_0_10878 < _zz_dataOut_payload_0_10830);
  assign _zz_dataOut_payload_0_11282 = (_zz_dataOut_payload_0_11281 ? _zz_dataOut_payload_0_10878 : _zz_dataOut_payload_0_10830);
  assign _zz_dataOut_payload_0_11283 = (_zz_dataOut_payload_0_11281 ? _zz_dataOut_payload_0_10830 : _zz_dataOut_payload_0_10878);
  assign _zz_dataOut_payload_0_11284 = (_zz_dataOut_payload_0_10875 < _zz_dataOut_payload_0_10827);
  assign _zz_dataOut_payload_0_11285 = (_zz_dataOut_payload_0_11284 ? _zz_dataOut_payload_0_10875 : _zz_dataOut_payload_0_10827);
  assign _zz_dataOut_payload_0_11286 = (_zz_dataOut_payload_0_11284 ? _zz_dataOut_payload_0_10827 : _zz_dataOut_payload_0_10875);
  assign _zz_dataOut_payload_0_11287 = (_zz_dataOut_payload_0_10872 < _zz_dataOut_payload_0_10824);
  assign _zz_dataOut_payload_0_11288 = (_zz_dataOut_payload_0_11287 ? _zz_dataOut_payload_0_10872 : _zz_dataOut_payload_0_10824);
  assign _zz_dataOut_payload_0_11289 = (_zz_dataOut_payload_0_11287 ? _zz_dataOut_payload_0_10824 : _zz_dataOut_payload_0_10872);
  assign _zz_dataOut_payload_0_11290 = (_zz_dataOut_payload_0_10869 < _zz_dataOut_payload_0_10821);
  assign _zz_dataOut_payload_0_11291 = (_zz_dataOut_payload_0_11290 ? _zz_dataOut_payload_0_10869 : _zz_dataOut_payload_0_10821);
  assign _zz_dataOut_payload_0_11292 = (_zz_dataOut_payload_0_11290 ? _zz_dataOut_payload_0_10821 : _zz_dataOut_payload_0_10869);
  assign _zz_dataOut_payload_0_11293 = (_zz_dataOut_payload_0_10866 < _zz_dataOut_payload_0_10818);
  assign _zz_dataOut_payload_0_11294 = (_zz_dataOut_payload_0_11293 ? _zz_dataOut_payload_0_10866 : _zz_dataOut_payload_0_10818);
  assign _zz_dataOut_payload_0_11295 = (_zz_dataOut_payload_0_11293 ? _zz_dataOut_payload_0_10818 : _zz_dataOut_payload_0_10866);
  assign _zz_dataOut_payload_0_11296 = (_zz_dataOut_payload_0_11249 < _zz_dataOut_payload_0_11273);
  assign _zz_dataOut_payload_0_11297 = (_zz_dataOut_payload_0_11296 ? _zz_dataOut_payload_0_11249 : _zz_dataOut_payload_0_11273);
  assign _zz_dataOut_payload_0_11298 = (_zz_dataOut_payload_0_11296 ? _zz_dataOut_payload_0_11273 : _zz_dataOut_payload_0_11249);
  assign _zz_dataOut_payload_0_11299 = (_zz_dataOut_payload_0_11252 < _zz_dataOut_payload_0_11276);
  assign _zz_dataOut_payload_0_11300 = (_zz_dataOut_payload_0_11299 ? _zz_dataOut_payload_0_11252 : _zz_dataOut_payload_0_11276);
  assign _zz_dataOut_payload_0_11301 = (_zz_dataOut_payload_0_11299 ? _zz_dataOut_payload_0_11276 : _zz_dataOut_payload_0_11252);
  assign _zz_dataOut_payload_0_11302 = (_zz_dataOut_payload_0_11255 < _zz_dataOut_payload_0_11279);
  assign _zz_dataOut_payload_0_11303 = (_zz_dataOut_payload_0_11302 ? _zz_dataOut_payload_0_11255 : _zz_dataOut_payload_0_11279);
  assign _zz_dataOut_payload_0_11304 = (_zz_dataOut_payload_0_11302 ? _zz_dataOut_payload_0_11279 : _zz_dataOut_payload_0_11255);
  assign _zz_dataOut_payload_0_11305 = (_zz_dataOut_payload_0_11258 < _zz_dataOut_payload_0_11282);
  assign _zz_dataOut_payload_0_11306 = (_zz_dataOut_payload_0_11305 ? _zz_dataOut_payload_0_11258 : _zz_dataOut_payload_0_11282);
  assign _zz_dataOut_payload_0_11307 = (_zz_dataOut_payload_0_11305 ? _zz_dataOut_payload_0_11282 : _zz_dataOut_payload_0_11258);
  assign _zz_dataOut_payload_0_11308 = (_zz_dataOut_payload_0_11261 < _zz_dataOut_payload_0_11285);
  assign _zz_dataOut_payload_0_11309 = (_zz_dataOut_payload_0_11308 ? _zz_dataOut_payload_0_11261 : _zz_dataOut_payload_0_11285);
  assign _zz_dataOut_payload_0_11310 = (_zz_dataOut_payload_0_11308 ? _zz_dataOut_payload_0_11285 : _zz_dataOut_payload_0_11261);
  assign _zz_dataOut_payload_0_11311 = (_zz_dataOut_payload_0_11264 < _zz_dataOut_payload_0_11288);
  assign _zz_dataOut_payload_0_11312 = (_zz_dataOut_payload_0_11311 ? _zz_dataOut_payload_0_11264 : _zz_dataOut_payload_0_11288);
  assign _zz_dataOut_payload_0_11313 = (_zz_dataOut_payload_0_11311 ? _zz_dataOut_payload_0_11288 : _zz_dataOut_payload_0_11264);
  assign _zz_dataOut_payload_0_11314 = (_zz_dataOut_payload_0_11267 < _zz_dataOut_payload_0_11291);
  assign _zz_dataOut_payload_0_11315 = (_zz_dataOut_payload_0_11314 ? _zz_dataOut_payload_0_11267 : _zz_dataOut_payload_0_11291);
  assign _zz_dataOut_payload_0_11316 = (_zz_dataOut_payload_0_11314 ? _zz_dataOut_payload_0_11291 : _zz_dataOut_payload_0_11267);
  assign _zz_dataOut_payload_0_11317 = (_zz_dataOut_payload_0_11270 < _zz_dataOut_payload_0_11294);
  assign _zz_dataOut_payload_0_11318 = (_zz_dataOut_payload_0_11317 ? _zz_dataOut_payload_0_11270 : _zz_dataOut_payload_0_11294);
  assign _zz_dataOut_payload_0_11319 = (_zz_dataOut_payload_0_11317 ? _zz_dataOut_payload_0_11294 : _zz_dataOut_payload_0_11270);
  assign _zz_dataOut_payload_0_11320 = (_zz_dataOut_payload_0_11297 < _zz_dataOut_payload_0_11309);
  assign _zz_dataOut_payload_0_11321 = (_zz_dataOut_payload_0_11320 ? _zz_dataOut_payload_0_11297 : _zz_dataOut_payload_0_11309);
  assign _zz_dataOut_payload_0_11322 = (_zz_dataOut_payload_0_11320 ? _zz_dataOut_payload_0_11309 : _zz_dataOut_payload_0_11297);
  assign _zz_dataOut_payload_0_11323 = (_zz_dataOut_payload_0_11300 < _zz_dataOut_payload_0_11312);
  assign _zz_dataOut_payload_0_11324 = (_zz_dataOut_payload_0_11323 ? _zz_dataOut_payload_0_11300 : _zz_dataOut_payload_0_11312);
  assign _zz_dataOut_payload_0_11325 = (_zz_dataOut_payload_0_11323 ? _zz_dataOut_payload_0_11312 : _zz_dataOut_payload_0_11300);
  assign _zz_dataOut_payload_0_11326 = (_zz_dataOut_payload_0_11303 < _zz_dataOut_payload_0_11315);
  assign _zz_dataOut_payload_0_11327 = (_zz_dataOut_payload_0_11326 ? _zz_dataOut_payload_0_11303 : _zz_dataOut_payload_0_11315);
  assign _zz_dataOut_payload_0_11328 = (_zz_dataOut_payload_0_11326 ? _zz_dataOut_payload_0_11315 : _zz_dataOut_payload_0_11303);
  assign _zz_dataOut_payload_0_11329 = (_zz_dataOut_payload_0_11306 < _zz_dataOut_payload_0_11318);
  assign _zz_dataOut_payload_0_11330 = (_zz_dataOut_payload_0_11329 ? _zz_dataOut_payload_0_11306 : _zz_dataOut_payload_0_11318);
  assign _zz_dataOut_payload_0_11331 = (_zz_dataOut_payload_0_11329 ? _zz_dataOut_payload_0_11318 : _zz_dataOut_payload_0_11306);
  assign _zz_dataOut_payload_0_11332 = (_zz_dataOut_payload_0_11321 < _zz_dataOut_payload_0_11327);
  assign _zz_dataOut_payload_0_11333 = (_zz_dataOut_payload_0_11332 ? _zz_dataOut_payload_0_11321 : _zz_dataOut_payload_0_11327);
  assign _zz_dataOut_payload_0_11334 = (_zz_dataOut_payload_0_11332 ? _zz_dataOut_payload_0_11327 : _zz_dataOut_payload_0_11321);
  assign _zz_dataOut_payload_0_11335 = (_zz_dataOut_payload_0_11324 < _zz_dataOut_payload_0_11330);
  assign _zz_dataOut_payload_0_11336 = (_zz_dataOut_payload_0_11335 ? _zz_dataOut_payload_0_11324 : _zz_dataOut_payload_0_11330);
  assign _zz_dataOut_payload_0_11337 = (_zz_dataOut_payload_0_11335 ? _zz_dataOut_payload_0_11330 : _zz_dataOut_payload_0_11324);
  assign _zz_dataOut_payload_0_11338 = (_zz_dataOut_payload_0_11333 < _zz_dataOut_payload_0_11336);
  assign _zz_dataOut_payload_0_11339 = (_zz_dataOut_payload_0_11334 < _zz_dataOut_payload_0_11337);
  assign _zz_dataOut_payload_0_11344 = (_zz_dataOut_payload_0_11322 < _zz_dataOut_payload_0_11328);
  assign _zz_dataOut_payload_0_11345 = (_zz_dataOut_payload_0_11344 ? _zz_dataOut_payload_0_11322 : _zz_dataOut_payload_0_11328);
  assign _zz_dataOut_payload_0_11346 = (_zz_dataOut_payload_0_11344 ? _zz_dataOut_payload_0_11328 : _zz_dataOut_payload_0_11322);
  assign _zz_dataOut_payload_0_11347 = (_zz_dataOut_payload_0_11325 < _zz_dataOut_payload_0_11331);
  assign _zz_dataOut_payload_0_11348 = (_zz_dataOut_payload_0_11347 ? _zz_dataOut_payload_0_11325 : _zz_dataOut_payload_0_11331);
  assign _zz_dataOut_payload_0_11349 = (_zz_dataOut_payload_0_11347 ? _zz_dataOut_payload_0_11331 : _zz_dataOut_payload_0_11325);
  assign _zz_dataOut_payload_0_11350 = (_zz_dataOut_payload_0_11345 < _zz_dataOut_payload_0_11348);
  assign _zz_dataOut_payload_0_11351 = (_zz_dataOut_payload_0_11346 < _zz_dataOut_payload_0_11349);
  assign _zz_dataOut_payload_0_11364 = (_zz_dataOut_payload_0_11298 < _zz_dataOut_payload_0_11310);
  assign _zz_dataOut_payload_0_11365 = (_zz_dataOut_payload_0_11364 ? _zz_dataOut_payload_0_11298 : _zz_dataOut_payload_0_11310);
  assign _zz_dataOut_payload_0_11366 = (_zz_dataOut_payload_0_11364 ? _zz_dataOut_payload_0_11310 : _zz_dataOut_payload_0_11298);
  assign _zz_dataOut_payload_0_11367 = (_zz_dataOut_payload_0_11301 < _zz_dataOut_payload_0_11313);
  assign _zz_dataOut_payload_0_11368 = (_zz_dataOut_payload_0_11367 ? _zz_dataOut_payload_0_11301 : _zz_dataOut_payload_0_11313);
  assign _zz_dataOut_payload_0_11369 = (_zz_dataOut_payload_0_11367 ? _zz_dataOut_payload_0_11313 : _zz_dataOut_payload_0_11301);
  assign _zz_dataOut_payload_0_11370 = (_zz_dataOut_payload_0_11304 < _zz_dataOut_payload_0_11316);
  assign _zz_dataOut_payload_0_11371 = (_zz_dataOut_payload_0_11370 ? _zz_dataOut_payload_0_11304 : _zz_dataOut_payload_0_11316);
  assign _zz_dataOut_payload_0_11372 = (_zz_dataOut_payload_0_11370 ? _zz_dataOut_payload_0_11316 : _zz_dataOut_payload_0_11304);
  assign _zz_dataOut_payload_0_11373 = (_zz_dataOut_payload_0_11307 < _zz_dataOut_payload_0_11319);
  assign _zz_dataOut_payload_0_11374 = (_zz_dataOut_payload_0_11373 ? _zz_dataOut_payload_0_11307 : _zz_dataOut_payload_0_11319);
  assign _zz_dataOut_payload_0_11375 = (_zz_dataOut_payload_0_11373 ? _zz_dataOut_payload_0_11319 : _zz_dataOut_payload_0_11307);
  assign _zz_dataOut_payload_0_11376 = (_zz_dataOut_payload_0_11365 < _zz_dataOut_payload_0_11371);
  assign _zz_dataOut_payload_0_11377 = (_zz_dataOut_payload_0_11376 ? _zz_dataOut_payload_0_11365 : _zz_dataOut_payload_0_11371);
  assign _zz_dataOut_payload_0_11378 = (_zz_dataOut_payload_0_11376 ? _zz_dataOut_payload_0_11371 : _zz_dataOut_payload_0_11365);
  assign _zz_dataOut_payload_0_11379 = (_zz_dataOut_payload_0_11368 < _zz_dataOut_payload_0_11374);
  assign _zz_dataOut_payload_0_11380 = (_zz_dataOut_payload_0_11379 ? _zz_dataOut_payload_0_11368 : _zz_dataOut_payload_0_11374);
  assign _zz_dataOut_payload_0_11381 = (_zz_dataOut_payload_0_11379 ? _zz_dataOut_payload_0_11374 : _zz_dataOut_payload_0_11368);
  assign _zz_dataOut_payload_0_11382 = (_zz_dataOut_payload_0_11377 < _zz_dataOut_payload_0_11380);
  assign _zz_dataOut_payload_0_11383 = (_zz_dataOut_payload_0_11378 < _zz_dataOut_payload_0_11381);
  assign _zz_dataOut_payload_0_11388 = (_zz_dataOut_payload_0_11366 < _zz_dataOut_payload_0_11372);
  assign _zz_dataOut_payload_0_11389 = (_zz_dataOut_payload_0_11388 ? _zz_dataOut_payload_0_11366 : _zz_dataOut_payload_0_11372);
  assign _zz_dataOut_payload_0_11390 = (_zz_dataOut_payload_0_11388 ? _zz_dataOut_payload_0_11372 : _zz_dataOut_payload_0_11366);
  assign _zz_dataOut_payload_0_11391 = (_zz_dataOut_payload_0_11369 < _zz_dataOut_payload_0_11375);
  assign _zz_dataOut_payload_0_11392 = (_zz_dataOut_payload_0_11391 ? _zz_dataOut_payload_0_11369 : _zz_dataOut_payload_0_11375);
  assign _zz_dataOut_payload_0_11393 = (_zz_dataOut_payload_0_11391 ? _zz_dataOut_payload_0_11375 : _zz_dataOut_payload_0_11369);
  assign _zz_dataOut_payload_0_11394 = (_zz_dataOut_payload_0_11389 < _zz_dataOut_payload_0_11392);
  assign _zz_dataOut_payload_0_11395 = (_zz_dataOut_payload_0_11390 < _zz_dataOut_payload_0_11393);
  assign _zz_dataOut_payload_0_11424 = (_zz_dataOut_payload_0_11250 < _zz_dataOut_payload_0_11274);
  assign _zz_dataOut_payload_0_11425 = (_zz_dataOut_payload_0_11424 ? _zz_dataOut_payload_0_11250 : _zz_dataOut_payload_0_11274);
  assign _zz_dataOut_payload_0_11426 = (_zz_dataOut_payload_0_11424 ? _zz_dataOut_payload_0_11274 : _zz_dataOut_payload_0_11250);
  assign _zz_dataOut_payload_0_11427 = (_zz_dataOut_payload_0_11253 < _zz_dataOut_payload_0_11277);
  assign _zz_dataOut_payload_0_11428 = (_zz_dataOut_payload_0_11427 ? _zz_dataOut_payload_0_11253 : _zz_dataOut_payload_0_11277);
  assign _zz_dataOut_payload_0_11429 = (_zz_dataOut_payload_0_11427 ? _zz_dataOut_payload_0_11277 : _zz_dataOut_payload_0_11253);
  assign _zz_dataOut_payload_0_11430 = (_zz_dataOut_payload_0_11256 < _zz_dataOut_payload_0_11280);
  assign _zz_dataOut_payload_0_11431 = (_zz_dataOut_payload_0_11430 ? _zz_dataOut_payload_0_11256 : _zz_dataOut_payload_0_11280);
  assign _zz_dataOut_payload_0_11432 = (_zz_dataOut_payload_0_11430 ? _zz_dataOut_payload_0_11280 : _zz_dataOut_payload_0_11256);
  assign _zz_dataOut_payload_0_11433 = (_zz_dataOut_payload_0_11259 < _zz_dataOut_payload_0_11283);
  assign _zz_dataOut_payload_0_11434 = (_zz_dataOut_payload_0_11433 ? _zz_dataOut_payload_0_11259 : _zz_dataOut_payload_0_11283);
  assign _zz_dataOut_payload_0_11435 = (_zz_dataOut_payload_0_11433 ? _zz_dataOut_payload_0_11283 : _zz_dataOut_payload_0_11259);
  assign _zz_dataOut_payload_0_11436 = (_zz_dataOut_payload_0_11262 < _zz_dataOut_payload_0_11286);
  assign _zz_dataOut_payload_0_11437 = (_zz_dataOut_payload_0_11436 ? _zz_dataOut_payload_0_11262 : _zz_dataOut_payload_0_11286);
  assign _zz_dataOut_payload_0_11438 = (_zz_dataOut_payload_0_11436 ? _zz_dataOut_payload_0_11286 : _zz_dataOut_payload_0_11262);
  assign _zz_dataOut_payload_0_11439 = (_zz_dataOut_payload_0_11265 < _zz_dataOut_payload_0_11289);
  assign _zz_dataOut_payload_0_11440 = (_zz_dataOut_payload_0_11439 ? _zz_dataOut_payload_0_11265 : _zz_dataOut_payload_0_11289);
  assign _zz_dataOut_payload_0_11441 = (_zz_dataOut_payload_0_11439 ? _zz_dataOut_payload_0_11289 : _zz_dataOut_payload_0_11265);
  assign _zz_dataOut_payload_0_11442 = (_zz_dataOut_payload_0_11268 < _zz_dataOut_payload_0_11292);
  assign _zz_dataOut_payload_0_11443 = (_zz_dataOut_payload_0_11442 ? _zz_dataOut_payload_0_11268 : _zz_dataOut_payload_0_11292);
  assign _zz_dataOut_payload_0_11444 = (_zz_dataOut_payload_0_11442 ? _zz_dataOut_payload_0_11292 : _zz_dataOut_payload_0_11268);
  assign _zz_dataOut_payload_0_11445 = (_zz_dataOut_payload_0_11271 < _zz_dataOut_payload_0_11295);
  assign _zz_dataOut_payload_0_11446 = (_zz_dataOut_payload_0_11445 ? _zz_dataOut_payload_0_11271 : _zz_dataOut_payload_0_11295);
  assign _zz_dataOut_payload_0_11447 = (_zz_dataOut_payload_0_11445 ? _zz_dataOut_payload_0_11295 : _zz_dataOut_payload_0_11271);
  assign _zz_dataOut_payload_0_11448 = (_zz_dataOut_payload_0_11425 < _zz_dataOut_payload_0_11437);
  assign _zz_dataOut_payload_0_11449 = (_zz_dataOut_payload_0_11448 ? _zz_dataOut_payload_0_11425 : _zz_dataOut_payload_0_11437);
  assign _zz_dataOut_payload_0_11450 = (_zz_dataOut_payload_0_11448 ? _zz_dataOut_payload_0_11437 : _zz_dataOut_payload_0_11425);
  assign _zz_dataOut_payload_0_11451 = (_zz_dataOut_payload_0_11428 < _zz_dataOut_payload_0_11440);
  assign _zz_dataOut_payload_0_11452 = (_zz_dataOut_payload_0_11451 ? _zz_dataOut_payload_0_11428 : _zz_dataOut_payload_0_11440);
  assign _zz_dataOut_payload_0_11453 = (_zz_dataOut_payload_0_11451 ? _zz_dataOut_payload_0_11440 : _zz_dataOut_payload_0_11428);
  assign _zz_dataOut_payload_0_11454 = (_zz_dataOut_payload_0_11431 < _zz_dataOut_payload_0_11443);
  assign _zz_dataOut_payload_0_11455 = (_zz_dataOut_payload_0_11454 ? _zz_dataOut_payload_0_11431 : _zz_dataOut_payload_0_11443);
  assign _zz_dataOut_payload_0_11456 = (_zz_dataOut_payload_0_11454 ? _zz_dataOut_payload_0_11443 : _zz_dataOut_payload_0_11431);
  assign _zz_dataOut_payload_0_11457 = (_zz_dataOut_payload_0_11434 < _zz_dataOut_payload_0_11446);
  assign _zz_dataOut_payload_0_11458 = (_zz_dataOut_payload_0_11457 ? _zz_dataOut_payload_0_11434 : _zz_dataOut_payload_0_11446);
  assign _zz_dataOut_payload_0_11459 = (_zz_dataOut_payload_0_11457 ? _zz_dataOut_payload_0_11446 : _zz_dataOut_payload_0_11434);
  assign _zz_dataOut_payload_0_11460 = (_zz_dataOut_payload_0_11449 < _zz_dataOut_payload_0_11455);
  assign _zz_dataOut_payload_0_11461 = (_zz_dataOut_payload_0_11460 ? _zz_dataOut_payload_0_11449 : _zz_dataOut_payload_0_11455);
  assign _zz_dataOut_payload_0_11462 = (_zz_dataOut_payload_0_11460 ? _zz_dataOut_payload_0_11455 : _zz_dataOut_payload_0_11449);
  assign _zz_dataOut_payload_0_11463 = (_zz_dataOut_payload_0_11452 < _zz_dataOut_payload_0_11458);
  assign _zz_dataOut_payload_0_11464 = (_zz_dataOut_payload_0_11463 ? _zz_dataOut_payload_0_11452 : _zz_dataOut_payload_0_11458);
  assign _zz_dataOut_payload_0_11465 = (_zz_dataOut_payload_0_11463 ? _zz_dataOut_payload_0_11458 : _zz_dataOut_payload_0_11452);
  assign _zz_dataOut_payload_0_11466 = (_zz_dataOut_payload_0_11461 < _zz_dataOut_payload_0_11464);
  assign _zz_dataOut_payload_0_11467 = (_zz_dataOut_payload_0_11462 < _zz_dataOut_payload_0_11465);
  assign _zz_dataOut_payload_0_11472 = (_zz_dataOut_payload_0_11450 < _zz_dataOut_payload_0_11456);
  assign _zz_dataOut_payload_0_11473 = (_zz_dataOut_payload_0_11472 ? _zz_dataOut_payload_0_11450 : _zz_dataOut_payload_0_11456);
  assign _zz_dataOut_payload_0_11474 = (_zz_dataOut_payload_0_11472 ? _zz_dataOut_payload_0_11456 : _zz_dataOut_payload_0_11450);
  assign _zz_dataOut_payload_0_11475 = (_zz_dataOut_payload_0_11453 < _zz_dataOut_payload_0_11459);
  assign _zz_dataOut_payload_0_11476 = (_zz_dataOut_payload_0_11475 ? _zz_dataOut_payload_0_11453 : _zz_dataOut_payload_0_11459);
  assign _zz_dataOut_payload_0_11477 = (_zz_dataOut_payload_0_11475 ? _zz_dataOut_payload_0_11459 : _zz_dataOut_payload_0_11453);
  assign _zz_dataOut_payload_0_11478 = (_zz_dataOut_payload_0_11473 < _zz_dataOut_payload_0_11476);
  assign _zz_dataOut_payload_0_11479 = (_zz_dataOut_payload_0_11474 < _zz_dataOut_payload_0_11477);
  assign _zz_dataOut_payload_0_11492 = (_zz_dataOut_payload_0_11426 < _zz_dataOut_payload_0_11438);
  assign _zz_dataOut_payload_0_11493 = (_zz_dataOut_payload_0_11492 ? _zz_dataOut_payload_0_11426 : _zz_dataOut_payload_0_11438);
  assign _zz_dataOut_payload_0_11494 = (_zz_dataOut_payload_0_11492 ? _zz_dataOut_payload_0_11438 : _zz_dataOut_payload_0_11426);
  assign _zz_dataOut_payload_0_11495 = (_zz_dataOut_payload_0_11429 < _zz_dataOut_payload_0_11441);
  assign _zz_dataOut_payload_0_11496 = (_zz_dataOut_payload_0_11495 ? _zz_dataOut_payload_0_11429 : _zz_dataOut_payload_0_11441);
  assign _zz_dataOut_payload_0_11497 = (_zz_dataOut_payload_0_11495 ? _zz_dataOut_payload_0_11441 : _zz_dataOut_payload_0_11429);
  assign _zz_dataOut_payload_0_11498 = (_zz_dataOut_payload_0_11432 < _zz_dataOut_payload_0_11444);
  assign _zz_dataOut_payload_0_11499 = (_zz_dataOut_payload_0_11498 ? _zz_dataOut_payload_0_11432 : _zz_dataOut_payload_0_11444);
  assign _zz_dataOut_payload_0_11500 = (_zz_dataOut_payload_0_11498 ? _zz_dataOut_payload_0_11444 : _zz_dataOut_payload_0_11432);
  assign _zz_dataOut_payload_0_11501 = (_zz_dataOut_payload_0_11435 < _zz_dataOut_payload_0_11447);
  assign _zz_dataOut_payload_0_11502 = (_zz_dataOut_payload_0_11501 ? _zz_dataOut_payload_0_11435 : _zz_dataOut_payload_0_11447);
  assign _zz_dataOut_payload_0_11503 = (_zz_dataOut_payload_0_11501 ? _zz_dataOut_payload_0_11447 : _zz_dataOut_payload_0_11435);
  assign _zz_dataOut_payload_0_11504 = (_zz_dataOut_payload_0_11493 < _zz_dataOut_payload_0_11499);
  assign _zz_dataOut_payload_0_11505 = (_zz_dataOut_payload_0_11504 ? _zz_dataOut_payload_0_11493 : _zz_dataOut_payload_0_11499);
  assign _zz_dataOut_payload_0_11506 = (_zz_dataOut_payload_0_11504 ? _zz_dataOut_payload_0_11499 : _zz_dataOut_payload_0_11493);
  assign _zz_dataOut_payload_0_11507 = (_zz_dataOut_payload_0_11496 < _zz_dataOut_payload_0_11502);
  assign _zz_dataOut_payload_0_11508 = (_zz_dataOut_payload_0_11507 ? _zz_dataOut_payload_0_11496 : _zz_dataOut_payload_0_11502);
  assign _zz_dataOut_payload_0_11509 = (_zz_dataOut_payload_0_11507 ? _zz_dataOut_payload_0_11502 : _zz_dataOut_payload_0_11496);
  assign _zz_dataOut_payload_0_11510 = (_zz_dataOut_payload_0_11505 < _zz_dataOut_payload_0_11508);
  assign _zz_dataOut_payload_0_11511 = (_zz_dataOut_payload_0_11506 < _zz_dataOut_payload_0_11509);
  assign _zz_dataOut_payload_0_11516 = (_zz_dataOut_payload_0_11494 < _zz_dataOut_payload_0_11500);
  assign _zz_dataOut_payload_0_11517 = (_zz_dataOut_payload_0_11516 ? _zz_dataOut_payload_0_11494 : _zz_dataOut_payload_0_11500);
  assign _zz_dataOut_payload_0_11518 = (_zz_dataOut_payload_0_11516 ? _zz_dataOut_payload_0_11500 : _zz_dataOut_payload_0_11494);
  assign _zz_dataOut_payload_0_11519 = (_zz_dataOut_payload_0_11497 < _zz_dataOut_payload_0_11503);
  assign _zz_dataOut_payload_0_11520 = (_zz_dataOut_payload_0_11519 ? _zz_dataOut_payload_0_11497 : _zz_dataOut_payload_0_11503);
  assign _zz_dataOut_payload_0_11521 = (_zz_dataOut_payload_0_11519 ? _zz_dataOut_payload_0_11503 : _zz_dataOut_payload_0_11497);
  assign _zz_dataOut_payload_0_11522 = (_zz_dataOut_payload_0_11517 < _zz_dataOut_payload_0_11520);
  assign _zz_dataOut_payload_0_11523 = (_zz_dataOut_payload_0_11518 < _zz_dataOut_payload_0_11521);
  assign _zz_dataOut_payload_0_11904 = (_zz_dataOut_payload_0_11648 < _zz_dataOut_payload_0_11775);
  assign _zz_dataOut_payload_0_11905 = (_zz_dataOut_payload_0_11904 ? _zz_dataOut_payload_0_11648 : _zz_dataOut_payload_0_11775);
  assign _zz_dataOut_payload_0_11906 = (_zz_dataOut_payload_0_11904 ? _zz_dataOut_payload_0_11775 : _zz_dataOut_payload_0_11648);
  assign _zz_dataOut_payload_0_11907 = (_zz_dataOut_payload_0_11649 < _zz_dataOut_payload_0_11774);
  assign _zz_dataOut_payload_0_11908 = (_zz_dataOut_payload_0_11907 ? _zz_dataOut_payload_0_11649 : _zz_dataOut_payload_0_11774);
  assign _zz_dataOut_payload_0_11909 = (_zz_dataOut_payload_0_11907 ? _zz_dataOut_payload_0_11774 : _zz_dataOut_payload_0_11649);
  assign _zz_dataOut_payload_0_11910 = (_zz_dataOut_payload_0_11650 < _zz_dataOut_payload_0_11773);
  assign _zz_dataOut_payload_0_11911 = (_zz_dataOut_payload_0_11910 ? _zz_dataOut_payload_0_11650 : _zz_dataOut_payload_0_11773);
  assign _zz_dataOut_payload_0_11912 = (_zz_dataOut_payload_0_11910 ? _zz_dataOut_payload_0_11773 : _zz_dataOut_payload_0_11650);
  assign _zz_dataOut_payload_0_11913 = (_zz_dataOut_payload_0_11651 < _zz_dataOut_payload_0_11772);
  assign _zz_dataOut_payload_0_11914 = (_zz_dataOut_payload_0_11913 ? _zz_dataOut_payload_0_11651 : _zz_dataOut_payload_0_11772);
  assign _zz_dataOut_payload_0_11915 = (_zz_dataOut_payload_0_11913 ? _zz_dataOut_payload_0_11772 : _zz_dataOut_payload_0_11651);
  assign _zz_dataOut_payload_0_11916 = (_zz_dataOut_payload_0_11652 < _zz_dataOut_payload_0_11771);
  assign _zz_dataOut_payload_0_11917 = (_zz_dataOut_payload_0_11916 ? _zz_dataOut_payload_0_11652 : _zz_dataOut_payload_0_11771);
  assign _zz_dataOut_payload_0_11918 = (_zz_dataOut_payload_0_11916 ? _zz_dataOut_payload_0_11771 : _zz_dataOut_payload_0_11652);
  assign _zz_dataOut_payload_0_11919 = (_zz_dataOut_payload_0_11653 < _zz_dataOut_payload_0_11770);
  assign _zz_dataOut_payload_0_11920 = (_zz_dataOut_payload_0_11919 ? _zz_dataOut_payload_0_11653 : _zz_dataOut_payload_0_11770);
  assign _zz_dataOut_payload_0_11921 = (_zz_dataOut_payload_0_11919 ? _zz_dataOut_payload_0_11770 : _zz_dataOut_payload_0_11653);
  assign _zz_dataOut_payload_0_11922 = (_zz_dataOut_payload_0_11654 < _zz_dataOut_payload_0_11769);
  assign _zz_dataOut_payload_0_11923 = (_zz_dataOut_payload_0_11922 ? _zz_dataOut_payload_0_11654 : _zz_dataOut_payload_0_11769);
  assign _zz_dataOut_payload_0_11924 = (_zz_dataOut_payload_0_11922 ? _zz_dataOut_payload_0_11769 : _zz_dataOut_payload_0_11654);
  assign _zz_dataOut_payload_0_11925 = (_zz_dataOut_payload_0_11655 < _zz_dataOut_payload_0_11768);
  assign _zz_dataOut_payload_0_11926 = (_zz_dataOut_payload_0_11925 ? _zz_dataOut_payload_0_11655 : _zz_dataOut_payload_0_11768);
  assign _zz_dataOut_payload_0_11927 = (_zz_dataOut_payload_0_11925 ? _zz_dataOut_payload_0_11768 : _zz_dataOut_payload_0_11655);
  assign _zz_dataOut_payload_0_11928 = (_zz_dataOut_payload_0_11656 < _zz_dataOut_payload_0_11767);
  assign _zz_dataOut_payload_0_11929 = (_zz_dataOut_payload_0_11928 ? _zz_dataOut_payload_0_11656 : _zz_dataOut_payload_0_11767);
  assign _zz_dataOut_payload_0_11930 = (_zz_dataOut_payload_0_11928 ? _zz_dataOut_payload_0_11767 : _zz_dataOut_payload_0_11656);
  assign _zz_dataOut_payload_0_11931 = (_zz_dataOut_payload_0_11657 < _zz_dataOut_payload_0_11766);
  assign _zz_dataOut_payload_0_11932 = (_zz_dataOut_payload_0_11931 ? _zz_dataOut_payload_0_11657 : _zz_dataOut_payload_0_11766);
  assign _zz_dataOut_payload_0_11933 = (_zz_dataOut_payload_0_11931 ? _zz_dataOut_payload_0_11766 : _zz_dataOut_payload_0_11657);
  assign _zz_dataOut_payload_0_11934 = (_zz_dataOut_payload_0_11658 < _zz_dataOut_payload_0_11765);
  assign _zz_dataOut_payload_0_11935 = (_zz_dataOut_payload_0_11934 ? _zz_dataOut_payload_0_11658 : _zz_dataOut_payload_0_11765);
  assign _zz_dataOut_payload_0_11936 = (_zz_dataOut_payload_0_11934 ? _zz_dataOut_payload_0_11765 : _zz_dataOut_payload_0_11658);
  assign _zz_dataOut_payload_0_11937 = (_zz_dataOut_payload_0_11659 < _zz_dataOut_payload_0_11764);
  assign _zz_dataOut_payload_0_11938 = (_zz_dataOut_payload_0_11937 ? _zz_dataOut_payload_0_11659 : _zz_dataOut_payload_0_11764);
  assign _zz_dataOut_payload_0_11939 = (_zz_dataOut_payload_0_11937 ? _zz_dataOut_payload_0_11764 : _zz_dataOut_payload_0_11659);
  assign _zz_dataOut_payload_0_11940 = (_zz_dataOut_payload_0_11660 < _zz_dataOut_payload_0_11763);
  assign _zz_dataOut_payload_0_11941 = (_zz_dataOut_payload_0_11940 ? _zz_dataOut_payload_0_11660 : _zz_dataOut_payload_0_11763);
  assign _zz_dataOut_payload_0_11942 = (_zz_dataOut_payload_0_11940 ? _zz_dataOut_payload_0_11763 : _zz_dataOut_payload_0_11660);
  assign _zz_dataOut_payload_0_11943 = (_zz_dataOut_payload_0_11661 < _zz_dataOut_payload_0_11762);
  assign _zz_dataOut_payload_0_11944 = (_zz_dataOut_payload_0_11943 ? _zz_dataOut_payload_0_11661 : _zz_dataOut_payload_0_11762);
  assign _zz_dataOut_payload_0_11945 = (_zz_dataOut_payload_0_11943 ? _zz_dataOut_payload_0_11762 : _zz_dataOut_payload_0_11661);
  assign _zz_dataOut_payload_0_11946 = (_zz_dataOut_payload_0_11662 < _zz_dataOut_payload_0_11761);
  assign _zz_dataOut_payload_0_11947 = (_zz_dataOut_payload_0_11946 ? _zz_dataOut_payload_0_11662 : _zz_dataOut_payload_0_11761);
  assign _zz_dataOut_payload_0_11948 = (_zz_dataOut_payload_0_11946 ? _zz_dataOut_payload_0_11761 : _zz_dataOut_payload_0_11662);
  assign _zz_dataOut_payload_0_11949 = (_zz_dataOut_payload_0_11663 < _zz_dataOut_payload_0_11760);
  assign _zz_dataOut_payload_0_11950 = (_zz_dataOut_payload_0_11949 ? _zz_dataOut_payload_0_11663 : _zz_dataOut_payload_0_11760);
  assign _zz_dataOut_payload_0_11951 = (_zz_dataOut_payload_0_11949 ? _zz_dataOut_payload_0_11760 : _zz_dataOut_payload_0_11663);
  assign _zz_dataOut_payload_0_11952 = (_zz_dataOut_payload_0_11664 < _zz_dataOut_payload_0_11759);
  assign _zz_dataOut_payload_0_11953 = (_zz_dataOut_payload_0_11952 ? _zz_dataOut_payload_0_11664 : _zz_dataOut_payload_0_11759);
  assign _zz_dataOut_payload_0_11954 = (_zz_dataOut_payload_0_11952 ? _zz_dataOut_payload_0_11759 : _zz_dataOut_payload_0_11664);
  assign _zz_dataOut_payload_0_11955 = (_zz_dataOut_payload_0_11665 < _zz_dataOut_payload_0_11758);
  assign _zz_dataOut_payload_0_11956 = (_zz_dataOut_payload_0_11955 ? _zz_dataOut_payload_0_11665 : _zz_dataOut_payload_0_11758);
  assign _zz_dataOut_payload_0_11957 = (_zz_dataOut_payload_0_11955 ? _zz_dataOut_payload_0_11758 : _zz_dataOut_payload_0_11665);
  assign _zz_dataOut_payload_0_11958 = (_zz_dataOut_payload_0_11666 < _zz_dataOut_payload_0_11757);
  assign _zz_dataOut_payload_0_11959 = (_zz_dataOut_payload_0_11958 ? _zz_dataOut_payload_0_11666 : _zz_dataOut_payload_0_11757);
  assign _zz_dataOut_payload_0_11960 = (_zz_dataOut_payload_0_11958 ? _zz_dataOut_payload_0_11757 : _zz_dataOut_payload_0_11666);
  assign _zz_dataOut_payload_0_11961 = (_zz_dataOut_payload_0_11667 < _zz_dataOut_payload_0_11756);
  assign _zz_dataOut_payload_0_11962 = (_zz_dataOut_payload_0_11961 ? _zz_dataOut_payload_0_11667 : _zz_dataOut_payload_0_11756);
  assign _zz_dataOut_payload_0_11963 = (_zz_dataOut_payload_0_11961 ? _zz_dataOut_payload_0_11756 : _zz_dataOut_payload_0_11667);
  assign _zz_dataOut_payload_0_11964 = (_zz_dataOut_payload_0_11668 < _zz_dataOut_payload_0_11755);
  assign _zz_dataOut_payload_0_11965 = (_zz_dataOut_payload_0_11964 ? _zz_dataOut_payload_0_11668 : _zz_dataOut_payload_0_11755);
  assign _zz_dataOut_payload_0_11966 = (_zz_dataOut_payload_0_11964 ? _zz_dataOut_payload_0_11755 : _zz_dataOut_payload_0_11668);
  assign _zz_dataOut_payload_0_11967 = (_zz_dataOut_payload_0_11669 < _zz_dataOut_payload_0_11754);
  assign _zz_dataOut_payload_0_11968 = (_zz_dataOut_payload_0_11967 ? _zz_dataOut_payload_0_11669 : _zz_dataOut_payload_0_11754);
  assign _zz_dataOut_payload_0_11969 = (_zz_dataOut_payload_0_11967 ? _zz_dataOut_payload_0_11754 : _zz_dataOut_payload_0_11669);
  assign _zz_dataOut_payload_0_11970 = (_zz_dataOut_payload_0_11670 < _zz_dataOut_payload_0_11753);
  assign _zz_dataOut_payload_0_11971 = (_zz_dataOut_payload_0_11970 ? _zz_dataOut_payload_0_11670 : _zz_dataOut_payload_0_11753);
  assign _zz_dataOut_payload_0_11972 = (_zz_dataOut_payload_0_11970 ? _zz_dataOut_payload_0_11753 : _zz_dataOut_payload_0_11670);
  assign _zz_dataOut_payload_0_11973 = (_zz_dataOut_payload_0_11671 < _zz_dataOut_payload_0_11752);
  assign _zz_dataOut_payload_0_11974 = (_zz_dataOut_payload_0_11973 ? _zz_dataOut_payload_0_11671 : _zz_dataOut_payload_0_11752);
  assign _zz_dataOut_payload_0_11975 = (_zz_dataOut_payload_0_11973 ? _zz_dataOut_payload_0_11752 : _zz_dataOut_payload_0_11671);
  assign _zz_dataOut_payload_0_11976 = (_zz_dataOut_payload_0_11672 < _zz_dataOut_payload_0_11751);
  assign _zz_dataOut_payload_0_11977 = (_zz_dataOut_payload_0_11976 ? _zz_dataOut_payload_0_11672 : _zz_dataOut_payload_0_11751);
  assign _zz_dataOut_payload_0_11978 = (_zz_dataOut_payload_0_11976 ? _zz_dataOut_payload_0_11751 : _zz_dataOut_payload_0_11672);
  assign _zz_dataOut_payload_0_11979 = (_zz_dataOut_payload_0_11673 < _zz_dataOut_payload_0_11750);
  assign _zz_dataOut_payload_0_11980 = (_zz_dataOut_payload_0_11979 ? _zz_dataOut_payload_0_11673 : _zz_dataOut_payload_0_11750);
  assign _zz_dataOut_payload_0_11981 = (_zz_dataOut_payload_0_11979 ? _zz_dataOut_payload_0_11750 : _zz_dataOut_payload_0_11673);
  assign _zz_dataOut_payload_0_11982 = (_zz_dataOut_payload_0_11674 < _zz_dataOut_payload_0_11749);
  assign _zz_dataOut_payload_0_11983 = (_zz_dataOut_payload_0_11982 ? _zz_dataOut_payload_0_11674 : _zz_dataOut_payload_0_11749);
  assign _zz_dataOut_payload_0_11984 = (_zz_dataOut_payload_0_11982 ? _zz_dataOut_payload_0_11749 : _zz_dataOut_payload_0_11674);
  assign _zz_dataOut_payload_0_11985 = (_zz_dataOut_payload_0_11675 < _zz_dataOut_payload_0_11748);
  assign _zz_dataOut_payload_0_11986 = (_zz_dataOut_payload_0_11985 ? _zz_dataOut_payload_0_11675 : _zz_dataOut_payload_0_11748);
  assign _zz_dataOut_payload_0_11987 = (_zz_dataOut_payload_0_11985 ? _zz_dataOut_payload_0_11748 : _zz_dataOut_payload_0_11675);
  assign _zz_dataOut_payload_0_11988 = (_zz_dataOut_payload_0_11676 < _zz_dataOut_payload_0_11747);
  assign _zz_dataOut_payload_0_11989 = (_zz_dataOut_payload_0_11988 ? _zz_dataOut_payload_0_11676 : _zz_dataOut_payload_0_11747);
  assign _zz_dataOut_payload_0_11990 = (_zz_dataOut_payload_0_11988 ? _zz_dataOut_payload_0_11747 : _zz_dataOut_payload_0_11676);
  assign _zz_dataOut_payload_0_11991 = (_zz_dataOut_payload_0_11677 < _zz_dataOut_payload_0_11746);
  assign _zz_dataOut_payload_0_11992 = (_zz_dataOut_payload_0_11991 ? _zz_dataOut_payload_0_11677 : _zz_dataOut_payload_0_11746);
  assign _zz_dataOut_payload_0_11993 = (_zz_dataOut_payload_0_11991 ? _zz_dataOut_payload_0_11746 : _zz_dataOut_payload_0_11677);
  assign _zz_dataOut_payload_0_11994 = (_zz_dataOut_payload_0_11678 < _zz_dataOut_payload_0_11745);
  assign _zz_dataOut_payload_0_11995 = (_zz_dataOut_payload_0_11994 ? _zz_dataOut_payload_0_11678 : _zz_dataOut_payload_0_11745);
  assign _zz_dataOut_payload_0_11996 = (_zz_dataOut_payload_0_11994 ? _zz_dataOut_payload_0_11745 : _zz_dataOut_payload_0_11678);
  assign _zz_dataOut_payload_0_11997 = (_zz_dataOut_payload_0_11679 < _zz_dataOut_payload_0_11744);
  assign _zz_dataOut_payload_0_11998 = (_zz_dataOut_payload_0_11997 ? _zz_dataOut_payload_0_11679 : _zz_dataOut_payload_0_11744);
  assign _zz_dataOut_payload_0_11999 = (_zz_dataOut_payload_0_11997 ? _zz_dataOut_payload_0_11744 : _zz_dataOut_payload_0_11679);
  assign _zz_dataOut_payload_0_12000 = (_zz_dataOut_payload_0_11680 < _zz_dataOut_payload_0_11743);
  assign _zz_dataOut_payload_0_12001 = (_zz_dataOut_payload_0_12000 ? _zz_dataOut_payload_0_11680 : _zz_dataOut_payload_0_11743);
  assign _zz_dataOut_payload_0_12002 = (_zz_dataOut_payload_0_12000 ? _zz_dataOut_payload_0_11743 : _zz_dataOut_payload_0_11680);
  assign _zz_dataOut_payload_0_12003 = (_zz_dataOut_payload_0_11681 < _zz_dataOut_payload_0_11742);
  assign _zz_dataOut_payload_0_12004 = (_zz_dataOut_payload_0_12003 ? _zz_dataOut_payload_0_11681 : _zz_dataOut_payload_0_11742);
  assign _zz_dataOut_payload_0_12005 = (_zz_dataOut_payload_0_12003 ? _zz_dataOut_payload_0_11742 : _zz_dataOut_payload_0_11681);
  assign _zz_dataOut_payload_0_12006 = (_zz_dataOut_payload_0_11682 < _zz_dataOut_payload_0_11741);
  assign _zz_dataOut_payload_0_12007 = (_zz_dataOut_payload_0_12006 ? _zz_dataOut_payload_0_11682 : _zz_dataOut_payload_0_11741);
  assign _zz_dataOut_payload_0_12008 = (_zz_dataOut_payload_0_12006 ? _zz_dataOut_payload_0_11741 : _zz_dataOut_payload_0_11682);
  assign _zz_dataOut_payload_0_12009 = (_zz_dataOut_payload_0_11683 < _zz_dataOut_payload_0_11740);
  assign _zz_dataOut_payload_0_12010 = (_zz_dataOut_payload_0_12009 ? _zz_dataOut_payload_0_11683 : _zz_dataOut_payload_0_11740);
  assign _zz_dataOut_payload_0_12011 = (_zz_dataOut_payload_0_12009 ? _zz_dataOut_payload_0_11740 : _zz_dataOut_payload_0_11683);
  assign _zz_dataOut_payload_0_12012 = (_zz_dataOut_payload_0_11684 < _zz_dataOut_payload_0_11739);
  assign _zz_dataOut_payload_0_12013 = (_zz_dataOut_payload_0_12012 ? _zz_dataOut_payload_0_11684 : _zz_dataOut_payload_0_11739);
  assign _zz_dataOut_payload_0_12014 = (_zz_dataOut_payload_0_12012 ? _zz_dataOut_payload_0_11739 : _zz_dataOut_payload_0_11684);
  assign _zz_dataOut_payload_0_12015 = (_zz_dataOut_payload_0_11685 < _zz_dataOut_payload_0_11738);
  assign _zz_dataOut_payload_0_12016 = (_zz_dataOut_payload_0_12015 ? _zz_dataOut_payload_0_11685 : _zz_dataOut_payload_0_11738);
  assign _zz_dataOut_payload_0_12017 = (_zz_dataOut_payload_0_12015 ? _zz_dataOut_payload_0_11738 : _zz_dataOut_payload_0_11685);
  assign _zz_dataOut_payload_0_12018 = (_zz_dataOut_payload_0_11686 < _zz_dataOut_payload_0_11737);
  assign _zz_dataOut_payload_0_12019 = (_zz_dataOut_payload_0_12018 ? _zz_dataOut_payload_0_11686 : _zz_dataOut_payload_0_11737);
  assign _zz_dataOut_payload_0_12020 = (_zz_dataOut_payload_0_12018 ? _zz_dataOut_payload_0_11737 : _zz_dataOut_payload_0_11686);
  assign _zz_dataOut_payload_0_12021 = (_zz_dataOut_payload_0_11687 < _zz_dataOut_payload_0_11736);
  assign _zz_dataOut_payload_0_12022 = (_zz_dataOut_payload_0_12021 ? _zz_dataOut_payload_0_11687 : _zz_dataOut_payload_0_11736);
  assign _zz_dataOut_payload_0_12023 = (_zz_dataOut_payload_0_12021 ? _zz_dataOut_payload_0_11736 : _zz_dataOut_payload_0_11687);
  assign _zz_dataOut_payload_0_12024 = (_zz_dataOut_payload_0_11688 < _zz_dataOut_payload_0_11735);
  assign _zz_dataOut_payload_0_12025 = (_zz_dataOut_payload_0_12024 ? _zz_dataOut_payload_0_11688 : _zz_dataOut_payload_0_11735);
  assign _zz_dataOut_payload_0_12026 = (_zz_dataOut_payload_0_12024 ? _zz_dataOut_payload_0_11735 : _zz_dataOut_payload_0_11688);
  assign _zz_dataOut_payload_0_12027 = (_zz_dataOut_payload_0_11689 < _zz_dataOut_payload_0_11734);
  assign _zz_dataOut_payload_0_12028 = (_zz_dataOut_payload_0_12027 ? _zz_dataOut_payload_0_11689 : _zz_dataOut_payload_0_11734);
  assign _zz_dataOut_payload_0_12029 = (_zz_dataOut_payload_0_12027 ? _zz_dataOut_payload_0_11734 : _zz_dataOut_payload_0_11689);
  assign _zz_dataOut_payload_0_12030 = (_zz_dataOut_payload_0_11690 < _zz_dataOut_payload_0_11733);
  assign _zz_dataOut_payload_0_12031 = (_zz_dataOut_payload_0_12030 ? _zz_dataOut_payload_0_11690 : _zz_dataOut_payload_0_11733);
  assign _zz_dataOut_payload_0_12032 = (_zz_dataOut_payload_0_12030 ? _zz_dataOut_payload_0_11733 : _zz_dataOut_payload_0_11690);
  assign _zz_dataOut_payload_0_12033 = (_zz_dataOut_payload_0_11691 < _zz_dataOut_payload_0_11732);
  assign _zz_dataOut_payload_0_12034 = (_zz_dataOut_payload_0_12033 ? _zz_dataOut_payload_0_11691 : _zz_dataOut_payload_0_11732);
  assign _zz_dataOut_payload_0_12035 = (_zz_dataOut_payload_0_12033 ? _zz_dataOut_payload_0_11732 : _zz_dataOut_payload_0_11691);
  assign _zz_dataOut_payload_0_12036 = (_zz_dataOut_payload_0_11692 < _zz_dataOut_payload_0_11731);
  assign _zz_dataOut_payload_0_12037 = (_zz_dataOut_payload_0_12036 ? _zz_dataOut_payload_0_11692 : _zz_dataOut_payload_0_11731);
  assign _zz_dataOut_payload_0_12038 = (_zz_dataOut_payload_0_12036 ? _zz_dataOut_payload_0_11731 : _zz_dataOut_payload_0_11692);
  assign _zz_dataOut_payload_0_12039 = (_zz_dataOut_payload_0_11693 < _zz_dataOut_payload_0_11730);
  assign _zz_dataOut_payload_0_12040 = (_zz_dataOut_payload_0_12039 ? _zz_dataOut_payload_0_11693 : _zz_dataOut_payload_0_11730);
  assign _zz_dataOut_payload_0_12041 = (_zz_dataOut_payload_0_12039 ? _zz_dataOut_payload_0_11730 : _zz_dataOut_payload_0_11693);
  assign _zz_dataOut_payload_0_12042 = (_zz_dataOut_payload_0_11694 < _zz_dataOut_payload_0_11729);
  assign _zz_dataOut_payload_0_12043 = (_zz_dataOut_payload_0_12042 ? _zz_dataOut_payload_0_11694 : _zz_dataOut_payload_0_11729);
  assign _zz_dataOut_payload_0_12044 = (_zz_dataOut_payload_0_12042 ? _zz_dataOut_payload_0_11729 : _zz_dataOut_payload_0_11694);
  assign _zz_dataOut_payload_0_12045 = (_zz_dataOut_payload_0_11695 < _zz_dataOut_payload_0_11728);
  assign _zz_dataOut_payload_0_12046 = (_zz_dataOut_payload_0_12045 ? _zz_dataOut_payload_0_11695 : _zz_dataOut_payload_0_11728);
  assign _zz_dataOut_payload_0_12047 = (_zz_dataOut_payload_0_12045 ? _zz_dataOut_payload_0_11728 : _zz_dataOut_payload_0_11695);
  assign _zz_dataOut_payload_0_12048 = (_zz_dataOut_payload_0_11696 < _zz_dataOut_payload_0_11727);
  assign _zz_dataOut_payload_0_12049 = (_zz_dataOut_payload_0_12048 ? _zz_dataOut_payload_0_11696 : _zz_dataOut_payload_0_11727);
  assign _zz_dataOut_payload_0_12050 = (_zz_dataOut_payload_0_12048 ? _zz_dataOut_payload_0_11727 : _zz_dataOut_payload_0_11696);
  assign _zz_dataOut_payload_0_12051 = (_zz_dataOut_payload_0_11697 < _zz_dataOut_payload_0_11726);
  assign _zz_dataOut_payload_0_12052 = (_zz_dataOut_payload_0_12051 ? _zz_dataOut_payload_0_11697 : _zz_dataOut_payload_0_11726);
  assign _zz_dataOut_payload_0_12053 = (_zz_dataOut_payload_0_12051 ? _zz_dataOut_payload_0_11726 : _zz_dataOut_payload_0_11697);
  assign _zz_dataOut_payload_0_12054 = (_zz_dataOut_payload_0_11698 < _zz_dataOut_payload_0_11725);
  assign _zz_dataOut_payload_0_12055 = (_zz_dataOut_payload_0_12054 ? _zz_dataOut_payload_0_11698 : _zz_dataOut_payload_0_11725);
  assign _zz_dataOut_payload_0_12056 = (_zz_dataOut_payload_0_12054 ? _zz_dataOut_payload_0_11725 : _zz_dataOut_payload_0_11698);
  assign _zz_dataOut_payload_0_12057 = (_zz_dataOut_payload_0_11699 < _zz_dataOut_payload_0_11724);
  assign _zz_dataOut_payload_0_12058 = (_zz_dataOut_payload_0_12057 ? _zz_dataOut_payload_0_11699 : _zz_dataOut_payload_0_11724);
  assign _zz_dataOut_payload_0_12059 = (_zz_dataOut_payload_0_12057 ? _zz_dataOut_payload_0_11724 : _zz_dataOut_payload_0_11699);
  assign _zz_dataOut_payload_0_12060 = (_zz_dataOut_payload_0_11700 < _zz_dataOut_payload_0_11723);
  assign _zz_dataOut_payload_0_12061 = (_zz_dataOut_payload_0_12060 ? _zz_dataOut_payload_0_11700 : _zz_dataOut_payload_0_11723);
  assign _zz_dataOut_payload_0_12062 = (_zz_dataOut_payload_0_12060 ? _zz_dataOut_payload_0_11723 : _zz_dataOut_payload_0_11700);
  assign _zz_dataOut_payload_0_12063 = (_zz_dataOut_payload_0_11701 < _zz_dataOut_payload_0_11722);
  assign _zz_dataOut_payload_0_12064 = (_zz_dataOut_payload_0_12063 ? _zz_dataOut_payload_0_11701 : _zz_dataOut_payload_0_11722);
  assign _zz_dataOut_payload_0_12065 = (_zz_dataOut_payload_0_12063 ? _zz_dataOut_payload_0_11722 : _zz_dataOut_payload_0_11701);
  assign _zz_dataOut_payload_0_12066 = (_zz_dataOut_payload_0_11702 < _zz_dataOut_payload_0_11721);
  assign _zz_dataOut_payload_0_12067 = (_zz_dataOut_payload_0_12066 ? _zz_dataOut_payload_0_11702 : _zz_dataOut_payload_0_11721);
  assign _zz_dataOut_payload_0_12068 = (_zz_dataOut_payload_0_12066 ? _zz_dataOut_payload_0_11721 : _zz_dataOut_payload_0_11702);
  assign _zz_dataOut_payload_0_12069 = (_zz_dataOut_payload_0_11703 < _zz_dataOut_payload_0_11720);
  assign _zz_dataOut_payload_0_12070 = (_zz_dataOut_payload_0_12069 ? _zz_dataOut_payload_0_11703 : _zz_dataOut_payload_0_11720);
  assign _zz_dataOut_payload_0_12071 = (_zz_dataOut_payload_0_12069 ? _zz_dataOut_payload_0_11720 : _zz_dataOut_payload_0_11703);
  assign _zz_dataOut_payload_0_12072 = (_zz_dataOut_payload_0_11704 < _zz_dataOut_payload_0_11719);
  assign _zz_dataOut_payload_0_12073 = (_zz_dataOut_payload_0_12072 ? _zz_dataOut_payload_0_11704 : _zz_dataOut_payload_0_11719);
  assign _zz_dataOut_payload_0_12074 = (_zz_dataOut_payload_0_12072 ? _zz_dataOut_payload_0_11719 : _zz_dataOut_payload_0_11704);
  assign _zz_dataOut_payload_0_12075 = (_zz_dataOut_payload_0_11705 < _zz_dataOut_payload_0_11718);
  assign _zz_dataOut_payload_0_12076 = (_zz_dataOut_payload_0_12075 ? _zz_dataOut_payload_0_11705 : _zz_dataOut_payload_0_11718);
  assign _zz_dataOut_payload_0_12077 = (_zz_dataOut_payload_0_12075 ? _zz_dataOut_payload_0_11718 : _zz_dataOut_payload_0_11705);
  assign _zz_dataOut_payload_0_12078 = (_zz_dataOut_payload_0_11706 < _zz_dataOut_payload_0_11717);
  assign _zz_dataOut_payload_0_12079 = (_zz_dataOut_payload_0_12078 ? _zz_dataOut_payload_0_11706 : _zz_dataOut_payload_0_11717);
  assign _zz_dataOut_payload_0_12080 = (_zz_dataOut_payload_0_12078 ? _zz_dataOut_payload_0_11717 : _zz_dataOut_payload_0_11706);
  assign _zz_dataOut_payload_0_12081 = (_zz_dataOut_payload_0_11707 < _zz_dataOut_payload_0_11716);
  assign _zz_dataOut_payload_0_12082 = (_zz_dataOut_payload_0_12081 ? _zz_dataOut_payload_0_11707 : _zz_dataOut_payload_0_11716);
  assign _zz_dataOut_payload_0_12083 = (_zz_dataOut_payload_0_12081 ? _zz_dataOut_payload_0_11716 : _zz_dataOut_payload_0_11707);
  assign _zz_dataOut_payload_0_12084 = (_zz_dataOut_payload_0_11708 < _zz_dataOut_payload_0_11715);
  assign _zz_dataOut_payload_0_12085 = (_zz_dataOut_payload_0_12084 ? _zz_dataOut_payload_0_11708 : _zz_dataOut_payload_0_11715);
  assign _zz_dataOut_payload_0_12086 = (_zz_dataOut_payload_0_12084 ? _zz_dataOut_payload_0_11715 : _zz_dataOut_payload_0_11708);
  assign _zz_dataOut_payload_0_12087 = (_zz_dataOut_payload_0_11709 < _zz_dataOut_payload_0_11714);
  assign _zz_dataOut_payload_0_12088 = (_zz_dataOut_payload_0_12087 ? _zz_dataOut_payload_0_11709 : _zz_dataOut_payload_0_11714);
  assign _zz_dataOut_payload_0_12089 = (_zz_dataOut_payload_0_12087 ? _zz_dataOut_payload_0_11714 : _zz_dataOut_payload_0_11709);
  assign _zz_dataOut_payload_0_12090 = (_zz_dataOut_payload_0_11710 < _zz_dataOut_payload_0_11713);
  assign _zz_dataOut_payload_0_12091 = (_zz_dataOut_payload_0_12090 ? _zz_dataOut_payload_0_11710 : _zz_dataOut_payload_0_11713);
  assign _zz_dataOut_payload_0_12092 = (_zz_dataOut_payload_0_12090 ? _zz_dataOut_payload_0_11713 : _zz_dataOut_payload_0_11710);
  assign _zz_dataOut_payload_0_12093 = (_zz_dataOut_payload_0_11711 < _zz_dataOut_payload_0_11712);
  assign _zz_dataOut_payload_0_12094 = (_zz_dataOut_payload_0_12093 ? _zz_dataOut_payload_0_11711 : _zz_dataOut_payload_0_11712);
  assign _zz_dataOut_payload_0_12095 = (_zz_dataOut_payload_0_12093 ? _zz_dataOut_payload_0_11712 : _zz_dataOut_payload_0_11711);
  assign _zz_dataOut_payload_0_12096 = (_zz_dataOut_payload_0_11905 < _zz_dataOut_payload_0_12001);
  assign _zz_dataOut_payload_0_12097 = (_zz_dataOut_payload_0_12096 ? _zz_dataOut_payload_0_11905 : _zz_dataOut_payload_0_12001);
  assign _zz_dataOut_payload_0_12098 = (_zz_dataOut_payload_0_12096 ? _zz_dataOut_payload_0_12001 : _zz_dataOut_payload_0_11905);
  assign _zz_dataOut_payload_0_12099 = (_zz_dataOut_payload_0_11908 < _zz_dataOut_payload_0_12004);
  assign _zz_dataOut_payload_0_12100 = (_zz_dataOut_payload_0_12099 ? _zz_dataOut_payload_0_11908 : _zz_dataOut_payload_0_12004);
  assign _zz_dataOut_payload_0_12101 = (_zz_dataOut_payload_0_12099 ? _zz_dataOut_payload_0_12004 : _zz_dataOut_payload_0_11908);
  assign _zz_dataOut_payload_0_12102 = (_zz_dataOut_payload_0_11911 < _zz_dataOut_payload_0_12007);
  assign _zz_dataOut_payload_0_12103 = (_zz_dataOut_payload_0_12102 ? _zz_dataOut_payload_0_11911 : _zz_dataOut_payload_0_12007);
  assign _zz_dataOut_payload_0_12104 = (_zz_dataOut_payload_0_12102 ? _zz_dataOut_payload_0_12007 : _zz_dataOut_payload_0_11911);
  assign _zz_dataOut_payload_0_12105 = (_zz_dataOut_payload_0_11914 < _zz_dataOut_payload_0_12010);
  assign _zz_dataOut_payload_0_12106 = (_zz_dataOut_payload_0_12105 ? _zz_dataOut_payload_0_11914 : _zz_dataOut_payload_0_12010);
  assign _zz_dataOut_payload_0_12107 = (_zz_dataOut_payload_0_12105 ? _zz_dataOut_payload_0_12010 : _zz_dataOut_payload_0_11914);
  assign _zz_dataOut_payload_0_12108 = (_zz_dataOut_payload_0_11917 < _zz_dataOut_payload_0_12013);
  assign _zz_dataOut_payload_0_12109 = (_zz_dataOut_payload_0_12108 ? _zz_dataOut_payload_0_11917 : _zz_dataOut_payload_0_12013);
  assign _zz_dataOut_payload_0_12110 = (_zz_dataOut_payload_0_12108 ? _zz_dataOut_payload_0_12013 : _zz_dataOut_payload_0_11917);
  assign _zz_dataOut_payload_0_12111 = (_zz_dataOut_payload_0_11920 < _zz_dataOut_payload_0_12016);
  assign _zz_dataOut_payload_0_12112 = (_zz_dataOut_payload_0_12111 ? _zz_dataOut_payload_0_11920 : _zz_dataOut_payload_0_12016);
  assign _zz_dataOut_payload_0_12113 = (_zz_dataOut_payload_0_12111 ? _zz_dataOut_payload_0_12016 : _zz_dataOut_payload_0_11920);
  assign _zz_dataOut_payload_0_12114 = (_zz_dataOut_payload_0_11923 < _zz_dataOut_payload_0_12019);
  assign _zz_dataOut_payload_0_12115 = (_zz_dataOut_payload_0_12114 ? _zz_dataOut_payload_0_11923 : _zz_dataOut_payload_0_12019);
  assign _zz_dataOut_payload_0_12116 = (_zz_dataOut_payload_0_12114 ? _zz_dataOut_payload_0_12019 : _zz_dataOut_payload_0_11923);
  assign _zz_dataOut_payload_0_12117 = (_zz_dataOut_payload_0_11926 < _zz_dataOut_payload_0_12022);
  assign _zz_dataOut_payload_0_12118 = (_zz_dataOut_payload_0_12117 ? _zz_dataOut_payload_0_11926 : _zz_dataOut_payload_0_12022);
  assign _zz_dataOut_payload_0_12119 = (_zz_dataOut_payload_0_12117 ? _zz_dataOut_payload_0_12022 : _zz_dataOut_payload_0_11926);
  assign _zz_dataOut_payload_0_12120 = (_zz_dataOut_payload_0_11929 < _zz_dataOut_payload_0_12025);
  assign _zz_dataOut_payload_0_12121 = (_zz_dataOut_payload_0_12120 ? _zz_dataOut_payload_0_11929 : _zz_dataOut_payload_0_12025);
  assign _zz_dataOut_payload_0_12122 = (_zz_dataOut_payload_0_12120 ? _zz_dataOut_payload_0_12025 : _zz_dataOut_payload_0_11929);
  assign _zz_dataOut_payload_0_12123 = (_zz_dataOut_payload_0_11932 < _zz_dataOut_payload_0_12028);
  assign _zz_dataOut_payload_0_12124 = (_zz_dataOut_payload_0_12123 ? _zz_dataOut_payload_0_11932 : _zz_dataOut_payload_0_12028);
  assign _zz_dataOut_payload_0_12125 = (_zz_dataOut_payload_0_12123 ? _zz_dataOut_payload_0_12028 : _zz_dataOut_payload_0_11932);
  assign _zz_dataOut_payload_0_12126 = (_zz_dataOut_payload_0_11935 < _zz_dataOut_payload_0_12031);
  assign _zz_dataOut_payload_0_12127 = (_zz_dataOut_payload_0_12126 ? _zz_dataOut_payload_0_11935 : _zz_dataOut_payload_0_12031);
  assign _zz_dataOut_payload_0_12128 = (_zz_dataOut_payload_0_12126 ? _zz_dataOut_payload_0_12031 : _zz_dataOut_payload_0_11935);
  assign _zz_dataOut_payload_0_12129 = (_zz_dataOut_payload_0_11938 < _zz_dataOut_payload_0_12034);
  assign _zz_dataOut_payload_0_12130 = (_zz_dataOut_payload_0_12129 ? _zz_dataOut_payload_0_11938 : _zz_dataOut_payload_0_12034);
  assign _zz_dataOut_payload_0_12131 = (_zz_dataOut_payload_0_12129 ? _zz_dataOut_payload_0_12034 : _zz_dataOut_payload_0_11938);
  assign _zz_dataOut_payload_0_12132 = (_zz_dataOut_payload_0_11941 < _zz_dataOut_payload_0_12037);
  assign _zz_dataOut_payload_0_12133 = (_zz_dataOut_payload_0_12132 ? _zz_dataOut_payload_0_11941 : _zz_dataOut_payload_0_12037);
  assign _zz_dataOut_payload_0_12134 = (_zz_dataOut_payload_0_12132 ? _zz_dataOut_payload_0_12037 : _zz_dataOut_payload_0_11941);
  assign _zz_dataOut_payload_0_12135 = (_zz_dataOut_payload_0_11944 < _zz_dataOut_payload_0_12040);
  assign _zz_dataOut_payload_0_12136 = (_zz_dataOut_payload_0_12135 ? _zz_dataOut_payload_0_11944 : _zz_dataOut_payload_0_12040);
  assign _zz_dataOut_payload_0_12137 = (_zz_dataOut_payload_0_12135 ? _zz_dataOut_payload_0_12040 : _zz_dataOut_payload_0_11944);
  assign _zz_dataOut_payload_0_12138 = (_zz_dataOut_payload_0_11947 < _zz_dataOut_payload_0_12043);
  assign _zz_dataOut_payload_0_12139 = (_zz_dataOut_payload_0_12138 ? _zz_dataOut_payload_0_11947 : _zz_dataOut_payload_0_12043);
  assign _zz_dataOut_payload_0_12140 = (_zz_dataOut_payload_0_12138 ? _zz_dataOut_payload_0_12043 : _zz_dataOut_payload_0_11947);
  assign _zz_dataOut_payload_0_12141 = (_zz_dataOut_payload_0_11950 < _zz_dataOut_payload_0_12046);
  assign _zz_dataOut_payload_0_12142 = (_zz_dataOut_payload_0_12141 ? _zz_dataOut_payload_0_11950 : _zz_dataOut_payload_0_12046);
  assign _zz_dataOut_payload_0_12143 = (_zz_dataOut_payload_0_12141 ? _zz_dataOut_payload_0_12046 : _zz_dataOut_payload_0_11950);
  assign _zz_dataOut_payload_0_12144 = (_zz_dataOut_payload_0_11953 < _zz_dataOut_payload_0_12049);
  assign _zz_dataOut_payload_0_12145 = (_zz_dataOut_payload_0_12144 ? _zz_dataOut_payload_0_11953 : _zz_dataOut_payload_0_12049);
  assign _zz_dataOut_payload_0_12146 = (_zz_dataOut_payload_0_12144 ? _zz_dataOut_payload_0_12049 : _zz_dataOut_payload_0_11953);
  assign _zz_dataOut_payload_0_12147 = (_zz_dataOut_payload_0_11956 < _zz_dataOut_payload_0_12052);
  assign _zz_dataOut_payload_0_12148 = (_zz_dataOut_payload_0_12147 ? _zz_dataOut_payload_0_11956 : _zz_dataOut_payload_0_12052);
  assign _zz_dataOut_payload_0_12149 = (_zz_dataOut_payload_0_12147 ? _zz_dataOut_payload_0_12052 : _zz_dataOut_payload_0_11956);
  assign _zz_dataOut_payload_0_12150 = (_zz_dataOut_payload_0_11959 < _zz_dataOut_payload_0_12055);
  assign _zz_dataOut_payload_0_12151 = (_zz_dataOut_payload_0_12150 ? _zz_dataOut_payload_0_11959 : _zz_dataOut_payload_0_12055);
  assign _zz_dataOut_payload_0_12152 = (_zz_dataOut_payload_0_12150 ? _zz_dataOut_payload_0_12055 : _zz_dataOut_payload_0_11959);
  assign _zz_dataOut_payload_0_12153 = (_zz_dataOut_payload_0_11962 < _zz_dataOut_payload_0_12058);
  assign _zz_dataOut_payload_0_12154 = (_zz_dataOut_payload_0_12153 ? _zz_dataOut_payload_0_11962 : _zz_dataOut_payload_0_12058);
  assign _zz_dataOut_payload_0_12155 = (_zz_dataOut_payload_0_12153 ? _zz_dataOut_payload_0_12058 : _zz_dataOut_payload_0_11962);
  assign _zz_dataOut_payload_0_12156 = (_zz_dataOut_payload_0_11965 < _zz_dataOut_payload_0_12061);
  assign _zz_dataOut_payload_0_12157 = (_zz_dataOut_payload_0_12156 ? _zz_dataOut_payload_0_11965 : _zz_dataOut_payload_0_12061);
  assign _zz_dataOut_payload_0_12158 = (_zz_dataOut_payload_0_12156 ? _zz_dataOut_payload_0_12061 : _zz_dataOut_payload_0_11965);
  assign _zz_dataOut_payload_0_12159 = (_zz_dataOut_payload_0_11968 < _zz_dataOut_payload_0_12064);
  assign _zz_dataOut_payload_0_12160 = (_zz_dataOut_payload_0_12159 ? _zz_dataOut_payload_0_11968 : _zz_dataOut_payload_0_12064);
  assign _zz_dataOut_payload_0_12161 = (_zz_dataOut_payload_0_12159 ? _zz_dataOut_payload_0_12064 : _zz_dataOut_payload_0_11968);
  assign _zz_dataOut_payload_0_12162 = (_zz_dataOut_payload_0_11971 < _zz_dataOut_payload_0_12067);
  assign _zz_dataOut_payload_0_12163 = (_zz_dataOut_payload_0_12162 ? _zz_dataOut_payload_0_11971 : _zz_dataOut_payload_0_12067);
  assign _zz_dataOut_payload_0_12164 = (_zz_dataOut_payload_0_12162 ? _zz_dataOut_payload_0_12067 : _zz_dataOut_payload_0_11971);
  assign _zz_dataOut_payload_0_12165 = (_zz_dataOut_payload_0_11974 < _zz_dataOut_payload_0_12070);
  assign _zz_dataOut_payload_0_12166 = (_zz_dataOut_payload_0_12165 ? _zz_dataOut_payload_0_11974 : _zz_dataOut_payload_0_12070);
  assign _zz_dataOut_payload_0_12167 = (_zz_dataOut_payload_0_12165 ? _zz_dataOut_payload_0_12070 : _zz_dataOut_payload_0_11974);
  assign _zz_dataOut_payload_0_12168 = (_zz_dataOut_payload_0_11977 < _zz_dataOut_payload_0_12073);
  assign _zz_dataOut_payload_0_12169 = (_zz_dataOut_payload_0_12168 ? _zz_dataOut_payload_0_11977 : _zz_dataOut_payload_0_12073);
  assign _zz_dataOut_payload_0_12170 = (_zz_dataOut_payload_0_12168 ? _zz_dataOut_payload_0_12073 : _zz_dataOut_payload_0_11977);
  assign _zz_dataOut_payload_0_12171 = (_zz_dataOut_payload_0_11980 < _zz_dataOut_payload_0_12076);
  assign _zz_dataOut_payload_0_12172 = (_zz_dataOut_payload_0_12171 ? _zz_dataOut_payload_0_11980 : _zz_dataOut_payload_0_12076);
  assign _zz_dataOut_payload_0_12173 = (_zz_dataOut_payload_0_12171 ? _zz_dataOut_payload_0_12076 : _zz_dataOut_payload_0_11980);
  assign _zz_dataOut_payload_0_12174 = (_zz_dataOut_payload_0_11983 < _zz_dataOut_payload_0_12079);
  assign _zz_dataOut_payload_0_12175 = (_zz_dataOut_payload_0_12174 ? _zz_dataOut_payload_0_11983 : _zz_dataOut_payload_0_12079);
  assign _zz_dataOut_payload_0_12176 = (_zz_dataOut_payload_0_12174 ? _zz_dataOut_payload_0_12079 : _zz_dataOut_payload_0_11983);
  assign _zz_dataOut_payload_0_12177 = (_zz_dataOut_payload_0_11986 < _zz_dataOut_payload_0_12082);
  assign _zz_dataOut_payload_0_12178 = (_zz_dataOut_payload_0_12177 ? _zz_dataOut_payload_0_11986 : _zz_dataOut_payload_0_12082);
  assign _zz_dataOut_payload_0_12179 = (_zz_dataOut_payload_0_12177 ? _zz_dataOut_payload_0_12082 : _zz_dataOut_payload_0_11986);
  assign _zz_dataOut_payload_0_12180 = (_zz_dataOut_payload_0_11989 < _zz_dataOut_payload_0_12085);
  assign _zz_dataOut_payload_0_12181 = (_zz_dataOut_payload_0_12180 ? _zz_dataOut_payload_0_11989 : _zz_dataOut_payload_0_12085);
  assign _zz_dataOut_payload_0_12182 = (_zz_dataOut_payload_0_12180 ? _zz_dataOut_payload_0_12085 : _zz_dataOut_payload_0_11989);
  assign _zz_dataOut_payload_0_12183 = (_zz_dataOut_payload_0_11992 < _zz_dataOut_payload_0_12088);
  assign _zz_dataOut_payload_0_12184 = (_zz_dataOut_payload_0_12183 ? _zz_dataOut_payload_0_11992 : _zz_dataOut_payload_0_12088);
  assign _zz_dataOut_payload_0_12185 = (_zz_dataOut_payload_0_12183 ? _zz_dataOut_payload_0_12088 : _zz_dataOut_payload_0_11992);
  assign _zz_dataOut_payload_0_12186 = (_zz_dataOut_payload_0_11995 < _zz_dataOut_payload_0_12091);
  assign _zz_dataOut_payload_0_12187 = (_zz_dataOut_payload_0_12186 ? _zz_dataOut_payload_0_11995 : _zz_dataOut_payload_0_12091);
  assign _zz_dataOut_payload_0_12188 = (_zz_dataOut_payload_0_12186 ? _zz_dataOut_payload_0_12091 : _zz_dataOut_payload_0_11995);
  assign _zz_dataOut_payload_0_12189 = (_zz_dataOut_payload_0_11998 < _zz_dataOut_payload_0_12094);
  assign _zz_dataOut_payload_0_12190 = (_zz_dataOut_payload_0_12189 ? _zz_dataOut_payload_0_11998 : _zz_dataOut_payload_0_12094);
  assign _zz_dataOut_payload_0_12191 = (_zz_dataOut_payload_0_12189 ? _zz_dataOut_payload_0_12094 : _zz_dataOut_payload_0_11998);
  assign _zz_dataOut_payload_0_12192 = (_zz_dataOut_payload_0_12097 < _zz_dataOut_payload_0_12145);
  assign _zz_dataOut_payload_0_12193 = (_zz_dataOut_payload_0_12192 ? _zz_dataOut_payload_0_12097 : _zz_dataOut_payload_0_12145);
  assign _zz_dataOut_payload_0_12194 = (_zz_dataOut_payload_0_12192 ? _zz_dataOut_payload_0_12145 : _zz_dataOut_payload_0_12097);
  assign _zz_dataOut_payload_0_12195 = (_zz_dataOut_payload_0_12100 < _zz_dataOut_payload_0_12148);
  assign _zz_dataOut_payload_0_12196 = (_zz_dataOut_payload_0_12195 ? _zz_dataOut_payload_0_12100 : _zz_dataOut_payload_0_12148);
  assign _zz_dataOut_payload_0_12197 = (_zz_dataOut_payload_0_12195 ? _zz_dataOut_payload_0_12148 : _zz_dataOut_payload_0_12100);
  assign _zz_dataOut_payload_0_12198 = (_zz_dataOut_payload_0_12103 < _zz_dataOut_payload_0_12151);
  assign _zz_dataOut_payload_0_12199 = (_zz_dataOut_payload_0_12198 ? _zz_dataOut_payload_0_12103 : _zz_dataOut_payload_0_12151);
  assign _zz_dataOut_payload_0_12200 = (_zz_dataOut_payload_0_12198 ? _zz_dataOut_payload_0_12151 : _zz_dataOut_payload_0_12103);
  assign _zz_dataOut_payload_0_12201 = (_zz_dataOut_payload_0_12106 < _zz_dataOut_payload_0_12154);
  assign _zz_dataOut_payload_0_12202 = (_zz_dataOut_payload_0_12201 ? _zz_dataOut_payload_0_12106 : _zz_dataOut_payload_0_12154);
  assign _zz_dataOut_payload_0_12203 = (_zz_dataOut_payload_0_12201 ? _zz_dataOut_payload_0_12154 : _zz_dataOut_payload_0_12106);
  assign _zz_dataOut_payload_0_12204 = (_zz_dataOut_payload_0_12109 < _zz_dataOut_payload_0_12157);
  assign _zz_dataOut_payload_0_12205 = (_zz_dataOut_payload_0_12204 ? _zz_dataOut_payload_0_12109 : _zz_dataOut_payload_0_12157);
  assign _zz_dataOut_payload_0_12206 = (_zz_dataOut_payload_0_12204 ? _zz_dataOut_payload_0_12157 : _zz_dataOut_payload_0_12109);
  assign _zz_dataOut_payload_0_12207 = (_zz_dataOut_payload_0_12112 < _zz_dataOut_payload_0_12160);
  assign _zz_dataOut_payload_0_12208 = (_zz_dataOut_payload_0_12207 ? _zz_dataOut_payload_0_12112 : _zz_dataOut_payload_0_12160);
  assign _zz_dataOut_payload_0_12209 = (_zz_dataOut_payload_0_12207 ? _zz_dataOut_payload_0_12160 : _zz_dataOut_payload_0_12112);
  assign _zz_dataOut_payload_0_12210 = (_zz_dataOut_payload_0_12115 < _zz_dataOut_payload_0_12163);
  assign _zz_dataOut_payload_0_12211 = (_zz_dataOut_payload_0_12210 ? _zz_dataOut_payload_0_12115 : _zz_dataOut_payload_0_12163);
  assign _zz_dataOut_payload_0_12212 = (_zz_dataOut_payload_0_12210 ? _zz_dataOut_payload_0_12163 : _zz_dataOut_payload_0_12115);
  assign _zz_dataOut_payload_0_12213 = (_zz_dataOut_payload_0_12118 < _zz_dataOut_payload_0_12166);
  assign _zz_dataOut_payload_0_12214 = (_zz_dataOut_payload_0_12213 ? _zz_dataOut_payload_0_12118 : _zz_dataOut_payload_0_12166);
  assign _zz_dataOut_payload_0_12215 = (_zz_dataOut_payload_0_12213 ? _zz_dataOut_payload_0_12166 : _zz_dataOut_payload_0_12118);
  assign _zz_dataOut_payload_0_12216 = (_zz_dataOut_payload_0_12121 < _zz_dataOut_payload_0_12169);
  assign _zz_dataOut_payload_0_12217 = (_zz_dataOut_payload_0_12216 ? _zz_dataOut_payload_0_12121 : _zz_dataOut_payload_0_12169);
  assign _zz_dataOut_payload_0_12218 = (_zz_dataOut_payload_0_12216 ? _zz_dataOut_payload_0_12169 : _zz_dataOut_payload_0_12121);
  assign _zz_dataOut_payload_0_12219 = (_zz_dataOut_payload_0_12124 < _zz_dataOut_payload_0_12172);
  assign _zz_dataOut_payload_0_12220 = (_zz_dataOut_payload_0_12219 ? _zz_dataOut_payload_0_12124 : _zz_dataOut_payload_0_12172);
  assign _zz_dataOut_payload_0_12221 = (_zz_dataOut_payload_0_12219 ? _zz_dataOut_payload_0_12172 : _zz_dataOut_payload_0_12124);
  assign _zz_dataOut_payload_0_12222 = (_zz_dataOut_payload_0_12127 < _zz_dataOut_payload_0_12175);
  assign _zz_dataOut_payload_0_12223 = (_zz_dataOut_payload_0_12222 ? _zz_dataOut_payload_0_12127 : _zz_dataOut_payload_0_12175);
  assign _zz_dataOut_payload_0_12224 = (_zz_dataOut_payload_0_12222 ? _zz_dataOut_payload_0_12175 : _zz_dataOut_payload_0_12127);
  assign _zz_dataOut_payload_0_12225 = (_zz_dataOut_payload_0_12130 < _zz_dataOut_payload_0_12178);
  assign _zz_dataOut_payload_0_12226 = (_zz_dataOut_payload_0_12225 ? _zz_dataOut_payload_0_12130 : _zz_dataOut_payload_0_12178);
  assign _zz_dataOut_payload_0_12227 = (_zz_dataOut_payload_0_12225 ? _zz_dataOut_payload_0_12178 : _zz_dataOut_payload_0_12130);
  assign _zz_dataOut_payload_0_12228 = (_zz_dataOut_payload_0_12133 < _zz_dataOut_payload_0_12181);
  assign _zz_dataOut_payload_0_12229 = (_zz_dataOut_payload_0_12228 ? _zz_dataOut_payload_0_12133 : _zz_dataOut_payload_0_12181);
  assign _zz_dataOut_payload_0_12230 = (_zz_dataOut_payload_0_12228 ? _zz_dataOut_payload_0_12181 : _zz_dataOut_payload_0_12133);
  assign _zz_dataOut_payload_0_12231 = (_zz_dataOut_payload_0_12136 < _zz_dataOut_payload_0_12184);
  assign _zz_dataOut_payload_0_12232 = (_zz_dataOut_payload_0_12231 ? _zz_dataOut_payload_0_12136 : _zz_dataOut_payload_0_12184);
  assign _zz_dataOut_payload_0_12233 = (_zz_dataOut_payload_0_12231 ? _zz_dataOut_payload_0_12184 : _zz_dataOut_payload_0_12136);
  assign _zz_dataOut_payload_0_12234 = (_zz_dataOut_payload_0_12139 < _zz_dataOut_payload_0_12187);
  assign _zz_dataOut_payload_0_12235 = (_zz_dataOut_payload_0_12234 ? _zz_dataOut_payload_0_12139 : _zz_dataOut_payload_0_12187);
  assign _zz_dataOut_payload_0_12236 = (_zz_dataOut_payload_0_12234 ? _zz_dataOut_payload_0_12187 : _zz_dataOut_payload_0_12139);
  assign _zz_dataOut_payload_0_12237 = (_zz_dataOut_payload_0_12142 < _zz_dataOut_payload_0_12190);
  assign _zz_dataOut_payload_0_12238 = (_zz_dataOut_payload_0_12237 ? _zz_dataOut_payload_0_12142 : _zz_dataOut_payload_0_12190);
  assign _zz_dataOut_payload_0_12239 = (_zz_dataOut_payload_0_12237 ? _zz_dataOut_payload_0_12190 : _zz_dataOut_payload_0_12142);
  assign _zz_dataOut_payload_0_12240 = (_zz_dataOut_payload_0_12193 < _zz_dataOut_payload_0_12217);
  assign _zz_dataOut_payload_0_12241 = (_zz_dataOut_payload_0_12240 ? _zz_dataOut_payload_0_12193 : _zz_dataOut_payload_0_12217);
  assign _zz_dataOut_payload_0_12242 = (_zz_dataOut_payload_0_12240 ? _zz_dataOut_payload_0_12217 : _zz_dataOut_payload_0_12193);
  assign _zz_dataOut_payload_0_12243 = (_zz_dataOut_payload_0_12196 < _zz_dataOut_payload_0_12220);
  assign _zz_dataOut_payload_0_12244 = (_zz_dataOut_payload_0_12243 ? _zz_dataOut_payload_0_12196 : _zz_dataOut_payload_0_12220);
  assign _zz_dataOut_payload_0_12245 = (_zz_dataOut_payload_0_12243 ? _zz_dataOut_payload_0_12220 : _zz_dataOut_payload_0_12196);
  assign _zz_dataOut_payload_0_12246 = (_zz_dataOut_payload_0_12199 < _zz_dataOut_payload_0_12223);
  assign _zz_dataOut_payload_0_12247 = (_zz_dataOut_payload_0_12246 ? _zz_dataOut_payload_0_12199 : _zz_dataOut_payload_0_12223);
  assign _zz_dataOut_payload_0_12248 = (_zz_dataOut_payload_0_12246 ? _zz_dataOut_payload_0_12223 : _zz_dataOut_payload_0_12199);
  assign _zz_dataOut_payload_0_12249 = (_zz_dataOut_payload_0_12202 < _zz_dataOut_payload_0_12226);
  assign _zz_dataOut_payload_0_12250 = (_zz_dataOut_payload_0_12249 ? _zz_dataOut_payload_0_12202 : _zz_dataOut_payload_0_12226);
  assign _zz_dataOut_payload_0_12251 = (_zz_dataOut_payload_0_12249 ? _zz_dataOut_payload_0_12226 : _zz_dataOut_payload_0_12202);
  assign _zz_dataOut_payload_0_12252 = (_zz_dataOut_payload_0_12205 < _zz_dataOut_payload_0_12229);
  assign _zz_dataOut_payload_0_12253 = (_zz_dataOut_payload_0_12252 ? _zz_dataOut_payload_0_12205 : _zz_dataOut_payload_0_12229);
  assign _zz_dataOut_payload_0_12254 = (_zz_dataOut_payload_0_12252 ? _zz_dataOut_payload_0_12229 : _zz_dataOut_payload_0_12205);
  assign _zz_dataOut_payload_0_12255 = (_zz_dataOut_payload_0_12208 < _zz_dataOut_payload_0_12232);
  assign _zz_dataOut_payload_0_12256 = (_zz_dataOut_payload_0_12255 ? _zz_dataOut_payload_0_12208 : _zz_dataOut_payload_0_12232);
  assign _zz_dataOut_payload_0_12257 = (_zz_dataOut_payload_0_12255 ? _zz_dataOut_payload_0_12232 : _zz_dataOut_payload_0_12208);
  assign _zz_dataOut_payload_0_12258 = (_zz_dataOut_payload_0_12211 < _zz_dataOut_payload_0_12235);
  assign _zz_dataOut_payload_0_12259 = (_zz_dataOut_payload_0_12258 ? _zz_dataOut_payload_0_12211 : _zz_dataOut_payload_0_12235);
  assign _zz_dataOut_payload_0_12260 = (_zz_dataOut_payload_0_12258 ? _zz_dataOut_payload_0_12235 : _zz_dataOut_payload_0_12211);
  assign _zz_dataOut_payload_0_12261 = (_zz_dataOut_payload_0_12214 < _zz_dataOut_payload_0_12238);
  assign _zz_dataOut_payload_0_12262 = (_zz_dataOut_payload_0_12261 ? _zz_dataOut_payload_0_12214 : _zz_dataOut_payload_0_12238);
  assign _zz_dataOut_payload_0_12263 = (_zz_dataOut_payload_0_12261 ? _zz_dataOut_payload_0_12238 : _zz_dataOut_payload_0_12214);
  assign _zz_dataOut_payload_0_12264 = (_zz_dataOut_payload_0_12241 < _zz_dataOut_payload_0_12253);
  assign _zz_dataOut_payload_0_12265 = (_zz_dataOut_payload_0_12264 ? _zz_dataOut_payload_0_12241 : _zz_dataOut_payload_0_12253);
  assign _zz_dataOut_payload_0_12266 = (_zz_dataOut_payload_0_12264 ? _zz_dataOut_payload_0_12253 : _zz_dataOut_payload_0_12241);
  assign _zz_dataOut_payload_0_12267 = (_zz_dataOut_payload_0_12244 < _zz_dataOut_payload_0_12256);
  assign _zz_dataOut_payload_0_12268 = (_zz_dataOut_payload_0_12267 ? _zz_dataOut_payload_0_12244 : _zz_dataOut_payload_0_12256);
  assign _zz_dataOut_payload_0_12269 = (_zz_dataOut_payload_0_12267 ? _zz_dataOut_payload_0_12256 : _zz_dataOut_payload_0_12244);
  assign _zz_dataOut_payload_0_12270 = (_zz_dataOut_payload_0_12247 < _zz_dataOut_payload_0_12259);
  assign _zz_dataOut_payload_0_12271 = (_zz_dataOut_payload_0_12270 ? _zz_dataOut_payload_0_12247 : _zz_dataOut_payload_0_12259);
  assign _zz_dataOut_payload_0_12272 = (_zz_dataOut_payload_0_12270 ? _zz_dataOut_payload_0_12259 : _zz_dataOut_payload_0_12247);
  assign _zz_dataOut_payload_0_12273 = (_zz_dataOut_payload_0_12250 < _zz_dataOut_payload_0_12262);
  assign _zz_dataOut_payload_0_12274 = (_zz_dataOut_payload_0_12273 ? _zz_dataOut_payload_0_12250 : _zz_dataOut_payload_0_12262);
  assign _zz_dataOut_payload_0_12275 = (_zz_dataOut_payload_0_12273 ? _zz_dataOut_payload_0_12262 : _zz_dataOut_payload_0_12250);
  assign _zz_dataOut_payload_0_12276 = (_zz_dataOut_payload_0_12265 < _zz_dataOut_payload_0_12271);
  assign _zz_dataOut_payload_0_12277 = (_zz_dataOut_payload_0_12276 ? _zz_dataOut_payload_0_12265 : _zz_dataOut_payload_0_12271);
  assign _zz_dataOut_payload_0_12278 = (_zz_dataOut_payload_0_12276 ? _zz_dataOut_payload_0_12271 : _zz_dataOut_payload_0_12265);
  assign _zz_dataOut_payload_0_12279 = (_zz_dataOut_payload_0_12268 < _zz_dataOut_payload_0_12274);
  assign _zz_dataOut_payload_0_12280 = (_zz_dataOut_payload_0_12279 ? _zz_dataOut_payload_0_12268 : _zz_dataOut_payload_0_12274);
  assign _zz_dataOut_payload_0_12281 = (_zz_dataOut_payload_0_12279 ? _zz_dataOut_payload_0_12274 : _zz_dataOut_payload_0_12268);
  assign _zz_dataOut_payload_0_12282 = (_zz_dataOut_payload_0_12277 < _zz_dataOut_payload_0_12280);
  assign _zz_dataOut_payload_0_12283 = (_zz_dataOut_payload_0_12278 < _zz_dataOut_payload_0_12281);
  assign _zz_dataOut_payload_0_12288 = (_zz_dataOut_payload_0_12266 < _zz_dataOut_payload_0_12272);
  assign _zz_dataOut_payload_0_12289 = (_zz_dataOut_payload_0_12288 ? _zz_dataOut_payload_0_12266 : _zz_dataOut_payload_0_12272);
  assign _zz_dataOut_payload_0_12290 = (_zz_dataOut_payload_0_12288 ? _zz_dataOut_payload_0_12272 : _zz_dataOut_payload_0_12266);
  assign _zz_dataOut_payload_0_12291 = (_zz_dataOut_payload_0_12269 < _zz_dataOut_payload_0_12275);
  assign _zz_dataOut_payload_0_12292 = (_zz_dataOut_payload_0_12291 ? _zz_dataOut_payload_0_12269 : _zz_dataOut_payload_0_12275);
  assign _zz_dataOut_payload_0_12293 = (_zz_dataOut_payload_0_12291 ? _zz_dataOut_payload_0_12275 : _zz_dataOut_payload_0_12269);
  assign _zz_dataOut_payload_0_12294 = (_zz_dataOut_payload_0_12289 < _zz_dataOut_payload_0_12292);
  assign _zz_dataOut_payload_0_12295 = (_zz_dataOut_payload_0_12290 < _zz_dataOut_payload_0_12293);
  assign _zz_dataOut_payload_0_12308 = (_zz_dataOut_payload_0_12242 < _zz_dataOut_payload_0_12254);
  assign _zz_dataOut_payload_0_12309 = (_zz_dataOut_payload_0_12308 ? _zz_dataOut_payload_0_12242 : _zz_dataOut_payload_0_12254);
  assign _zz_dataOut_payload_0_12310 = (_zz_dataOut_payload_0_12308 ? _zz_dataOut_payload_0_12254 : _zz_dataOut_payload_0_12242);
  assign _zz_dataOut_payload_0_12311 = (_zz_dataOut_payload_0_12245 < _zz_dataOut_payload_0_12257);
  assign _zz_dataOut_payload_0_12312 = (_zz_dataOut_payload_0_12311 ? _zz_dataOut_payload_0_12245 : _zz_dataOut_payload_0_12257);
  assign _zz_dataOut_payload_0_12313 = (_zz_dataOut_payload_0_12311 ? _zz_dataOut_payload_0_12257 : _zz_dataOut_payload_0_12245);
  assign _zz_dataOut_payload_0_12314 = (_zz_dataOut_payload_0_12248 < _zz_dataOut_payload_0_12260);
  assign _zz_dataOut_payload_0_12315 = (_zz_dataOut_payload_0_12314 ? _zz_dataOut_payload_0_12248 : _zz_dataOut_payload_0_12260);
  assign _zz_dataOut_payload_0_12316 = (_zz_dataOut_payload_0_12314 ? _zz_dataOut_payload_0_12260 : _zz_dataOut_payload_0_12248);
  assign _zz_dataOut_payload_0_12317 = (_zz_dataOut_payload_0_12251 < _zz_dataOut_payload_0_12263);
  assign _zz_dataOut_payload_0_12318 = (_zz_dataOut_payload_0_12317 ? _zz_dataOut_payload_0_12251 : _zz_dataOut_payload_0_12263);
  assign _zz_dataOut_payload_0_12319 = (_zz_dataOut_payload_0_12317 ? _zz_dataOut_payload_0_12263 : _zz_dataOut_payload_0_12251);
  assign _zz_dataOut_payload_0_12320 = (_zz_dataOut_payload_0_12309 < _zz_dataOut_payload_0_12315);
  assign _zz_dataOut_payload_0_12321 = (_zz_dataOut_payload_0_12320 ? _zz_dataOut_payload_0_12309 : _zz_dataOut_payload_0_12315);
  assign _zz_dataOut_payload_0_12322 = (_zz_dataOut_payload_0_12320 ? _zz_dataOut_payload_0_12315 : _zz_dataOut_payload_0_12309);
  assign _zz_dataOut_payload_0_12323 = (_zz_dataOut_payload_0_12312 < _zz_dataOut_payload_0_12318);
  assign _zz_dataOut_payload_0_12324 = (_zz_dataOut_payload_0_12323 ? _zz_dataOut_payload_0_12312 : _zz_dataOut_payload_0_12318);
  assign _zz_dataOut_payload_0_12325 = (_zz_dataOut_payload_0_12323 ? _zz_dataOut_payload_0_12318 : _zz_dataOut_payload_0_12312);
  assign _zz_dataOut_payload_0_12326 = (_zz_dataOut_payload_0_12321 < _zz_dataOut_payload_0_12324);
  assign _zz_dataOut_payload_0_12327 = (_zz_dataOut_payload_0_12322 < _zz_dataOut_payload_0_12325);
  assign _zz_dataOut_payload_0_12332 = (_zz_dataOut_payload_0_12310 < _zz_dataOut_payload_0_12316);
  assign _zz_dataOut_payload_0_12333 = (_zz_dataOut_payload_0_12332 ? _zz_dataOut_payload_0_12310 : _zz_dataOut_payload_0_12316);
  assign _zz_dataOut_payload_0_12334 = (_zz_dataOut_payload_0_12332 ? _zz_dataOut_payload_0_12316 : _zz_dataOut_payload_0_12310);
  assign _zz_dataOut_payload_0_12335 = (_zz_dataOut_payload_0_12313 < _zz_dataOut_payload_0_12319);
  assign _zz_dataOut_payload_0_12336 = (_zz_dataOut_payload_0_12335 ? _zz_dataOut_payload_0_12313 : _zz_dataOut_payload_0_12319);
  assign _zz_dataOut_payload_0_12337 = (_zz_dataOut_payload_0_12335 ? _zz_dataOut_payload_0_12319 : _zz_dataOut_payload_0_12313);
  assign _zz_dataOut_payload_0_12338 = (_zz_dataOut_payload_0_12333 < _zz_dataOut_payload_0_12336);
  assign _zz_dataOut_payload_0_12339 = (_zz_dataOut_payload_0_12334 < _zz_dataOut_payload_0_12337);
  assign _zz_dataOut_payload_0_12368 = (_zz_dataOut_payload_0_12194 < _zz_dataOut_payload_0_12218);
  assign _zz_dataOut_payload_0_12369 = (_zz_dataOut_payload_0_12368 ? _zz_dataOut_payload_0_12194 : _zz_dataOut_payload_0_12218);
  assign _zz_dataOut_payload_0_12370 = (_zz_dataOut_payload_0_12368 ? _zz_dataOut_payload_0_12218 : _zz_dataOut_payload_0_12194);
  assign _zz_dataOut_payload_0_12371 = (_zz_dataOut_payload_0_12197 < _zz_dataOut_payload_0_12221);
  assign _zz_dataOut_payload_0_12372 = (_zz_dataOut_payload_0_12371 ? _zz_dataOut_payload_0_12197 : _zz_dataOut_payload_0_12221);
  assign _zz_dataOut_payload_0_12373 = (_zz_dataOut_payload_0_12371 ? _zz_dataOut_payload_0_12221 : _zz_dataOut_payload_0_12197);
  assign _zz_dataOut_payload_0_12374 = (_zz_dataOut_payload_0_12200 < _zz_dataOut_payload_0_12224);
  assign _zz_dataOut_payload_0_12375 = (_zz_dataOut_payload_0_12374 ? _zz_dataOut_payload_0_12200 : _zz_dataOut_payload_0_12224);
  assign _zz_dataOut_payload_0_12376 = (_zz_dataOut_payload_0_12374 ? _zz_dataOut_payload_0_12224 : _zz_dataOut_payload_0_12200);
  assign _zz_dataOut_payload_0_12377 = (_zz_dataOut_payload_0_12203 < _zz_dataOut_payload_0_12227);
  assign _zz_dataOut_payload_0_12378 = (_zz_dataOut_payload_0_12377 ? _zz_dataOut_payload_0_12203 : _zz_dataOut_payload_0_12227);
  assign _zz_dataOut_payload_0_12379 = (_zz_dataOut_payload_0_12377 ? _zz_dataOut_payload_0_12227 : _zz_dataOut_payload_0_12203);
  assign _zz_dataOut_payload_0_12380 = (_zz_dataOut_payload_0_12206 < _zz_dataOut_payload_0_12230);
  assign _zz_dataOut_payload_0_12381 = (_zz_dataOut_payload_0_12380 ? _zz_dataOut_payload_0_12206 : _zz_dataOut_payload_0_12230);
  assign _zz_dataOut_payload_0_12382 = (_zz_dataOut_payload_0_12380 ? _zz_dataOut_payload_0_12230 : _zz_dataOut_payload_0_12206);
  assign _zz_dataOut_payload_0_12383 = (_zz_dataOut_payload_0_12209 < _zz_dataOut_payload_0_12233);
  assign _zz_dataOut_payload_0_12384 = (_zz_dataOut_payload_0_12383 ? _zz_dataOut_payload_0_12209 : _zz_dataOut_payload_0_12233);
  assign _zz_dataOut_payload_0_12385 = (_zz_dataOut_payload_0_12383 ? _zz_dataOut_payload_0_12233 : _zz_dataOut_payload_0_12209);
  assign _zz_dataOut_payload_0_12386 = (_zz_dataOut_payload_0_12212 < _zz_dataOut_payload_0_12236);
  assign _zz_dataOut_payload_0_12387 = (_zz_dataOut_payload_0_12386 ? _zz_dataOut_payload_0_12212 : _zz_dataOut_payload_0_12236);
  assign _zz_dataOut_payload_0_12388 = (_zz_dataOut_payload_0_12386 ? _zz_dataOut_payload_0_12236 : _zz_dataOut_payload_0_12212);
  assign _zz_dataOut_payload_0_12389 = (_zz_dataOut_payload_0_12215 < _zz_dataOut_payload_0_12239);
  assign _zz_dataOut_payload_0_12390 = (_zz_dataOut_payload_0_12389 ? _zz_dataOut_payload_0_12215 : _zz_dataOut_payload_0_12239);
  assign _zz_dataOut_payload_0_12391 = (_zz_dataOut_payload_0_12389 ? _zz_dataOut_payload_0_12239 : _zz_dataOut_payload_0_12215);
  assign _zz_dataOut_payload_0_12392 = (_zz_dataOut_payload_0_12369 < _zz_dataOut_payload_0_12381);
  assign _zz_dataOut_payload_0_12393 = (_zz_dataOut_payload_0_12392 ? _zz_dataOut_payload_0_12369 : _zz_dataOut_payload_0_12381);
  assign _zz_dataOut_payload_0_12394 = (_zz_dataOut_payload_0_12392 ? _zz_dataOut_payload_0_12381 : _zz_dataOut_payload_0_12369);
  assign _zz_dataOut_payload_0_12395 = (_zz_dataOut_payload_0_12372 < _zz_dataOut_payload_0_12384);
  assign _zz_dataOut_payload_0_12396 = (_zz_dataOut_payload_0_12395 ? _zz_dataOut_payload_0_12372 : _zz_dataOut_payload_0_12384);
  assign _zz_dataOut_payload_0_12397 = (_zz_dataOut_payload_0_12395 ? _zz_dataOut_payload_0_12384 : _zz_dataOut_payload_0_12372);
  assign _zz_dataOut_payload_0_12398 = (_zz_dataOut_payload_0_12375 < _zz_dataOut_payload_0_12387);
  assign _zz_dataOut_payload_0_12399 = (_zz_dataOut_payload_0_12398 ? _zz_dataOut_payload_0_12375 : _zz_dataOut_payload_0_12387);
  assign _zz_dataOut_payload_0_12400 = (_zz_dataOut_payload_0_12398 ? _zz_dataOut_payload_0_12387 : _zz_dataOut_payload_0_12375);
  assign _zz_dataOut_payload_0_12401 = (_zz_dataOut_payload_0_12378 < _zz_dataOut_payload_0_12390);
  assign _zz_dataOut_payload_0_12402 = (_zz_dataOut_payload_0_12401 ? _zz_dataOut_payload_0_12378 : _zz_dataOut_payload_0_12390);
  assign _zz_dataOut_payload_0_12403 = (_zz_dataOut_payload_0_12401 ? _zz_dataOut_payload_0_12390 : _zz_dataOut_payload_0_12378);
  assign _zz_dataOut_payload_0_12404 = (_zz_dataOut_payload_0_12393 < _zz_dataOut_payload_0_12399);
  assign _zz_dataOut_payload_0_12405 = (_zz_dataOut_payload_0_12404 ? _zz_dataOut_payload_0_12393 : _zz_dataOut_payload_0_12399);
  assign _zz_dataOut_payload_0_12406 = (_zz_dataOut_payload_0_12404 ? _zz_dataOut_payload_0_12399 : _zz_dataOut_payload_0_12393);
  assign _zz_dataOut_payload_0_12407 = (_zz_dataOut_payload_0_12396 < _zz_dataOut_payload_0_12402);
  assign _zz_dataOut_payload_0_12408 = (_zz_dataOut_payload_0_12407 ? _zz_dataOut_payload_0_12396 : _zz_dataOut_payload_0_12402);
  assign _zz_dataOut_payload_0_12409 = (_zz_dataOut_payload_0_12407 ? _zz_dataOut_payload_0_12402 : _zz_dataOut_payload_0_12396);
  assign _zz_dataOut_payload_0_12410 = (_zz_dataOut_payload_0_12405 < _zz_dataOut_payload_0_12408);
  assign _zz_dataOut_payload_0_12411 = (_zz_dataOut_payload_0_12406 < _zz_dataOut_payload_0_12409);
  assign _zz_dataOut_payload_0_12416 = (_zz_dataOut_payload_0_12394 < _zz_dataOut_payload_0_12400);
  assign _zz_dataOut_payload_0_12417 = (_zz_dataOut_payload_0_12416 ? _zz_dataOut_payload_0_12394 : _zz_dataOut_payload_0_12400);
  assign _zz_dataOut_payload_0_12418 = (_zz_dataOut_payload_0_12416 ? _zz_dataOut_payload_0_12400 : _zz_dataOut_payload_0_12394);
  assign _zz_dataOut_payload_0_12419 = (_zz_dataOut_payload_0_12397 < _zz_dataOut_payload_0_12403);
  assign _zz_dataOut_payload_0_12420 = (_zz_dataOut_payload_0_12419 ? _zz_dataOut_payload_0_12397 : _zz_dataOut_payload_0_12403);
  assign _zz_dataOut_payload_0_12421 = (_zz_dataOut_payload_0_12419 ? _zz_dataOut_payload_0_12403 : _zz_dataOut_payload_0_12397);
  assign _zz_dataOut_payload_0_12422 = (_zz_dataOut_payload_0_12417 < _zz_dataOut_payload_0_12420);
  assign _zz_dataOut_payload_0_12423 = (_zz_dataOut_payload_0_12418 < _zz_dataOut_payload_0_12421);
  assign _zz_dataOut_payload_0_12436 = (_zz_dataOut_payload_0_12370 < _zz_dataOut_payload_0_12382);
  assign _zz_dataOut_payload_0_12437 = (_zz_dataOut_payload_0_12436 ? _zz_dataOut_payload_0_12370 : _zz_dataOut_payload_0_12382);
  assign _zz_dataOut_payload_0_12438 = (_zz_dataOut_payload_0_12436 ? _zz_dataOut_payload_0_12382 : _zz_dataOut_payload_0_12370);
  assign _zz_dataOut_payload_0_12439 = (_zz_dataOut_payload_0_12373 < _zz_dataOut_payload_0_12385);
  assign _zz_dataOut_payload_0_12440 = (_zz_dataOut_payload_0_12439 ? _zz_dataOut_payload_0_12373 : _zz_dataOut_payload_0_12385);
  assign _zz_dataOut_payload_0_12441 = (_zz_dataOut_payload_0_12439 ? _zz_dataOut_payload_0_12385 : _zz_dataOut_payload_0_12373);
  assign _zz_dataOut_payload_0_12442 = (_zz_dataOut_payload_0_12376 < _zz_dataOut_payload_0_12388);
  assign _zz_dataOut_payload_0_12443 = (_zz_dataOut_payload_0_12442 ? _zz_dataOut_payload_0_12376 : _zz_dataOut_payload_0_12388);
  assign _zz_dataOut_payload_0_12444 = (_zz_dataOut_payload_0_12442 ? _zz_dataOut_payload_0_12388 : _zz_dataOut_payload_0_12376);
  assign _zz_dataOut_payload_0_12445 = (_zz_dataOut_payload_0_12379 < _zz_dataOut_payload_0_12391);
  assign _zz_dataOut_payload_0_12446 = (_zz_dataOut_payload_0_12445 ? _zz_dataOut_payload_0_12379 : _zz_dataOut_payload_0_12391);
  assign _zz_dataOut_payload_0_12447 = (_zz_dataOut_payload_0_12445 ? _zz_dataOut_payload_0_12391 : _zz_dataOut_payload_0_12379);
  assign _zz_dataOut_payload_0_12448 = (_zz_dataOut_payload_0_12437 < _zz_dataOut_payload_0_12443);
  assign _zz_dataOut_payload_0_12449 = (_zz_dataOut_payload_0_12448 ? _zz_dataOut_payload_0_12437 : _zz_dataOut_payload_0_12443);
  assign _zz_dataOut_payload_0_12450 = (_zz_dataOut_payload_0_12448 ? _zz_dataOut_payload_0_12443 : _zz_dataOut_payload_0_12437);
  assign _zz_dataOut_payload_0_12451 = (_zz_dataOut_payload_0_12440 < _zz_dataOut_payload_0_12446);
  assign _zz_dataOut_payload_0_12452 = (_zz_dataOut_payload_0_12451 ? _zz_dataOut_payload_0_12440 : _zz_dataOut_payload_0_12446);
  assign _zz_dataOut_payload_0_12453 = (_zz_dataOut_payload_0_12451 ? _zz_dataOut_payload_0_12446 : _zz_dataOut_payload_0_12440);
  assign _zz_dataOut_payload_0_12454 = (_zz_dataOut_payload_0_12449 < _zz_dataOut_payload_0_12452);
  assign _zz_dataOut_payload_0_12455 = (_zz_dataOut_payload_0_12450 < _zz_dataOut_payload_0_12453);
  assign _zz_dataOut_payload_0_12460 = (_zz_dataOut_payload_0_12438 < _zz_dataOut_payload_0_12444);
  assign _zz_dataOut_payload_0_12461 = (_zz_dataOut_payload_0_12460 ? _zz_dataOut_payload_0_12438 : _zz_dataOut_payload_0_12444);
  assign _zz_dataOut_payload_0_12462 = (_zz_dataOut_payload_0_12460 ? _zz_dataOut_payload_0_12444 : _zz_dataOut_payload_0_12438);
  assign _zz_dataOut_payload_0_12463 = (_zz_dataOut_payload_0_12441 < _zz_dataOut_payload_0_12447);
  assign _zz_dataOut_payload_0_12464 = (_zz_dataOut_payload_0_12463 ? _zz_dataOut_payload_0_12441 : _zz_dataOut_payload_0_12447);
  assign _zz_dataOut_payload_0_12465 = (_zz_dataOut_payload_0_12463 ? _zz_dataOut_payload_0_12447 : _zz_dataOut_payload_0_12441);
  assign _zz_dataOut_payload_0_12466 = (_zz_dataOut_payload_0_12461 < _zz_dataOut_payload_0_12464);
  assign _zz_dataOut_payload_0_12467 = (_zz_dataOut_payload_0_12462 < _zz_dataOut_payload_0_12465);
  assign _zz_dataOut_payload_0_12528 = (_zz_dataOut_payload_0_12098 < _zz_dataOut_payload_0_12146);
  assign _zz_dataOut_payload_0_12529 = (_zz_dataOut_payload_0_12528 ? _zz_dataOut_payload_0_12098 : _zz_dataOut_payload_0_12146);
  assign _zz_dataOut_payload_0_12530 = (_zz_dataOut_payload_0_12528 ? _zz_dataOut_payload_0_12146 : _zz_dataOut_payload_0_12098);
  assign _zz_dataOut_payload_0_12531 = (_zz_dataOut_payload_0_12101 < _zz_dataOut_payload_0_12149);
  assign _zz_dataOut_payload_0_12532 = (_zz_dataOut_payload_0_12531 ? _zz_dataOut_payload_0_12101 : _zz_dataOut_payload_0_12149);
  assign _zz_dataOut_payload_0_12533 = (_zz_dataOut_payload_0_12531 ? _zz_dataOut_payload_0_12149 : _zz_dataOut_payload_0_12101);
  assign _zz_dataOut_payload_0_12534 = (_zz_dataOut_payload_0_12104 < _zz_dataOut_payload_0_12152);
  assign _zz_dataOut_payload_0_12535 = (_zz_dataOut_payload_0_12534 ? _zz_dataOut_payload_0_12104 : _zz_dataOut_payload_0_12152);
  assign _zz_dataOut_payload_0_12536 = (_zz_dataOut_payload_0_12534 ? _zz_dataOut_payload_0_12152 : _zz_dataOut_payload_0_12104);
  assign _zz_dataOut_payload_0_12537 = (_zz_dataOut_payload_0_12107 < _zz_dataOut_payload_0_12155);
  assign _zz_dataOut_payload_0_12538 = (_zz_dataOut_payload_0_12537 ? _zz_dataOut_payload_0_12107 : _zz_dataOut_payload_0_12155);
  assign _zz_dataOut_payload_0_12539 = (_zz_dataOut_payload_0_12537 ? _zz_dataOut_payload_0_12155 : _zz_dataOut_payload_0_12107);
  assign _zz_dataOut_payload_0_12540 = (_zz_dataOut_payload_0_12110 < _zz_dataOut_payload_0_12158);
  assign _zz_dataOut_payload_0_12541 = (_zz_dataOut_payload_0_12540 ? _zz_dataOut_payload_0_12110 : _zz_dataOut_payload_0_12158);
  assign _zz_dataOut_payload_0_12542 = (_zz_dataOut_payload_0_12540 ? _zz_dataOut_payload_0_12158 : _zz_dataOut_payload_0_12110);
  assign _zz_dataOut_payload_0_12543 = (_zz_dataOut_payload_0_12113 < _zz_dataOut_payload_0_12161);
  assign _zz_dataOut_payload_0_12544 = (_zz_dataOut_payload_0_12543 ? _zz_dataOut_payload_0_12113 : _zz_dataOut_payload_0_12161);
  assign _zz_dataOut_payload_0_12545 = (_zz_dataOut_payload_0_12543 ? _zz_dataOut_payload_0_12161 : _zz_dataOut_payload_0_12113);
  assign _zz_dataOut_payload_0_12546 = (_zz_dataOut_payload_0_12116 < _zz_dataOut_payload_0_12164);
  assign _zz_dataOut_payload_0_12547 = (_zz_dataOut_payload_0_12546 ? _zz_dataOut_payload_0_12116 : _zz_dataOut_payload_0_12164);
  assign _zz_dataOut_payload_0_12548 = (_zz_dataOut_payload_0_12546 ? _zz_dataOut_payload_0_12164 : _zz_dataOut_payload_0_12116);
  assign _zz_dataOut_payload_0_12549 = (_zz_dataOut_payload_0_12119 < _zz_dataOut_payload_0_12167);
  assign _zz_dataOut_payload_0_12550 = (_zz_dataOut_payload_0_12549 ? _zz_dataOut_payload_0_12119 : _zz_dataOut_payload_0_12167);
  assign _zz_dataOut_payload_0_12551 = (_zz_dataOut_payload_0_12549 ? _zz_dataOut_payload_0_12167 : _zz_dataOut_payload_0_12119);
  assign _zz_dataOut_payload_0_12552 = (_zz_dataOut_payload_0_12122 < _zz_dataOut_payload_0_12170);
  assign _zz_dataOut_payload_0_12553 = (_zz_dataOut_payload_0_12552 ? _zz_dataOut_payload_0_12122 : _zz_dataOut_payload_0_12170);
  assign _zz_dataOut_payload_0_12554 = (_zz_dataOut_payload_0_12552 ? _zz_dataOut_payload_0_12170 : _zz_dataOut_payload_0_12122);
  assign _zz_dataOut_payload_0_12555 = (_zz_dataOut_payload_0_12125 < _zz_dataOut_payload_0_12173);
  assign _zz_dataOut_payload_0_12556 = (_zz_dataOut_payload_0_12555 ? _zz_dataOut_payload_0_12125 : _zz_dataOut_payload_0_12173);
  assign _zz_dataOut_payload_0_12557 = (_zz_dataOut_payload_0_12555 ? _zz_dataOut_payload_0_12173 : _zz_dataOut_payload_0_12125);
  assign _zz_dataOut_payload_0_12558 = (_zz_dataOut_payload_0_12128 < _zz_dataOut_payload_0_12176);
  assign _zz_dataOut_payload_0_12559 = (_zz_dataOut_payload_0_12558 ? _zz_dataOut_payload_0_12128 : _zz_dataOut_payload_0_12176);
  assign _zz_dataOut_payload_0_12560 = (_zz_dataOut_payload_0_12558 ? _zz_dataOut_payload_0_12176 : _zz_dataOut_payload_0_12128);
  assign _zz_dataOut_payload_0_12561 = (_zz_dataOut_payload_0_12131 < _zz_dataOut_payload_0_12179);
  assign _zz_dataOut_payload_0_12562 = (_zz_dataOut_payload_0_12561 ? _zz_dataOut_payload_0_12131 : _zz_dataOut_payload_0_12179);
  assign _zz_dataOut_payload_0_12563 = (_zz_dataOut_payload_0_12561 ? _zz_dataOut_payload_0_12179 : _zz_dataOut_payload_0_12131);
  assign _zz_dataOut_payload_0_12564 = (_zz_dataOut_payload_0_12134 < _zz_dataOut_payload_0_12182);
  assign _zz_dataOut_payload_0_12565 = (_zz_dataOut_payload_0_12564 ? _zz_dataOut_payload_0_12134 : _zz_dataOut_payload_0_12182);
  assign _zz_dataOut_payload_0_12566 = (_zz_dataOut_payload_0_12564 ? _zz_dataOut_payload_0_12182 : _zz_dataOut_payload_0_12134);
  assign _zz_dataOut_payload_0_12567 = (_zz_dataOut_payload_0_12137 < _zz_dataOut_payload_0_12185);
  assign _zz_dataOut_payload_0_12568 = (_zz_dataOut_payload_0_12567 ? _zz_dataOut_payload_0_12137 : _zz_dataOut_payload_0_12185);
  assign _zz_dataOut_payload_0_12569 = (_zz_dataOut_payload_0_12567 ? _zz_dataOut_payload_0_12185 : _zz_dataOut_payload_0_12137);
  assign _zz_dataOut_payload_0_12570 = (_zz_dataOut_payload_0_12140 < _zz_dataOut_payload_0_12188);
  assign _zz_dataOut_payload_0_12571 = (_zz_dataOut_payload_0_12570 ? _zz_dataOut_payload_0_12140 : _zz_dataOut_payload_0_12188);
  assign _zz_dataOut_payload_0_12572 = (_zz_dataOut_payload_0_12570 ? _zz_dataOut_payload_0_12188 : _zz_dataOut_payload_0_12140);
  assign _zz_dataOut_payload_0_12573 = (_zz_dataOut_payload_0_12143 < _zz_dataOut_payload_0_12191);
  assign _zz_dataOut_payload_0_12574 = (_zz_dataOut_payload_0_12573 ? _zz_dataOut_payload_0_12143 : _zz_dataOut_payload_0_12191);
  assign _zz_dataOut_payload_0_12575 = (_zz_dataOut_payload_0_12573 ? _zz_dataOut_payload_0_12191 : _zz_dataOut_payload_0_12143);
  assign _zz_dataOut_payload_0_12576 = (_zz_dataOut_payload_0_12529 < _zz_dataOut_payload_0_12553);
  assign _zz_dataOut_payload_0_12577 = (_zz_dataOut_payload_0_12576 ? _zz_dataOut_payload_0_12529 : _zz_dataOut_payload_0_12553);
  assign _zz_dataOut_payload_0_12578 = (_zz_dataOut_payload_0_12576 ? _zz_dataOut_payload_0_12553 : _zz_dataOut_payload_0_12529);
  assign _zz_dataOut_payload_0_12579 = (_zz_dataOut_payload_0_12532 < _zz_dataOut_payload_0_12556);
  assign _zz_dataOut_payload_0_12580 = (_zz_dataOut_payload_0_12579 ? _zz_dataOut_payload_0_12532 : _zz_dataOut_payload_0_12556);
  assign _zz_dataOut_payload_0_12581 = (_zz_dataOut_payload_0_12579 ? _zz_dataOut_payload_0_12556 : _zz_dataOut_payload_0_12532);
  assign _zz_dataOut_payload_0_12582 = (_zz_dataOut_payload_0_12535 < _zz_dataOut_payload_0_12559);
  assign _zz_dataOut_payload_0_12583 = (_zz_dataOut_payload_0_12582 ? _zz_dataOut_payload_0_12535 : _zz_dataOut_payload_0_12559);
  assign _zz_dataOut_payload_0_12584 = (_zz_dataOut_payload_0_12582 ? _zz_dataOut_payload_0_12559 : _zz_dataOut_payload_0_12535);
  assign _zz_dataOut_payload_0_12585 = (_zz_dataOut_payload_0_12538 < _zz_dataOut_payload_0_12562);
  assign _zz_dataOut_payload_0_12586 = (_zz_dataOut_payload_0_12585 ? _zz_dataOut_payload_0_12538 : _zz_dataOut_payload_0_12562);
  assign _zz_dataOut_payload_0_12587 = (_zz_dataOut_payload_0_12585 ? _zz_dataOut_payload_0_12562 : _zz_dataOut_payload_0_12538);
  assign _zz_dataOut_payload_0_12588 = (_zz_dataOut_payload_0_12541 < _zz_dataOut_payload_0_12565);
  assign _zz_dataOut_payload_0_12589 = (_zz_dataOut_payload_0_12588 ? _zz_dataOut_payload_0_12541 : _zz_dataOut_payload_0_12565);
  assign _zz_dataOut_payload_0_12590 = (_zz_dataOut_payload_0_12588 ? _zz_dataOut_payload_0_12565 : _zz_dataOut_payload_0_12541);
  assign _zz_dataOut_payload_0_12591 = (_zz_dataOut_payload_0_12544 < _zz_dataOut_payload_0_12568);
  assign _zz_dataOut_payload_0_12592 = (_zz_dataOut_payload_0_12591 ? _zz_dataOut_payload_0_12544 : _zz_dataOut_payload_0_12568);
  assign _zz_dataOut_payload_0_12593 = (_zz_dataOut_payload_0_12591 ? _zz_dataOut_payload_0_12568 : _zz_dataOut_payload_0_12544);
  assign _zz_dataOut_payload_0_12594 = (_zz_dataOut_payload_0_12547 < _zz_dataOut_payload_0_12571);
  assign _zz_dataOut_payload_0_12595 = (_zz_dataOut_payload_0_12594 ? _zz_dataOut_payload_0_12547 : _zz_dataOut_payload_0_12571);
  assign _zz_dataOut_payload_0_12596 = (_zz_dataOut_payload_0_12594 ? _zz_dataOut_payload_0_12571 : _zz_dataOut_payload_0_12547);
  assign _zz_dataOut_payload_0_12597 = (_zz_dataOut_payload_0_12550 < _zz_dataOut_payload_0_12574);
  assign _zz_dataOut_payload_0_12598 = (_zz_dataOut_payload_0_12597 ? _zz_dataOut_payload_0_12550 : _zz_dataOut_payload_0_12574);
  assign _zz_dataOut_payload_0_12599 = (_zz_dataOut_payload_0_12597 ? _zz_dataOut_payload_0_12574 : _zz_dataOut_payload_0_12550);
  assign _zz_dataOut_payload_0_12600 = (_zz_dataOut_payload_0_12577 < _zz_dataOut_payload_0_12589);
  assign _zz_dataOut_payload_0_12601 = (_zz_dataOut_payload_0_12600 ? _zz_dataOut_payload_0_12577 : _zz_dataOut_payload_0_12589);
  assign _zz_dataOut_payload_0_12602 = (_zz_dataOut_payload_0_12600 ? _zz_dataOut_payload_0_12589 : _zz_dataOut_payload_0_12577);
  assign _zz_dataOut_payload_0_12603 = (_zz_dataOut_payload_0_12580 < _zz_dataOut_payload_0_12592);
  assign _zz_dataOut_payload_0_12604 = (_zz_dataOut_payload_0_12603 ? _zz_dataOut_payload_0_12580 : _zz_dataOut_payload_0_12592);
  assign _zz_dataOut_payload_0_12605 = (_zz_dataOut_payload_0_12603 ? _zz_dataOut_payload_0_12592 : _zz_dataOut_payload_0_12580);
  assign _zz_dataOut_payload_0_12606 = (_zz_dataOut_payload_0_12583 < _zz_dataOut_payload_0_12595);
  assign _zz_dataOut_payload_0_12607 = (_zz_dataOut_payload_0_12606 ? _zz_dataOut_payload_0_12583 : _zz_dataOut_payload_0_12595);
  assign _zz_dataOut_payload_0_12608 = (_zz_dataOut_payload_0_12606 ? _zz_dataOut_payload_0_12595 : _zz_dataOut_payload_0_12583);
  assign _zz_dataOut_payload_0_12609 = (_zz_dataOut_payload_0_12586 < _zz_dataOut_payload_0_12598);
  assign _zz_dataOut_payload_0_12610 = (_zz_dataOut_payload_0_12609 ? _zz_dataOut_payload_0_12586 : _zz_dataOut_payload_0_12598);
  assign _zz_dataOut_payload_0_12611 = (_zz_dataOut_payload_0_12609 ? _zz_dataOut_payload_0_12598 : _zz_dataOut_payload_0_12586);
  assign _zz_dataOut_payload_0_12612 = (_zz_dataOut_payload_0_12601 < _zz_dataOut_payload_0_12607);
  assign _zz_dataOut_payload_0_12613 = (_zz_dataOut_payload_0_12612 ? _zz_dataOut_payload_0_12601 : _zz_dataOut_payload_0_12607);
  assign _zz_dataOut_payload_0_12614 = (_zz_dataOut_payload_0_12612 ? _zz_dataOut_payload_0_12607 : _zz_dataOut_payload_0_12601);
  assign _zz_dataOut_payload_0_12615 = (_zz_dataOut_payload_0_12604 < _zz_dataOut_payload_0_12610);
  assign _zz_dataOut_payload_0_12616 = (_zz_dataOut_payload_0_12615 ? _zz_dataOut_payload_0_12604 : _zz_dataOut_payload_0_12610);
  assign _zz_dataOut_payload_0_12617 = (_zz_dataOut_payload_0_12615 ? _zz_dataOut_payload_0_12610 : _zz_dataOut_payload_0_12604);
  assign _zz_dataOut_payload_0_12618 = (_zz_dataOut_payload_0_12613 < _zz_dataOut_payload_0_12616);
  assign _zz_dataOut_payload_0_12619 = (_zz_dataOut_payload_0_12614 < _zz_dataOut_payload_0_12617);
  assign _zz_dataOut_payload_0_12624 = (_zz_dataOut_payload_0_12602 < _zz_dataOut_payload_0_12608);
  assign _zz_dataOut_payload_0_12625 = (_zz_dataOut_payload_0_12624 ? _zz_dataOut_payload_0_12602 : _zz_dataOut_payload_0_12608);
  assign _zz_dataOut_payload_0_12626 = (_zz_dataOut_payload_0_12624 ? _zz_dataOut_payload_0_12608 : _zz_dataOut_payload_0_12602);
  assign _zz_dataOut_payload_0_12627 = (_zz_dataOut_payload_0_12605 < _zz_dataOut_payload_0_12611);
  assign _zz_dataOut_payload_0_12628 = (_zz_dataOut_payload_0_12627 ? _zz_dataOut_payload_0_12605 : _zz_dataOut_payload_0_12611);
  assign _zz_dataOut_payload_0_12629 = (_zz_dataOut_payload_0_12627 ? _zz_dataOut_payload_0_12611 : _zz_dataOut_payload_0_12605);
  assign _zz_dataOut_payload_0_12630 = (_zz_dataOut_payload_0_12625 < _zz_dataOut_payload_0_12628);
  assign _zz_dataOut_payload_0_12631 = (_zz_dataOut_payload_0_12626 < _zz_dataOut_payload_0_12629);
  assign _zz_dataOut_payload_0_12644 = (_zz_dataOut_payload_0_12578 < _zz_dataOut_payload_0_12590);
  assign _zz_dataOut_payload_0_12645 = (_zz_dataOut_payload_0_12644 ? _zz_dataOut_payload_0_12578 : _zz_dataOut_payload_0_12590);
  assign _zz_dataOut_payload_0_12646 = (_zz_dataOut_payload_0_12644 ? _zz_dataOut_payload_0_12590 : _zz_dataOut_payload_0_12578);
  assign _zz_dataOut_payload_0_12647 = (_zz_dataOut_payload_0_12581 < _zz_dataOut_payload_0_12593);
  assign _zz_dataOut_payload_0_12648 = (_zz_dataOut_payload_0_12647 ? _zz_dataOut_payload_0_12581 : _zz_dataOut_payload_0_12593);
  assign _zz_dataOut_payload_0_12649 = (_zz_dataOut_payload_0_12647 ? _zz_dataOut_payload_0_12593 : _zz_dataOut_payload_0_12581);
  assign _zz_dataOut_payload_0_12650 = (_zz_dataOut_payload_0_12584 < _zz_dataOut_payload_0_12596);
  assign _zz_dataOut_payload_0_12651 = (_zz_dataOut_payload_0_12650 ? _zz_dataOut_payload_0_12584 : _zz_dataOut_payload_0_12596);
  assign _zz_dataOut_payload_0_12652 = (_zz_dataOut_payload_0_12650 ? _zz_dataOut_payload_0_12596 : _zz_dataOut_payload_0_12584);
  assign _zz_dataOut_payload_0_12653 = (_zz_dataOut_payload_0_12587 < _zz_dataOut_payload_0_12599);
  assign _zz_dataOut_payload_0_12654 = (_zz_dataOut_payload_0_12653 ? _zz_dataOut_payload_0_12587 : _zz_dataOut_payload_0_12599);
  assign _zz_dataOut_payload_0_12655 = (_zz_dataOut_payload_0_12653 ? _zz_dataOut_payload_0_12599 : _zz_dataOut_payload_0_12587);
  assign _zz_dataOut_payload_0_12656 = (_zz_dataOut_payload_0_12645 < _zz_dataOut_payload_0_12651);
  assign _zz_dataOut_payload_0_12657 = (_zz_dataOut_payload_0_12656 ? _zz_dataOut_payload_0_12645 : _zz_dataOut_payload_0_12651);
  assign _zz_dataOut_payload_0_12658 = (_zz_dataOut_payload_0_12656 ? _zz_dataOut_payload_0_12651 : _zz_dataOut_payload_0_12645);
  assign _zz_dataOut_payload_0_12659 = (_zz_dataOut_payload_0_12648 < _zz_dataOut_payload_0_12654);
  assign _zz_dataOut_payload_0_12660 = (_zz_dataOut_payload_0_12659 ? _zz_dataOut_payload_0_12648 : _zz_dataOut_payload_0_12654);
  assign _zz_dataOut_payload_0_12661 = (_zz_dataOut_payload_0_12659 ? _zz_dataOut_payload_0_12654 : _zz_dataOut_payload_0_12648);
  assign _zz_dataOut_payload_0_12662 = (_zz_dataOut_payload_0_12657 < _zz_dataOut_payload_0_12660);
  assign _zz_dataOut_payload_0_12663 = (_zz_dataOut_payload_0_12658 < _zz_dataOut_payload_0_12661);
  assign _zz_dataOut_payload_0_12668 = (_zz_dataOut_payload_0_12646 < _zz_dataOut_payload_0_12652);
  assign _zz_dataOut_payload_0_12669 = (_zz_dataOut_payload_0_12668 ? _zz_dataOut_payload_0_12646 : _zz_dataOut_payload_0_12652);
  assign _zz_dataOut_payload_0_12670 = (_zz_dataOut_payload_0_12668 ? _zz_dataOut_payload_0_12652 : _zz_dataOut_payload_0_12646);
  assign _zz_dataOut_payload_0_12671 = (_zz_dataOut_payload_0_12649 < _zz_dataOut_payload_0_12655);
  assign _zz_dataOut_payload_0_12672 = (_zz_dataOut_payload_0_12671 ? _zz_dataOut_payload_0_12649 : _zz_dataOut_payload_0_12655);
  assign _zz_dataOut_payload_0_12673 = (_zz_dataOut_payload_0_12671 ? _zz_dataOut_payload_0_12655 : _zz_dataOut_payload_0_12649);
  assign _zz_dataOut_payload_0_12674 = (_zz_dataOut_payload_0_12669 < _zz_dataOut_payload_0_12672);
  assign _zz_dataOut_payload_0_12675 = (_zz_dataOut_payload_0_12670 < _zz_dataOut_payload_0_12673);
  assign _zz_dataOut_payload_0_12704 = (_zz_dataOut_payload_0_12530 < _zz_dataOut_payload_0_12554);
  assign _zz_dataOut_payload_0_12705 = (_zz_dataOut_payload_0_12704 ? _zz_dataOut_payload_0_12530 : _zz_dataOut_payload_0_12554);
  assign _zz_dataOut_payload_0_12706 = (_zz_dataOut_payload_0_12704 ? _zz_dataOut_payload_0_12554 : _zz_dataOut_payload_0_12530);
  assign _zz_dataOut_payload_0_12707 = (_zz_dataOut_payload_0_12533 < _zz_dataOut_payload_0_12557);
  assign _zz_dataOut_payload_0_12708 = (_zz_dataOut_payload_0_12707 ? _zz_dataOut_payload_0_12533 : _zz_dataOut_payload_0_12557);
  assign _zz_dataOut_payload_0_12709 = (_zz_dataOut_payload_0_12707 ? _zz_dataOut_payload_0_12557 : _zz_dataOut_payload_0_12533);
  assign _zz_dataOut_payload_0_12710 = (_zz_dataOut_payload_0_12536 < _zz_dataOut_payload_0_12560);
  assign _zz_dataOut_payload_0_12711 = (_zz_dataOut_payload_0_12710 ? _zz_dataOut_payload_0_12536 : _zz_dataOut_payload_0_12560);
  assign _zz_dataOut_payload_0_12712 = (_zz_dataOut_payload_0_12710 ? _zz_dataOut_payload_0_12560 : _zz_dataOut_payload_0_12536);
  assign _zz_dataOut_payload_0_12713 = (_zz_dataOut_payload_0_12539 < _zz_dataOut_payload_0_12563);
  assign _zz_dataOut_payload_0_12714 = (_zz_dataOut_payload_0_12713 ? _zz_dataOut_payload_0_12539 : _zz_dataOut_payload_0_12563);
  assign _zz_dataOut_payload_0_12715 = (_zz_dataOut_payload_0_12713 ? _zz_dataOut_payload_0_12563 : _zz_dataOut_payload_0_12539);
  assign _zz_dataOut_payload_0_12716 = (_zz_dataOut_payload_0_12542 < _zz_dataOut_payload_0_12566);
  assign _zz_dataOut_payload_0_12717 = (_zz_dataOut_payload_0_12716 ? _zz_dataOut_payload_0_12542 : _zz_dataOut_payload_0_12566);
  assign _zz_dataOut_payload_0_12718 = (_zz_dataOut_payload_0_12716 ? _zz_dataOut_payload_0_12566 : _zz_dataOut_payload_0_12542);
  assign _zz_dataOut_payload_0_12719 = (_zz_dataOut_payload_0_12545 < _zz_dataOut_payload_0_12569);
  assign _zz_dataOut_payload_0_12720 = (_zz_dataOut_payload_0_12719 ? _zz_dataOut_payload_0_12545 : _zz_dataOut_payload_0_12569);
  assign _zz_dataOut_payload_0_12721 = (_zz_dataOut_payload_0_12719 ? _zz_dataOut_payload_0_12569 : _zz_dataOut_payload_0_12545);
  assign _zz_dataOut_payload_0_12722 = (_zz_dataOut_payload_0_12548 < _zz_dataOut_payload_0_12572);
  assign _zz_dataOut_payload_0_12723 = (_zz_dataOut_payload_0_12722 ? _zz_dataOut_payload_0_12548 : _zz_dataOut_payload_0_12572);
  assign _zz_dataOut_payload_0_12724 = (_zz_dataOut_payload_0_12722 ? _zz_dataOut_payload_0_12572 : _zz_dataOut_payload_0_12548);
  assign _zz_dataOut_payload_0_12725 = (_zz_dataOut_payload_0_12551 < _zz_dataOut_payload_0_12575);
  assign _zz_dataOut_payload_0_12726 = (_zz_dataOut_payload_0_12725 ? _zz_dataOut_payload_0_12551 : _zz_dataOut_payload_0_12575);
  assign _zz_dataOut_payload_0_12727 = (_zz_dataOut_payload_0_12725 ? _zz_dataOut_payload_0_12575 : _zz_dataOut_payload_0_12551);
  assign _zz_dataOut_payload_0_12728 = (_zz_dataOut_payload_0_12705 < _zz_dataOut_payload_0_12717);
  assign _zz_dataOut_payload_0_12729 = (_zz_dataOut_payload_0_12728 ? _zz_dataOut_payload_0_12705 : _zz_dataOut_payload_0_12717);
  assign _zz_dataOut_payload_0_12730 = (_zz_dataOut_payload_0_12728 ? _zz_dataOut_payload_0_12717 : _zz_dataOut_payload_0_12705);
  assign _zz_dataOut_payload_0_12731 = (_zz_dataOut_payload_0_12708 < _zz_dataOut_payload_0_12720);
  assign _zz_dataOut_payload_0_12732 = (_zz_dataOut_payload_0_12731 ? _zz_dataOut_payload_0_12708 : _zz_dataOut_payload_0_12720);
  assign _zz_dataOut_payload_0_12733 = (_zz_dataOut_payload_0_12731 ? _zz_dataOut_payload_0_12720 : _zz_dataOut_payload_0_12708);
  assign _zz_dataOut_payload_0_12734 = (_zz_dataOut_payload_0_12711 < _zz_dataOut_payload_0_12723);
  assign _zz_dataOut_payload_0_12735 = (_zz_dataOut_payload_0_12734 ? _zz_dataOut_payload_0_12711 : _zz_dataOut_payload_0_12723);
  assign _zz_dataOut_payload_0_12736 = (_zz_dataOut_payload_0_12734 ? _zz_dataOut_payload_0_12723 : _zz_dataOut_payload_0_12711);
  assign _zz_dataOut_payload_0_12737 = (_zz_dataOut_payload_0_12714 < _zz_dataOut_payload_0_12726);
  assign _zz_dataOut_payload_0_12738 = (_zz_dataOut_payload_0_12737 ? _zz_dataOut_payload_0_12714 : _zz_dataOut_payload_0_12726);
  assign _zz_dataOut_payload_0_12739 = (_zz_dataOut_payload_0_12737 ? _zz_dataOut_payload_0_12726 : _zz_dataOut_payload_0_12714);
  assign _zz_dataOut_payload_0_12740 = (_zz_dataOut_payload_0_12729 < _zz_dataOut_payload_0_12735);
  assign _zz_dataOut_payload_0_12741 = (_zz_dataOut_payload_0_12740 ? _zz_dataOut_payload_0_12729 : _zz_dataOut_payload_0_12735);
  assign _zz_dataOut_payload_0_12742 = (_zz_dataOut_payload_0_12740 ? _zz_dataOut_payload_0_12735 : _zz_dataOut_payload_0_12729);
  assign _zz_dataOut_payload_0_12743 = (_zz_dataOut_payload_0_12732 < _zz_dataOut_payload_0_12738);
  assign _zz_dataOut_payload_0_12744 = (_zz_dataOut_payload_0_12743 ? _zz_dataOut_payload_0_12732 : _zz_dataOut_payload_0_12738);
  assign _zz_dataOut_payload_0_12745 = (_zz_dataOut_payload_0_12743 ? _zz_dataOut_payload_0_12738 : _zz_dataOut_payload_0_12732);
  assign _zz_dataOut_payload_0_12746 = (_zz_dataOut_payload_0_12741 < _zz_dataOut_payload_0_12744);
  assign _zz_dataOut_payload_0_12747 = (_zz_dataOut_payload_0_12742 < _zz_dataOut_payload_0_12745);
  assign _zz_dataOut_payload_0_12752 = (_zz_dataOut_payload_0_12730 < _zz_dataOut_payload_0_12736);
  assign _zz_dataOut_payload_0_12753 = (_zz_dataOut_payload_0_12752 ? _zz_dataOut_payload_0_12730 : _zz_dataOut_payload_0_12736);
  assign _zz_dataOut_payload_0_12754 = (_zz_dataOut_payload_0_12752 ? _zz_dataOut_payload_0_12736 : _zz_dataOut_payload_0_12730);
  assign _zz_dataOut_payload_0_12755 = (_zz_dataOut_payload_0_12733 < _zz_dataOut_payload_0_12739);
  assign _zz_dataOut_payload_0_12756 = (_zz_dataOut_payload_0_12755 ? _zz_dataOut_payload_0_12733 : _zz_dataOut_payload_0_12739);
  assign _zz_dataOut_payload_0_12757 = (_zz_dataOut_payload_0_12755 ? _zz_dataOut_payload_0_12739 : _zz_dataOut_payload_0_12733);
  assign _zz_dataOut_payload_0_12758 = (_zz_dataOut_payload_0_12753 < _zz_dataOut_payload_0_12756);
  assign _zz_dataOut_payload_0_12759 = (_zz_dataOut_payload_0_12754 < _zz_dataOut_payload_0_12757);
  assign _zz_dataOut_payload_0_12772 = (_zz_dataOut_payload_0_12706 < _zz_dataOut_payload_0_12718);
  assign _zz_dataOut_payload_0_12773 = (_zz_dataOut_payload_0_12772 ? _zz_dataOut_payload_0_12706 : _zz_dataOut_payload_0_12718);
  assign _zz_dataOut_payload_0_12774 = (_zz_dataOut_payload_0_12772 ? _zz_dataOut_payload_0_12718 : _zz_dataOut_payload_0_12706);
  assign _zz_dataOut_payload_0_12775 = (_zz_dataOut_payload_0_12709 < _zz_dataOut_payload_0_12721);
  assign _zz_dataOut_payload_0_12776 = (_zz_dataOut_payload_0_12775 ? _zz_dataOut_payload_0_12709 : _zz_dataOut_payload_0_12721);
  assign _zz_dataOut_payload_0_12777 = (_zz_dataOut_payload_0_12775 ? _zz_dataOut_payload_0_12721 : _zz_dataOut_payload_0_12709);
  assign _zz_dataOut_payload_0_12778 = (_zz_dataOut_payload_0_12712 < _zz_dataOut_payload_0_12724);
  assign _zz_dataOut_payload_0_12779 = (_zz_dataOut_payload_0_12778 ? _zz_dataOut_payload_0_12712 : _zz_dataOut_payload_0_12724);
  assign _zz_dataOut_payload_0_12780 = (_zz_dataOut_payload_0_12778 ? _zz_dataOut_payload_0_12724 : _zz_dataOut_payload_0_12712);
  assign _zz_dataOut_payload_0_12781 = (_zz_dataOut_payload_0_12715 < _zz_dataOut_payload_0_12727);
  assign _zz_dataOut_payload_0_12782 = (_zz_dataOut_payload_0_12781 ? _zz_dataOut_payload_0_12715 : _zz_dataOut_payload_0_12727);
  assign _zz_dataOut_payload_0_12783 = (_zz_dataOut_payload_0_12781 ? _zz_dataOut_payload_0_12727 : _zz_dataOut_payload_0_12715);
  assign _zz_dataOut_payload_0_12784 = (_zz_dataOut_payload_0_12773 < _zz_dataOut_payload_0_12779);
  assign _zz_dataOut_payload_0_12785 = (_zz_dataOut_payload_0_12784 ? _zz_dataOut_payload_0_12773 : _zz_dataOut_payload_0_12779);
  assign _zz_dataOut_payload_0_12786 = (_zz_dataOut_payload_0_12784 ? _zz_dataOut_payload_0_12779 : _zz_dataOut_payload_0_12773);
  assign _zz_dataOut_payload_0_12787 = (_zz_dataOut_payload_0_12776 < _zz_dataOut_payload_0_12782);
  assign _zz_dataOut_payload_0_12788 = (_zz_dataOut_payload_0_12787 ? _zz_dataOut_payload_0_12776 : _zz_dataOut_payload_0_12782);
  assign _zz_dataOut_payload_0_12789 = (_zz_dataOut_payload_0_12787 ? _zz_dataOut_payload_0_12782 : _zz_dataOut_payload_0_12776);
  assign _zz_dataOut_payload_0_12790 = (_zz_dataOut_payload_0_12785 < _zz_dataOut_payload_0_12788);
  assign _zz_dataOut_payload_0_12791 = (_zz_dataOut_payload_0_12786 < _zz_dataOut_payload_0_12789);
  assign _zz_dataOut_payload_0_12796 = (_zz_dataOut_payload_0_12774 < _zz_dataOut_payload_0_12780);
  assign _zz_dataOut_payload_0_12797 = (_zz_dataOut_payload_0_12796 ? _zz_dataOut_payload_0_12774 : _zz_dataOut_payload_0_12780);
  assign _zz_dataOut_payload_0_12798 = (_zz_dataOut_payload_0_12796 ? _zz_dataOut_payload_0_12780 : _zz_dataOut_payload_0_12774);
  assign _zz_dataOut_payload_0_12799 = (_zz_dataOut_payload_0_12777 < _zz_dataOut_payload_0_12783);
  assign _zz_dataOut_payload_0_12800 = (_zz_dataOut_payload_0_12799 ? _zz_dataOut_payload_0_12777 : _zz_dataOut_payload_0_12783);
  assign _zz_dataOut_payload_0_12801 = (_zz_dataOut_payload_0_12799 ? _zz_dataOut_payload_0_12783 : _zz_dataOut_payload_0_12777);
  assign _zz_dataOut_payload_0_12802 = (_zz_dataOut_payload_0_12797 < _zz_dataOut_payload_0_12800);
  assign _zz_dataOut_payload_0_12803 = (_zz_dataOut_payload_0_12798 < _zz_dataOut_payload_0_12801);
  assign _zz_dataOut_payload_0_12928 = (_zz_dataOut_payload_0_12095 < _zz_dataOut_payload_0_11999);
  assign _zz_dataOut_payload_0_12929 = (_zz_dataOut_payload_0_12928 ? _zz_dataOut_payload_0_12095 : _zz_dataOut_payload_0_11999);
  assign _zz_dataOut_payload_0_12930 = (_zz_dataOut_payload_0_12928 ? _zz_dataOut_payload_0_11999 : _zz_dataOut_payload_0_12095);
  assign _zz_dataOut_payload_0_12931 = (_zz_dataOut_payload_0_12092 < _zz_dataOut_payload_0_11996);
  assign _zz_dataOut_payload_0_12932 = (_zz_dataOut_payload_0_12931 ? _zz_dataOut_payload_0_12092 : _zz_dataOut_payload_0_11996);
  assign _zz_dataOut_payload_0_12933 = (_zz_dataOut_payload_0_12931 ? _zz_dataOut_payload_0_11996 : _zz_dataOut_payload_0_12092);
  assign _zz_dataOut_payload_0_12934 = (_zz_dataOut_payload_0_12089 < _zz_dataOut_payload_0_11993);
  assign _zz_dataOut_payload_0_12935 = (_zz_dataOut_payload_0_12934 ? _zz_dataOut_payload_0_12089 : _zz_dataOut_payload_0_11993);
  assign _zz_dataOut_payload_0_12936 = (_zz_dataOut_payload_0_12934 ? _zz_dataOut_payload_0_11993 : _zz_dataOut_payload_0_12089);
  assign _zz_dataOut_payload_0_12937 = (_zz_dataOut_payload_0_12086 < _zz_dataOut_payload_0_11990);
  assign _zz_dataOut_payload_0_12938 = (_zz_dataOut_payload_0_12937 ? _zz_dataOut_payload_0_12086 : _zz_dataOut_payload_0_11990);
  assign _zz_dataOut_payload_0_12939 = (_zz_dataOut_payload_0_12937 ? _zz_dataOut_payload_0_11990 : _zz_dataOut_payload_0_12086);
  assign _zz_dataOut_payload_0_12940 = (_zz_dataOut_payload_0_12083 < _zz_dataOut_payload_0_11987);
  assign _zz_dataOut_payload_0_12941 = (_zz_dataOut_payload_0_12940 ? _zz_dataOut_payload_0_12083 : _zz_dataOut_payload_0_11987);
  assign _zz_dataOut_payload_0_12942 = (_zz_dataOut_payload_0_12940 ? _zz_dataOut_payload_0_11987 : _zz_dataOut_payload_0_12083);
  assign _zz_dataOut_payload_0_12943 = (_zz_dataOut_payload_0_12080 < _zz_dataOut_payload_0_11984);
  assign _zz_dataOut_payload_0_12944 = (_zz_dataOut_payload_0_12943 ? _zz_dataOut_payload_0_12080 : _zz_dataOut_payload_0_11984);
  assign _zz_dataOut_payload_0_12945 = (_zz_dataOut_payload_0_12943 ? _zz_dataOut_payload_0_11984 : _zz_dataOut_payload_0_12080);
  assign _zz_dataOut_payload_0_12946 = (_zz_dataOut_payload_0_12077 < _zz_dataOut_payload_0_11981);
  assign _zz_dataOut_payload_0_12947 = (_zz_dataOut_payload_0_12946 ? _zz_dataOut_payload_0_12077 : _zz_dataOut_payload_0_11981);
  assign _zz_dataOut_payload_0_12948 = (_zz_dataOut_payload_0_12946 ? _zz_dataOut_payload_0_11981 : _zz_dataOut_payload_0_12077);
  assign _zz_dataOut_payload_0_12949 = (_zz_dataOut_payload_0_12074 < _zz_dataOut_payload_0_11978);
  assign _zz_dataOut_payload_0_12950 = (_zz_dataOut_payload_0_12949 ? _zz_dataOut_payload_0_12074 : _zz_dataOut_payload_0_11978);
  assign _zz_dataOut_payload_0_12951 = (_zz_dataOut_payload_0_12949 ? _zz_dataOut_payload_0_11978 : _zz_dataOut_payload_0_12074);
  assign _zz_dataOut_payload_0_12952 = (_zz_dataOut_payload_0_12071 < _zz_dataOut_payload_0_11975);
  assign _zz_dataOut_payload_0_12953 = (_zz_dataOut_payload_0_12952 ? _zz_dataOut_payload_0_12071 : _zz_dataOut_payload_0_11975);
  assign _zz_dataOut_payload_0_12954 = (_zz_dataOut_payload_0_12952 ? _zz_dataOut_payload_0_11975 : _zz_dataOut_payload_0_12071);
  assign _zz_dataOut_payload_0_12955 = (_zz_dataOut_payload_0_12068 < _zz_dataOut_payload_0_11972);
  assign _zz_dataOut_payload_0_12956 = (_zz_dataOut_payload_0_12955 ? _zz_dataOut_payload_0_12068 : _zz_dataOut_payload_0_11972);
  assign _zz_dataOut_payload_0_12957 = (_zz_dataOut_payload_0_12955 ? _zz_dataOut_payload_0_11972 : _zz_dataOut_payload_0_12068);
  assign _zz_dataOut_payload_0_12958 = (_zz_dataOut_payload_0_12065 < _zz_dataOut_payload_0_11969);
  assign _zz_dataOut_payload_0_12959 = (_zz_dataOut_payload_0_12958 ? _zz_dataOut_payload_0_12065 : _zz_dataOut_payload_0_11969);
  assign _zz_dataOut_payload_0_12960 = (_zz_dataOut_payload_0_12958 ? _zz_dataOut_payload_0_11969 : _zz_dataOut_payload_0_12065);
  assign _zz_dataOut_payload_0_12961 = (_zz_dataOut_payload_0_12062 < _zz_dataOut_payload_0_11966);
  assign _zz_dataOut_payload_0_12962 = (_zz_dataOut_payload_0_12961 ? _zz_dataOut_payload_0_12062 : _zz_dataOut_payload_0_11966);
  assign _zz_dataOut_payload_0_12963 = (_zz_dataOut_payload_0_12961 ? _zz_dataOut_payload_0_11966 : _zz_dataOut_payload_0_12062);
  assign _zz_dataOut_payload_0_12964 = (_zz_dataOut_payload_0_12059 < _zz_dataOut_payload_0_11963);
  assign _zz_dataOut_payload_0_12965 = (_zz_dataOut_payload_0_12964 ? _zz_dataOut_payload_0_12059 : _zz_dataOut_payload_0_11963);
  assign _zz_dataOut_payload_0_12966 = (_zz_dataOut_payload_0_12964 ? _zz_dataOut_payload_0_11963 : _zz_dataOut_payload_0_12059);
  assign _zz_dataOut_payload_0_12967 = (_zz_dataOut_payload_0_12056 < _zz_dataOut_payload_0_11960);
  assign _zz_dataOut_payload_0_12968 = (_zz_dataOut_payload_0_12967 ? _zz_dataOut_payload_0_12056 : _zz_dataOut_payload_0_11960);
  assign _zz_dataOut_payload_0_12969 = (_zz_dataOut_payload_0_12967 ? _zz_dataOut_payload_0_11960 : _zz_dataOut_payload_0_12056);
  assign _zz_dataOut_payload_0_12970 = (_zz_dataOut_payload_0_12053 < _zz_dataOut_payload_0_11957);
  assign _zz_dataOut_payload_0_12971 = (_zz_dataOut_payload_0_12970 ? _zz_dataOut_payload_0_12053 : _zz_dataOut_payload_0_11957);
  assign _zz_dataOut_payload_0_12972 = (_zz_dataOut_payload_0_12970 ? _zz_dataOut_payload_0_11957 : _zz_dataOut_payload_0_12053);
  assign _zz_dataOut_payload_0_12973 = (_zz_dataOut_payload_0_12050 < _zz_dataOut_payload_0_11954);
  assign _zz_dataOut_payload_0_12974 = (_zz_dataOut_payload_0_12973 ? _zz_dataOut_payload_0_12050 : _zz_dataOut_payload_0_11954);
  assign _zz_dataOut_payload_0_12975 = (_zz_dataOut_payload_0_12973 ? _zz_dataOut_payload_0_11954 : _zz_dataOut_payload_0_12050);
  assign _zz_dataOut_payload_0_12976 = (_zz_dataOut_payload_0_12047 < _zz_dataOut_payload_0_11951);
  assign _zz_dataOut_payload_0_12977 = (_zz_dataOut_payload_0_12976 ? _zz_dataOut_payload_0_12047 : _zz_dataOut_payload_0_11951);
  assign _zz_dataOut_payload_0_12978 = (_zz_dataOut_payload_0_12976 ? _zz_dataOut_payload_0_11951 : _zz_dataOut_payload_0_12047);
  assign _zz_dataOut_payload_0_12979 = (_zz_dataOut_payload_0_12044 < _zz_dataOut_payload_0_11948);
  assign _zz_dataOut_payload_0_12980 = (_zz_dataOut_payload_0_12979 ? _zz_dataOut_payload_0_12044 : _zz_dataOut_payload_0_11948);
  assign _zz_dataOut_payload_0_12981 = (_zz_dataOut_payload_0_12979 ? _zz_dataOut_payload_0_11948 : _zz_dataOut_payload_0_12044);
  assign _zz_dataOut_payload_0_12982 = (_zz_dataOut_payload_0_12041 < _zz_dataOut_payload_0_11945);
  assign _zz_dataOut_payload_0_12983 = (_zz_dataOut_payload_0_12982 ? _zz_dataOut_payload_0_12041 : _zz_dataOut_payload_0_11945);
  assign _zz_dataOut_payload_0_12984 = (_zz_dataOut_payload_0_12982 ? _zz_dataOut_payload_0_11945 : _zz_dataOut_payload_0_12041);
  assign _zz_dataOut_payload_0_12985 = (_zz_dataOut_payload_0_12038 < _zz_dataOut_payload_0_11942);
  assign _zz_dataOut_payload_0_12986 = (_zz_dataOut_payload_0_12985 ? _zz_dataOut_payload_0_12038 : _zz_dataOut_payload_0_11942);
  assign _zz_dataOut_payload_0_12987 = (_zz_dataOut_payload_0_12985 ? _zz_dataOut_payload_0_11942 : _zz_dataOut_payload_0_12038);
  assign _zz_dataOut_payload_0_12988 = (_zz_dataOut_payload_0_12035 < _zz_dataOut_payload_0_11939);
  assign _zz_dataOut_payload_0_12989 = (_zz_dataOut_payload_0_12988 ? _zz_dataOut_payload_0_12035 : _zz_dataOut_payload_0_11939);
  assign _zz_dataOut_payload_0_12990 = (_zz_dataOut_payload_0_12988 ? _zz_dataOut_payload_0_11939 : _zz_dataOut_payload_0_12035);
  assign _zz_dataOut_payload_0_12991 = (_zz_dataOut_payload_0_12032 < _zz_dataOut_payload_0_11936);
  assign _zz_dataOut_payload_0_12992 = (_zz_dataOut_payload_0_12991 ? _zz_dataOut_payload_0_12032 : _zz_dataOut_payload_0_11936);
  assign _zz_dataOut_payload_0_12993 = (_zz_dataOut_payload_0_12991 ? _zz_dataOut_payload_0_11936 : _zz_dataOut_payload_0_12032);
  assign _zz_dataOut_payload_0_12994 = (_zz_dataOut_payload_0_12029 < _zz_dataOut_payload_0_11933);
  assign _zz_dataOut_payload_0_12995 = (_zz_dataOut_payload_0_12994 ? _zz_dataOut_payload_0_12029 : _zz_dataOut_payload_0_11933);
  assign _zz_dataOut_payload_0_12996 = (_zz_dataOut_payload_0_12994 ? _zz_dataOut_payload_0_11933 : _zz_dataOut_payload_0_12029);
  assign _zz_dataOut_payload_0_12997 = (_zz_dataOut_payload_0_12026 < _zz_dataOut_payload_0_11930);
  assign _zz_dataOut_payload_0_12998 = (_zz_dataOut_payload_0_12997 ? _zz_dataOut_payload_0_12026 : _zz_dataOut_payload_0_11930);
  assign _zz_dataOut_payload_0_12999 = (_zz_dataOut_payload_0_12997 ? _zz_dataOut_payload_0_11930 : _zz_dataOut_payload_0_12026);
  assign _zz_dataOut_payload_0_13000 = (_zz_dataOut_payload_0_12023 < _zz_dataOut_payload_0_11927);
  assign _zz_dataOut_payload_0_13001 = (_zz_dataOut_payload_0_13000 ? _zz_dataOut_payload_0_12023 : _zz_dataOut_payload_0_11927);
  assign _zz_dataOut_payload_0_13002 = (_zz_dataOut_payload_0_13000 ? _zz_dataOut_payload_0_11927 : _zz_dataOut_payload_0_12023);
  assign _zz_dataOut_payload_0_13003 = (_zz_dataOut_payload_0_12020 < _zz_dataOut_payload_0_11924);
  assign _zz_dataOut_payload_0_13004 = (_zz_dataOut_payload_0_13003 ? _zz_dataOut_payload_0_12020 : _zz_dataOut_payload_0_11924);
  assign _zz_dataOut_payload_0_13005 = (_zz_dataOut_payload_0_13003 ? _zz_dataOut_payload_0_11924 : _zz_dataOut_payload_0_12020);
  assign _zz_dataOut_payload_0_13006 = (_zz_dataOut_payload_0_12017 < _zz_dataOut_payload_0_11921);
  assign _zz_dataOut_payload_0_13007 = (_zz_dataOut_payload_0_13006 ? _zz_dataOut_payload_0_12017 : _zz_dataOut_payload_0_11921);
  assign _zz_dataOut_payload_0_13008 = (_zz_dataOut_payload_0_13006 ? _zz_dataOut_payload_0_11921 : _zz_dataOut_payload_0_12017);
  assign _zz_dataOut_payload_0_13009 = (_zz_dataOut_payload_0_12014 < _zz_dataOut_payload_0_11918);
  assign _zz_dataOut_payload_0_13010 = (_zz_dataOut_payload_0_13009 ? _zz_dataOut_payload_0_12014 : _zz_dataOut_payload_0_11918);
  assign _zz_dataOut_payload_0_13011 = (_zz_dataOut_payload_0_13009 ? _zz_dataOut_payload_0_11918 : _zz_dataOut_payload_0_12014);
  assign _zz_dataOut_payload_0_13012 = (_zz_dataOut_payload_0_12011 < _zz_dataOut_payload_0_11915);
  assign _zz_dataOut_payload_0_13013 = (_zz_dataOut_payload_0_13012 ? _zz_dataOut_payload_0_12011 : _zz_dataOut_payload_0_11915);
  assign _zz_dataOut_payload_0_13014 = (_zz_dataOut_payload_0_13012 ? _zz_dataOut_payload_0_11915 : _zz_dataOut_payload_0_12011);
  assign _zz_dataOut_payload_0_13015 = (_zz_dataOut_payload_0_12008 < _zz_dataOut_payload_0_11912);
  assign _zz_dataOut_payload_0_13016 = (_zz_dataOut_payload_0_13015 ? _zz_dataOut_payload_0_12008 : _zz_dataOut_payload_0_11912);
  assign _zz_dataOut_payload_0_13017 = (_zz_dataOut_payload_0_13015 ? _zz_dataOut_payload_0_11912 : _zz_dataOut_payload_0_12008);
  assign _zz_dataOut_payload_0_13018 = (_zz_dataOut_payload_0_12005 < _zz_dataOut_payload_0_11909);
  assign _zz_dataOut_payload_0_13019 = (_zz_dataOut_payload_0_13018 ? _zz_dataOut_payload_0_12005 : _zz_dataOut_payload_0_11909);
  assign _zz_dataOut_payload_0_13020 = (_zz_dataOut_payload_0_13018 ? _zz_dataOut_payload_0_11909 : _zz_dataOut_payload_0_12005);
  assign _zz_dataOut_payload_0_13021 = (_zz_dataOut_payload_0_12002 < _zz_dataOut_payload_0_11906);
  assign _zz_dataOut_payload_0_13022 = (_zz_dataOut_payload_0_13021 ? _zz_dataOut_payload_0_12002 : _zz_dataOut_payload_0_11906);
  assign _zz_dataOut_payload_0_13023 = (_zz_dataOut_payload_0_13021 ? _zz_dataOut_payload_0_11906 : _zz_dataOut_payload_0_12002);
  assign _zz_dataOut_payload_0_13024 = (_zz_dataOut_payload_0_12929 < _zz_dataOut_payload_0_12977);
  assign _zz_dataOut_payload_0_13025 = (_zz_dataOut_payload_0_13024 ? _zz_dataOut_payload_0_12929 : _zz_dataOut_payload_0_12977);
  assign _zz_dataOut_payload_0_13026 = (_zz_dataOut_payload_0_13024 ? _zz_dataOut_payload_0_12977 : _zz_dataOut_payload_0_12929);
  assign _zz_dataOut_payload_0_13027 = (_zz_dataOut_payload_0_12932 < _zz_dataOut_payload_0_12980);
  assign _zz_dataOut_payload_0_13028 = (_zz_dataOut_payload_0_13027 ? _zz_dataOut_payload_0_12932 : _zz_dataOut_payload_0_12980);
  assign _zz_dataOut_payload_0_13029 = (_zz_dataOut_payload_0_13027 ? _zz_dataOut_payload_0_12980 : _zz_dataOut_payload_0_12932);
  assign _zz_dataOut_payload_0_13030 = (_zz_dataOut_payload_0_12935 < _zz_dataOut_payload_0_12983);
  assign _zz_dataOut_payload_0_13031 = (_zz_dataOut_payload_0_13030 ? _zz_dataOut_payload_0_12935 : _zz_dataOut_payload_0_12983);
  assign _zz_dataOut_payload_0_13032 = (_zz_dataOut_payload_0_13030 ? _zz_dataOut_payload_0_12983 : _zz_dataOut_payload_0_12935);
  assign _zz_dataOut_payload_0_13033 = (_zz_dataOut_payload_0_12938 < _zz_dataOut_payload_0_12986);
  assign _zz_dataOut_payload_0_13034 = (_zz_dataOut_payload_0_13033 ? _zz_dataOut_payload_0_12938 : _zz_dataOut_payload_0_12986);
  assign _zz_dataOut_payload_0_13035 = (_zz_dataOut_payload_0_13033 ? _zz_dataOut_payload_0_12986 : _zz_dataOut_payload_0_12938);
  assign _zz_dataOut_payload_0_13036 = (_zz_dataOut_payload_0_12941 < _zz_dataOut_payload_0_12989);
  assign _zz_dataOut_payload_0_13037 = (_zz_dataOut_payload_0_13036 ? _zz_dataOut_payload_0_12941 : _zz_dataOut_payload_0_12989);
  assign _zz_dataOut_payload_0_13038 = (_zz_dataOut_payload_0_13036 ? _zz_dataOut_payload_0_12989 : _zz_dataOut_payload_0_12941);
  assign _zz_dataOut_payload_0_13039 = (_zz_dataOut_payload_0_12944 < _zz_dataOut_payload_0_12992);
  assign _zz_dataOut_payload_0_13040 = (_zz_dataOut_payload_0_13039 ? _zz_dataOut_payload_0_12944 : _zz_dataOut_payload_0_12992);
  assign _zz_dataOut_payload_0_13041 = (_zz_dataOut_payload_0_13039 ? _zz_dataOut_payload_0_12992 : _zz_dataOut_payload_0_12944);
  assign _zz_dataOut_payload_0_13042 = (_zz_dataOut_payload_0_12947 < _zz_dataOut_payload_0_12995);
  assign _zz_dataOut_payload_0_13043 = (_zz_dataOut_payload_0_13042 ? _zz_dataOut_payload_0_12947 : _zz_dataOut_payload_0_12995);
  assign _zz_dataOut_payload_0_13044 = (_zz_dataOut_payload_0_13042 ? _zz_dataOut_payload_0_12995 : _zz_dataOut_payload_0_12947);
  assign _zz_dataOut_payload_0_13045 = (_zz_dataOut_payload_0_12950 < _zz_dataOut_payload_0_12998);
  assign _zz_dataOut_payload_0_13046 = (_zz_dataOut_payload_0_13045 ? _zz_dataOut_payload_0_12950 : _zz_dataOut_payload_0_12998);
  assign _zz_dataOut_payload_0_13047 = (_zz_dataOut_payload_0_13045 ? _zz_dataOut_payload_0_12998 : _zz_dataOut_payload_0_12950);
  assign _zz_dataOut_payload_0_13048 = (_zz_dataOut_payload_0_12953 < _zz_dataOut_payload_0_13001);
  assign _zz_dataOut_payload_0_13049 = (_zz_dataOut_payload_0_13048 ? _zz_dataOut_payload_0_12953 : _zz_dataOut_payload_0_13001);
  assign _zz_dataOut_payload_0_13050 = (_zz_dataOut_payload_0_13048 ? _zz_dataOut_payload_0_13001 : _zz_dataOut_payload_0_12953);
  assign _zz_dataOut_payload_0_13051 = (_zz_dataOut_payload_0_12956 < _zz_dataOut_payload_0_13004);
  assign _zz_dataOut_payload_0_13052 = (_zz_dataOut_payload_0_13051 ? _zz_dataOut_payload_0_12956 : _zz_dataOut_payload_0_13004);
  assign _zz_dataOut_payload_0_13053 = (_zz_dataOut_payload_0_13051 ? _zz_dataOut_payload_0_13004 : _zz_dataOut_payload_0_12956);
  assign _zz_dataOut_payload_0_13054 = (_zz_dataOut_payload_0_12959 < _zz_dataOut_payload_0_13007);
  assign _zz_dataOut_payload_0_13055 = (_zz_dataOut_payload_0_13054 ? _zz_dataOut_payload_0_12959 : _zz_dataOut_payload_0_13007);
  assign _zz_dataOut_payload_0_13056 = (_zz_dataOut_payload_0_13054 ? _zz_dataOut_payload_0_13007 : _zz_dataOut_payload_0_12959);
  assign _zz_dataOut_payload_0_13057 = (_zz_dataOut_payload_0_12962 < _zz_dataOut_payload_0_13010);
  assign _zz_dataOut_payload_0_13058 = (_zz_dataOut_payload_0_13057 ? _zz_dataOut_payload_0_12962 : _zz_dataOut_payload_0_13010);
  assign _zz_dataOut_payload_0_13059 = (_zz_dataOut_payload_0_13057 ? _zz_dataOut_payload_0_13010 : _zz_dataOut_payload_0_12962);
  assign _zz_dataOut_payload_0_13060 = (_zz_dataOut_payload_0_12965 < _zz_dataOut_payload_0_13013);
  assign _zz_dataOut_payload_0_13061 = (_zz_dataOut_payload_0_13060 ? _zz_dataOut_payload_0_12965 : _zz_dataOut_payload_0_13013);
  assign _zz_dataOut_payload_0_13062 = (_zz_dataOut_payload_0_13060 ? _zz_dataOut_payload_0_13013 : _zz_dataOut_payload_0_12965);
  assign _zz_dataOut_payload_0_13063 = (_zz_dataOut_payload_0_12968 < _zz_dataOut_payload_0_13016);
  assign _zz_dataOut_payload_0_13064 = (_zz_dataOut_payload_0_13063 ? _zz_dataOut_payload_0_12968 : _zz_dataOut_payload_0_13016);
  assign _zz_dataOut_payload_0_13065 = (_zz_dataOut_payload_0_13063 ? _zz_dataOut_payload_0_13016 : _zz_dataOut_payload_0_12968);
  assign _zz_dataOut_payload_0_13066 = (_zz_dataOut_payload_0_12971 < _zz_dataOut_payload_0_13019);
  assign _zz_dataOut_payload_0_13067 = (_zz_dataOut_payload_0_13066 ? _zz_dataOut_payload_0_12971 : _zz_dataOut_payload_0_13019);
  assign _zz_dataOut_payload_0_13068 = (_zz_dataOut_payload_0_13066 ? _zz_dataOut_payload_0_13019 : _zz_dataOut_payload_0_12971);
  assign _zz_dataOut_payload_0_13069 = (_zz_dataOut_payload_0_12974 < _zz_dataOut_payload_0_13022);
  assign _zz_dataOut_payload_0_13070 = (_zz_dataOut_payload_0_13069 ? _zz_dataOut_payload_0_12974 : _zz_dataOut_payload_0_13022);
  assign _zz_dataOut_payload_0_13071 = (_zz_dataOut_payload_0_13069 ? _zz_dataOut_payload_0_13022 : _zz_dataOut_payload_0_12974);
  assign _zz_dataOut_payload_0_13072 = (_zz_dataOut_payload_0_13025 < _zz_dataOut_payload_0_13049);
  assign _zz_dataOut_payload_0_13073 = (_zz_dataOut_payload_0_13072 ? _zz_dataOut_payload_0_13025 : _zz_dataOut_payload_0_13049);
  assign _zz_dataOut_payload_0_13074 = (_zz_dataOut_payload_0_13072 ? _zz_dataOut_payload_0_13049 : _zz_dataOut_payload_0_13025);
  assign _zz_dataOut_payload_0_13075 = (_zz_dataOut_payload_0_13028 < _zz_dataOut_payload_0_13052);
  assign _zz_dataOut_payload_0_13076 = (_zz_dataOut_payload_0_13075 ? _zz_dataOut_payload_0_13028 : _zz_dataOut_payload_0_13052);
  assign _zz_dataOut_payload_0_13077 = (_zz_dataOut_payload_0_13075 ? _zz_dataOut_payload_0_13052 : _zz_dataOut_payload_0_13028);
  assign _zz_dataOut_payload_0_13078 = (_zz_dataOut_payload_0_13031 < _zz_dataOut_payload_0_13055);
  assign _zz_dataOut_payload_0_13079 = (_zz_dataOut_payload_0_13078 ? _zz_dataOut_payload_0_13031 : _zz_dataOut_payload_0_13055);
  assign _zz_dataOut_payload_0_13080 = (_zz_dataOut_payload_0_13078 ? _zz_dataOut_payload_0_13055 : _zz_dataOut_payload_0_13031);
  assign _zz_dataOut_payload_0_13081 = (_zz_dataOut_payload_0_13034 < _zz_dataOut_payload_0_13058);
  assign _zz_dataOut_payload_0_13082 = (_zz_dataOut_payload_0_13081 ? _zz_dataOut_payload_0_13034 : _zz_dataOut_payload_0_13058);
  assign _zz_dataOut_payload_0_13083 = (_zz_dataOut_payload_0_13081 ? _zz_dataOut_payload_0_13058 : _zz_dataOut_payload_0_13034);
  assign _zz_dataOut_payload_0_13084 = (_zz_dataOut_payload_0_13037 < _zz_dataOut_payload_0_13061);
  assign _zz_dataOut_payload_0_13085 = (_zz_dataOut_payload_0_13084 ? _zz_dataOut_payload_0_13037 : _zz_dataOut_payload_0_13061);
  assign _zz_dataOut_payload_0_13086 = (_zz_dataOut_payload_0_13084 ? _zz_dataOut_payload_0_13061 : _zz_dataOut_payload_0_13037);
  assign _zz_dataOut_payload_0_13087 = (_zz_dataOut_payload_0_13040 < _zz_dataOut_payload_0_13064);
  assign _zz_dataOut_payload_0_13088 = (_zz_dataOut_payload_0_13087 ? _zz_dataOut_payload_0_13040 : _zz_dataOut_payload_0_13064);
  assign _zz_dataOut_payload_0_13089 = (_zz_dataOut_payload_0_13087 ? _zz_dataOut_payload_0_13064 : _zz_dataOut_payload_0_13040);
  assign _zz_dataOut_payload_0_13090 = (_zz_dataOut_payload_0_13043 < _zz_dataOut_payload_0_13067);
  assign _zz_dataOut_payload_0_13091 = (_zz_dataOut_payload_0_13090 ? _zz_dataOut_payload_0_13043 : _zz_dataOut_payload_0_13067);
  assign _zz_dataOut_payload_0_13092 = (_zz_dataOut_payload_0_13090 ? _zz_dataOut_payload_0_13067 : _zz_dataOut_payload_0_13043);
  assign _zz_dataOut_payload_0_13093 = (_zz_dataOut_payload_0_13046 < _zz_dataOut_payload_0_13070);
  assign _zz_dataOut_payload_0_13094 = (_zz_dataOut_payload_0_13093 ? _zz_dataOut_payload_0_13046 : _zz_dataOut_payload_0_13070);
  assign _zz_dataOut_payload_0_13095 = (_zz_dataOut_payload_0_13093 ? _zz_dataOut_payload_0_13070 : _zz_dataOut_payload_0_13046);
  assign _zz_dataOut_payload_0_13096 = (_zz_dataOut_payload_0_13073 < _zz_dataOut_payload_0_13085);
  assign _zz_dataOut_payload_0_13097 = (_zz_dataOut_payload_0_13096 ? _zz_dataOut_payload_0_13073 : _zz_dataOut_payload_0_13085);
  assign _zz_dataOut_payload_0_13098 = (_zz_dataOut_payload_0_13096 ? _zz_dataOut_payload_0_13085 : _zz_dataOut_payload_0_13073);
  assign _zz_dataOut_payload_0_13099 = (_zz_dataOut_payload_0_13076 < _zz_dataOut_payload_0_13088);
  assign _zz_dataOut_payload_0_13100 = (_zz_dataOut_payload_0_13099 ? _zz_dataOut_payload_0_13076 : _zz_dataOut_payload_0_13088);
  assign _zz_dataOut_payload_0_13101 = (_zz_dataOut_payload_0_13099 ? _zz_dataOut_payload_0_13088 : _zz_dataOut_payload_0_13076);
  assign _zz_dataOut_payload_0_13102 = (_zz_dataOut_payload_0_13079 < _zz_dataOut_payload_0_13091);
  assign _zz_dataOut_payload_0_13103 = (_zz_dataOut_payload_0_13102 ? _zz_dataOut_payload_0_13079 : _zz_dataOut_payload_0_13091);
  assign _zz_dataOut_payload_0_13104 = (_zz_dataOut_payload_0_13102 ? _zz_dataOut_payload_0_13091 : _zz_dataOut_payload_0_13079);
  assign _zz_dataOut_payload_0_13105 = (_zz_dataOut_payload_0_13082 < _zz_dataOut_payload_0_13094);
  assign _zz_dataOut_payload_0_13106 = (_zz_dataOut_payload_0_13105 ? _zz_dataOut_payload_0_13082 : _zz_dataOut_payload_0_13094);
  assign _zz_dataOut_payload_0_13107 = (_zz_dataOut_payload_0_13105 ? _zz_dataOut_payload_0_13094 : _zz_dataOut_payload_0_13082);
  assign _zz_dataOut_payload_0_13108 = (_zz_dataOut_payload_0_13097 < _zz_dataOut_payload_0_13103);
  assign _zz_dataOut_payload_0_13109 = (_zz_dataOut_payload_0_13108 ? _zz_dataOut_payload_0_13097 : _zz_dataOut_payload_0_13103);
  assign _zz_dataOut_payload_0_13110 = (_zz_dataOut_payload_0_13108 ? _zz_dataOut_payload_0_13103 : _zz_dataOut_payload_0_13097);
  assign _zz_dataOut_payload_0_13111 = (_zz_dataOut_payload_0_13100 < _zz_dataOut_payload_0_13106);
  assign _zz_dataOut_payload_0_13112 = (_zz_dataOut_payload_0_13111 ? _zz_dataOut_payload_0_13100 : _zz_dataOut_payload_0_13106);
  assign _zz_dataOut_payload_0_13113 = (_zz_dataOut_payload_0_13111 ? _zz_dataOut_payload_0_13106 : _zz_dataOut_payload_0_13100);
  assign _zz_dataOut_payload_0_13114 = (_zz_dataOut_payload_0_13109 < _zz_dataOut_payload_0_13112);
  assign _zz_dataOut_payload_0_13115 = (_zz_dataOut_payload_0_13110 < _zz_dataOut_payload_0_13113);
  assign _zz_dataOut_payload_0_13120 = (_zz_dataOut_payload_0_13098 < _zz_dataOut_payload_0_13104);
  assign _zz_dataOut_payload_0_13121 = (_zz_dataOut_payload_0_13120 ? _zz_dataOut_payload_0_13098 : _zz_dataOut_payload_0_13104);
  assign _zz_dataOut_payload_0_13122 = (_zz_dataOut_payload_0_13120 ? _zz_dataOut_payload_0_13104 : _zz_dataOut_payload_0_13098);
  assign _zz_dataOut_payload_0_13123 = (_zz_dataOut_payload_0_13101 < _zz_dataOut_payload_0_13107);
  assign _zz_dataOut_payload_0_13124 = (_zz_dataOut_payload_0_13123 ? _zz_dataOut_payload_0_13101 : _zz_dataOut_payload_0_13107);
  assign _zz_dataOut_payload_0_13125 = (_zz_dataOut_payload_0_13123 ? _zz_dataOut_payload_0_13107 : _zz_dataOut_payload_0_13101);
  assign _zz_dataOut_payload_0_13126 = (_zz_dataOut_payload_0_13121 < _zz_dataOut_payload_0_13124);
  assign _zz_dataOut_payload_0_13127 = (_zz_dataOut_payload_0_13122 < _zz_dataOut_payload_0_13125);
  assign _zz_dataOut_payload_0_13140 = (_zz_dataOut_payload_0_13074 < _zz_dataOut_payload_0_13086);
  assign _zz_dataOut_payload_0_13141 = (_zz_dataOut_payload_0_13140 ? _zz_dataOut_payload_0_13074 : _zz_dataOut_payload_0_13086);
  assign _zz_dataOut_payload_0_13142 = (_zz_dataOut_payload_0_13140 ? _zz_dataOut_payload_0_13086 : _zz_dataOut_payload_0_13074);
  assign _zz_dataOut_payload_0_13143 = (_zz_dataOut_payload_0_13077 < _zz_dataOut_payload_0_13089);
  assign _zz_dataOut_payload_0_13144 = (_zz_dataOut_payload_0_13143 ? _zz_dataOut_payload_0_13077 : _zz_dataOut_payload_0_13089);
  assign _zz_dataOut_payload_0_13145 = (_zz_dataOut_payload_0_13143 ? _zz_dataOut_payload_0_13089 : _zz_dataOut_payload_0_13077);
  assign _zz_dataOut_payload_0_13146 = (_zz_dataOut_payload_0_13080 < _zz_dataOut_payload_0_13092);
  assign _zz_dataOut_payload_0_13147 = (_zz_dataOut_payload_0_13146 ? _zz_dataOut_payload_0_13080 : _zz_dataOut_payload_0_13092);
  assign _zz_dataOut_payload_0_13148 = (_zz_dataOut_payload_0_13146 ? _zz_dataOut_payload_0_13092 : _zz_dataOut_payload_0_13080);
  assign _zz_dataOut_payload_0_13149 = (_zz_dataOut_payload_0_13083 < _zz_dataOut_payload_0_13095);
  assign _zz_dataOut_payload_0_13150 = (_zz_dataOut_payload_0_13149 ? _zz_dataOut_payload_0_13083 : _zz_dataOut_payload_0_13095);
  assign _zz_dataOut_payload_0_13151 = (_zz_dataOut_payload_0_13149 ? _zz_dataOut_payload_0_13095 : _zz_dataOut_payload_0_13083);
  assign _zz_dataOut_payload_0_13152 = (_zz_dataOut_payload_0_13141 < _zz_dataOut_payload_0_13147);
  assign _zz_dataOut_payload_0_13153 = (_zz_dataOut_payload_0_13152 ? _zz_dataOut_payload_0_13141 : _zz_dataOut_payload_0_13147);
  assign _zz_dataOut_payload_0_13154 = (_zz_dataOut_payload_0_13152 ? _zz_dataOut_payload_0_13147 : _zz_dataOut_payload_0_13141);
  assign _zz_dataOut_payload_0_13155 = (_zz_dataOut_payload_0_13144 < _zz_dataOut_payload_0_13150);
  assign _zz_dataOut_payload_0_13156 = (_zz_dataOut_payload_0_13155 ? _zz_dataOut_payload_0_13144 : _zz_dataOut_payload_0_13150);
  assign _zz_dataOut_payload_0_13157 = (_zz_dataOut_payload_0_13155 ? _zz_dataOut_payload_0_13150 : _zz_dataOut_payload_0_13144);
  assign _zz_dataOut_payload_0_13158 = (_zz_dataOut_payload_0_13153 < _zz_dataOut_payload_0_13156);
  assign _zz_dataOut_payload_0_13159 = (_zz_dataOut_payload_0_13154 < _zz_dataOut_payload_0_13157);
  assign _zz_dataOut_payload_0_13164 = (_zz_dataOut_payload_0_13142 < _zz_dataOut_payload_0_13148);
  assign _zz_dataOut_payload_0_13165 = (_zz_dataOut_payload_0_13164 ? _zz_dataOut_payload_0_13142 : _zz_dataOut_payload_0_13148);
  assign _zz_dataOut_payload_0_13166 = (_zz_dataOut_payload_0_13164 ? _zz_dataOut_payload_0_13148 : _zz_dataOut_payload_0_13142);
  assign _zz_dataOut_payload_0_13167 = (_zz_dataOut_payload_0_13145 < _zz_dataOut_payload_0_13151);
  assign _zz_dataOut_payload_0_13168 = (_zz_dataOut_payload_0_13167 ? _zz_dataOut_payload_0_13145 : _zz_dataOut_payload_0_13151);
  assign _zz_dataOut_payload_0_13169 = (_zz_dataOut_payload_0_13167 ? _zz_dataOut_payload_0_13151 : _zz_dataOut_payload_0_13145);
  assign _zz_dataOut_payload_0_13170 = (_zz_dataOut_payload_0_13165 < _zz_dataOut_payload_0_13168);
  assign _zz_dataOut_payload_0_13171 = (_zz_dataOut_payload_0_13166 < _zz_dataOut_payload_0_13169);
  assign _zz_dataOut_payload_0_13200 = (_zz_dataOut_payload_0_13026 < _zz_dataOut_payload_0_13050);
  assign _zz_dataOut_payload_0_13201 = (_zz_dataOut_payload_0_13200 ? _zz_dataOut_payload_0_13026 : _zz_dataOut_payload_0_13050);
  assign _zz_dataOut_payload_0_13202 = (_zz_dataOut_payload_0_13200 ? _zz_dataOut_payload_0_13050 : _zz_dataOut_payload_0_13026);
  assign _zz_dataOut_payload_0_13203 = (_zz_dataOut_payload_0_13029 < _zz_dataOut_payload_0_13053);
  assign _zz_dataOut_payload_0_13204 = (_zz_dataOut_payload_0_13203 ? _zz_dataOut_payload_0_13029 : _zz_dataOut_payload_0_13053);
  assign _zz_dataOut_payload_0_13205 = (_zz_dataOut_payload_0_13203 ? _zz_dataOut_payload_0_13053 : _zz_dataOut_payload_0_13029);
  assign _zz_dataOut_payload_0_13206 = (_zz_dataOut_payload_0_13032 < _zz_dataOut_payload_0_13056);
  assign _zz_dataOut_payload_0_13207 = (_zz_dataOut_payload_0_13206 ? _zz_dataOut_payload_0_13032 : _zz_dataOut_payload_0_13056);
  assign _zz_dataOut_payload_0_13208 = (_zz_dataOut_payload_0_13206 ? _zz_dataOut_payload_0_13056 : _zz_dataOut_payload_0_13032);
  assign _zz_dataOut_payload_0_13209 = (_zz_dataOut_payload_0_13035 < _zz_dataOut_payload_0_13059);
  assign _zz_dataOut_payload_0_13210 = (_zz_dataOut_payload_0_13209 ? _zz_dataOut_payload_0_13035 : _zz_dataOut_payload_0_13059);
  assign _zz_dataOut_payload_0_13211 = (_zz_dataOut_payload_0_13209 ? _zz_dataOut_payload_0_13059 : _zz_dataOut_payload_0_13035);
  assign _zz_dataOut_payload_0_13212 = (_zz_dataOut_payload_0_13038 < _zz_dataOut_payload_0_13062);
  assign _zz_dataOut_payload_0_13213 = (_zz_dataOut_payload_0_13212 ? _zz_dataOut_payload_0_13038 : _zz_dataOut_payload_0_13062);
  assign _zz_dataOut_payload_0_13214 = (_zz_dataOut_payload_0_13212 ? _zz_dataOut_payload_0_13062 : _zz_dataOut_payload_0_13038);
  assign _zz_dataOut_payload_0_13215 = (_zz_dataOut_payload_0_13041 < _zz_dataOut_payload_0_13065);
  assign _zz_dataOut_payload_0_13216 = (_zz_dataOut_payload_0_13215 ? _zz_dataOut_payload_0_13041 : _zz_dataOut_payload_0_13065);
  assign _zz_dataOut_payload_0_13217 = (_zz_dataOut_payload_0_13215 ? _zz_dataOut_payload_0_13065 : _zz_dataOut_payload_0_13041);
  assign _zz_dataOut_payload_0_13218 = (_zz_dataOut_payload_0_13044 < _zz_dataOut_payload_0_13068);
  assign _zz_dataOut_payload_0_13219 = (_zz_dataOut_payload_0_13218 ? _zz_dataOut_payload_0_13044 : _zz_dataOut_payload_0_13068);
  assign _zz_dataOut_payload_0_13220 = (_zz_dataOut_payload_0_13218 ? _zz_dataOut_payload_0_13068 : _zz_dataOut_payload_0_13044);
  assign _zz_dataOut_payload_0_13221 = (_zz_dataOut_payload_0_13047 < _zz_dataOut_payload_0_13071);
  assign _zz_dataOut_payload_0_13222 = (_zz_dataOut_payload_0_13221 ? _zz_dataOut_payload_0_13047 : _zz_dataOut_payload_0_13071);
  assign _zz_dataOut_payload_0_13223 = (_zz_dataOut_payload_0_13221 ? _zz_dataOut_payload_0_13071 : _zz_dataOut_payload_0_13047);
  assign _zz_dataOut_payload_0_13224 = (_zz_dataOut_payload_0_13201 < _zz_dataOut_payload_0_13213);
  assign _zz_dataOut_payload_0_13225 = (_zz_dataOut_payload_0_13224 ? _zz_dataOut_payload_0_13201 : _zz_dataOut_payload_0_13213);
  assign _zz_dataOut_payload_0_13226 = (_zz_dataOut_payload_0_13224 ? _zz_dataOut_payload_0_13213 : _zz_dataOut_payload_0_13201);
  assign _zz_dataOut_payload_0_13227 = (_zz_dataOut_payload_0_13204 < _zz_dataOut_payload_0_13216);
  assign _zz_dataOut_payload_0_13228 = (_zz_dataOut_payload_0_13227 ? _zz_dataOut_payload_0_13204 : _zz_dataOut_payload_0_13216);
  assign _zz_dataOut_payload_0_13229 = (_zz_dataOut_payload_0_13227 ? _zz_dataOut_payload_0_13216 : _zz_dataOut_payload_0_13204);
  assign _zz_dataOut_payload_0_13230 = (_zz_dataOut_payload_0_13207 < _zz_dataOut_payload_0_13219);
  assign _zz_dataOut_payload_0_13231 = (_zz_dataOut_payload_0_13230 ? _zz_dataOut_payload_0_13207 : _zz_dataOut_payload_0_13219);
  assign _zz_dataOut_payload_0_13232 = (_zz_dataOut_payload_0_13230 ? _zz_dataOut_payload_0_13219 : _zz_dataOut_payload_0_13207);
  assign _zz_dataOut_payload_0_13233 = (_zz_dataOut_payload_0_13210 < _zz_dataOut_payload_0_13222);
  assign _zz_dataOut_payload_0_13234 = (_zz_dataOut_payload_0_13233 ? _zz_dataOut_payload_0_13210 : _zz_dataOut_payload_0_13222);
  assign _zz_dataOut_payload_0_13235 = (_zz_dataOut_payload_0_13233 ? _zz_dataOut_payload_0_13222 : _zz_dataOut_payload_0_13210);
  assign _zz_dataOut_payload_0_13236 = (_zz_dataOut_payload_0_13225 < _zz_dataOut_payload_0_13231);
  assign _zz_dataOut_payload_0_13237 = (_zz_dataOut_payload_0_13236 ? _zz_dataOut_payload_0_13225 : _zz_dataOut_payload_0_13231);
  assign _zz_dataOut_payload_0_13238 = (_zz_dataOut_payload_0_13236 ? _zz_dataOut_payload_0_13231 : _zz_dataOut_payload_0_13225);
  assign _zz_dataOut_payload_0_13239 = (_zz_dataOut_payload_0_13228 < _zz_dataOut_payload_0_13234);
  assign _zz_dataOut_payload_0_13240 = (_zz_dataOut_payload_0_13239 ? _zz_dataOut_payload_0_13228 : _zz_dataOut_payload_0_13234);
  assign _zz_dataOut_payload_0_13241 = (_zz_dataOut_payload_0_13239 ? _zz_dataOut_payload_0_13234 : _zz_dataOut_payload_0_13228);
  assign _zz_dataOut_payload_0_13242 = (_zz_dataOut_payload_0_13237 < _zz_dataOut_payload_0_13240);
  assign _zz_dataOut_payload_0_13243 = (_zz_dataOut_payload_0_13238 < _zz_dataOut_payload_0_13241);
  assign _zz_dataOut_payload_0_13248 = (_zz_dataOut_payload_0_13226 < _zz_dataOut_payload_0_13232);
  assign _zz_dataOut_payload_0_13249 = (_zz_dataOut_payload_0_13248 ? _zz_dataOut_payload_0_13226 : _zz_dataOut_payload_0_13232);
  assign _zz_dataOut_payload_0_13250 = (_zz_dataOut_payload_0_13248 ? _zz_dataOut_payload_0_13232 : _zz_dataOut_payload_0_13226);
  assign _zz_dataOut_payload_0_13251 = (_zz_dataOut_payload_0_13229 < _zz_dataOut_payload_0_13235);
  assign _zz_dataOut_payload_0_13252 = (_zz_dataOut_payload_0_13251 ? _zz_dataOut_payload_0_13229 : _zz_dataOut_payload_0_13235);
  assign _zz_dataOut_payload_0_13253 = (_zz_dataOut_payload_0_13251 ? _zz_dataOut_payload_0_13235 : _zz_dataOut_payload_0_13229);
  assign _zz_dataOut_payload_0_13254 = (_zz_dataOut_payload_0_13249 < _zz_dataOut_payload_0_13252);
  assign _zz_dataOut_payload_0_13255 = (_zz_dataOut_payload_0_13250 < _zz_dataOut_payload_0_13253);
  assign _zz_dataOut_payload_0_13268 = (_zz_dataOut_payload_0_13202 < _zz_dataOut_payload_0_13214);
  assign _zz_dataOut_payload_0_13269 = (_zz_dataOut_payload_0_13268 ? _zz_dataOut_payload_0_13202 : _zz_dataOut_payload_0_13214);
  assign _zz_dataOut_payload_0_13270 = (_zz_dataOut_payload_0_13268 ? _zz_dataOut_payload_0_13214 : _zz_dataOut_payload_0_13202);
  assign _zz_dataOut_payload_0_13271 = (_zz_dataOut_payload_0_13205 < _zz_dataOut_payload_0_13217);
  assign _zz_dataOut_payload_0_13272 = (_zz_dataOut_payload_0_13271 ? _zz_dataOut_payload_0_13205 : _zz_dataOut_payload_0_13217);
  assign _zz_dataOut_payload_0_13273 = (_zz_dataOut_payload_0_13271 ? _zz_dataOut_payload_0_13217 : _zz_dataOut_payload_0_13205);
  assign _zz_dataOut_payload_0_13274 = (_zz_dataOut_payload_0_13208 < _zz_dataOut_payload_0_13220);
  assign _zz_dataOut_payload_0_13275 = (_zz_dataOut_payload_0_13274 ? _zz_dataOut_payload_0_13208 : _zz_dataOut_payload_0_13220);
  assign _zz_dataOut_payload_0_13276 = (_zz_dataOut_payload_0_13274 ? _zz_dataOut_payload_0_13220 : _zz_dataOut_payload_0_13208);
  assign _zz_dataOut_payload_0_13277 = (_zz_dataOut_payload_0_13211 < _zz_dataOut_payload_0_13223);
  assign _zz_dataOut_payload_0_13278 = (_zz_dataOut_payload_0_13277 ? _zz_dataOut_payload_0_13211 : _zz_dataOut_payload_0_13223);
  assign _zz_dataOut_payload_0_13279 = (_zz_dataOut_payload_0_13277 ? _zz_dataOut_payload_0_13223 : _zz_dataOut_payload_0_13211);
  assign _zz_dataOut_payload_0_13280 = (_zz_dataOut_payload_0_13269 < _zz_dataOut_payload_0_13275);
  assign _zz_dataOut_payload_0_13281 = (_zz_dataOut_payload_0_13280 ? _zz_dataOut_payload_0_13269 : _zz_dataOut_payload_0_13275);
  assign _zz_dataOut_payload_0_13282 = (_zz_dataOut_payload_0_13280 ? _zz_dataOut_payload_0_13275 : _zz_dataOut_payload_0_13269);
  assign _zz_dataOut_payload_0_13283 = (_zz_dataOut_payload_0_13272 < _zz_dataOut_payload_0_13278);
  assign _zz_dataOut_payload_0_13284 = (_zz_dataOut_payload_0_13283 ? _zz_dataOut_payload_0_13272 : _zz_dataOut_payload_0_13278);
  assign _zz_dataOut_payload_0_13285 = (_zz_dataOut_payload_0_13283 ? _zz_dataOut_payload_0_13278 : _zz_dataOut_payload_0_13272);
  assign _zz_dataOut_payload_0_13286 = (_zz_dataOut_payload_0_13281 < _zz_dataOut_payload_0_13284);
  assign _zz_dataOut_payload_0_13287 = (_zz_dataOut_payload_0_13282 < _zz_dataOut_payload_0_13285);
  assign _zz_dataOut_payload_0_13292 = (_zz_dataOut_payload_0_13270 < _zz_dataOut_payload_0_13276);
  assign _zz_dataOut_payload_0_13293 = (_zz_dataOut_payload_0_13292 ? _zz_dataOut_payload_0_13270 : _zz_dataOut_payload_0_13276);
  assign _zz_dataOut_payload_0_13294 = (_zz_dataOut_payload_0_13292 ? _zz_dataOut_payload_0_13276 : _zz_dataOut_payload_0_13270);
  assign _zz_dataOut_payload_0_13295 = (_zz_dataOut_payload_0_13273 < _zz_dataOut_payload_0_13279);
  assign _zz_dataOut_payload_0_13296 = (_zz_dataOut_payload_0_13295 ? _zz_dataOut_payload_0_13273 : _zz_dataOut_payload_0_13279);
  assign _zz_dataOut_payload_0_13297 = (_zz_dataOut_payload_0_13295 ? _zz_dataOut_payload_0_13279 : _zz_dataOut_payload_0_13273);
  assign _zz_dataOut_payload_0_13298 = (_zz_dataOut_payload_0_13293 < _zz_dataOut_payload_0_13296);
  assign _zz_dataOut_payload_0_13299 = (_zz_dataOut_payload_0_13294 < _zz_dataOut_payload_0_13297);
  assign _zz_dataOut_payload_0_13360 = (_zz_dataOut_payload_0_12930 < _zz_dataOut_payload_0_12978);
  assign _zz_dataOut_payload_0_13361 = (_zz_dataOut_payload_0_13360 ? _zz_dataOut_payload_0_12930 : _zz_dataOut_payload_0_12978);
  assign _zz_dataOut_payload_0_13362 = (_zz_dataOut_payload_0_13360 ? _zz_dataOut_payload_0_12978 : _zz_dataOut_payload_0_12930);
  assign _zz_dataOut_payload_0_13363 = (_zz_dataOut_payload_0_12933 < _zz_dataOut_payload_0_12981);
  assign _zz_dataOut_payload_0_13364 = (_zz_dataOut_payload_0_13363 ? _zz_dataOut_payload_0_12933 : _zz_dataOut_payload_0_12981);
  assign _zz_dataOut_payload_0_13365 = (_zz_dataOut_payload_0_13363 ? _zz_dataOut_payload_0_12981 : _zz_dataOut_payload_0_12933);
  assign _zz_dataOut_payload_0_13366 = (_zz_dataOut_payload_0_12936 < _zz_dataOut_payload_0_12984);
  assign _zz_dataOut_payload_0_13367 = (_zz_dataOut_payload_0_13366 ? _zz_dataOut_payload_0_12936 : _zz_dataOut_payload_0_12984);
  assign _zz_dataOut_payload_0_13368 = (_zz_dataOut_payload_0_13366 ? _zz_dataOut_payload_0_12984 : _zz_dataOut_payload_0_12936);
  assign _zz_dataOut_payload_0_13369 = (_zz_dataOut_payload_0_12939 < _zz_dataOut_payload_0_12987);
  assign _zz_dataOut_payload_0_13370 = (_zz_dataOut_payload_0_13369 ? _zz_dataOut_payload_0_12939 : _zz_dataOut_payload_0_12987);
  assign _zz_dataOut_payload_0_13371 = (_zz_dataOut_payload_0_13369 ? _zz_dataOut_payload_0_12987 : _zz_dataOut_payload_0_12939);
  assign _zz_dataOut_payload_0_13372 = (_zz_dataOut_payload_0_12942 < _zz_dataOut_payload_0_12990);
  assign _zz_dataOut_payload_0_13373 = (_zz_dataOut_payload_0_13372 ? _zz_dataOut_payload_0_12942 : _zz_dataOut_payload_0_12990);
  assign _zz_dataOut_payload_0_13374 = (_zz_dataOut_payload_0_13372 ? _zz_dataOut_payload_0_12990 : _zz_dataOut_payload_0_12942);
  assign _zz_dataOut_payload_0_13375 = (_zz_dataOut_payload_0_12945 < _zz_dataOut_payload_0_12993);
  assign _zz_dataOut_payload_0_13376 = (_zz_dataOut_payload_0_13375 ? _zz_dataOut_payload_0_12945 : _zz_dataOut_payload_0_12993);
  assign _zz_dataOut_payload_0_13377 = (_zz_dataOut_payload_0_13375 ? _zz_dataOut_payload_0_12993 : _zz_dataOut_payload_0_12945);
  assign _zz_dataOut_payload_0_13378 = (_zz_dataOut_payload_0_12948 < _zz_dataOut_payload_0_12996);
  assign _zz_dataOut_payload_0_13379 = (_zz_dataOut_payload_0_13378 ? _zz_dataOut_payload_0_12948 : _zz_dataOut_payload_0_12996);
  assign _zz_dataOut_payload_0_13380 = (_zz_dataOut_payload_0_13378 ? _zz_dataOut_payload_0_12996 : _zz_dataOut_payload_0_12948);
  assign _zz_dataOut_payload_0_13381 = (_zz_dataOut_payload_0_12951 < _zz_dataOut_payload_0_12999);
  assign _zz_dataOut_payload_0_13382 = (_zz_dataOut_payload_0_13381 ? _zz_dataOut_payload_0_12951 : _zz_dataOut_payload_0_12999);
  assign _zz_dataOut_payload_0_13383 = (_zz_dataOut_payload_0_13381 ? _zz_dataOut_payload_0_12999 : _zz_dataOut_payload_0_12951);
  assign _zz_dataOut_payload_0_13384 = (_zz_dataOut_payload_0_12954 < _zz_dataOut_payload_0_13002);
  assign _zz_dataOut_payload_0_13385 = (_zz_dataOut_payload_0_13384 ? _zz_dataOut_payload_0_12954 : _zz_dataOut_payload_0_13002);
  assign _zz_dataOut_payload_0_13386 = (_zz_dataOut_payload_0_13384 ? _zz_dataOut_payload_0_13002 : _zz_dataOut_payload_0_12954);
  assign _zz_dataOut_payload_0_13387 = (_zz_dataOut_payload_0_12957 < _zz_dataOut_payload_0_13005);
  assign _zz_dataOut_payload_0_13388 = (_zz_dataOut_payload_0_13387 ? _zz_dataOut_payload_0_12957 : _zz_dataOut_payload_0_13005);
  assign _zz_dataOut_payload_0_13389 = (_zz_dataOut_payload_0_13387 ? _zz_dataOut_payload_0_13005 : _zz_dataOut_payload_0_12957);
  assign _zz_dataOut_payload_0_13390 = (_zz_dataOut_payload_0_12960 < _zz_dataOut_payload_0_13008);
  assign _zz_dataOut_payload_0_13391 = (_zz_dataOut_payload_0_13390 ? _zz_dataOut_payload_0_12960 : _zz_dataOut_payload_0_13008);
  assign _zz_dataOut_payload_0_13392 = (_zz_dataOut_payload_0_13390 ? _zz_dataOut_payload_0_13008 : _zz_dataOut_payload_0_12960);
  assign _zz_dataOut_payload_0_13393 = (_zz_dataOut_payload_0_12963 < _zz_dataOut_payload_0_13011);
  assign _zz_dataOut_payload_0_13394 = (_zz_dataOut_payload_0_13393 ? _zz_dataOut_payload_0_12963 : _zz_dataOut_payload_0_13011);
  assign _zz_dataOut_payload_0_13395 = (_zz_dataOut_payload_0_13393 ? _zz_dataOut_payload_0_13011 : _zz_dataOut_payload_0_12963);
  assign _zz_dataOut_payload_0_13396 = (_zz_dataOut_payload_0_12966 < _zz_dataOut_payload_0_13014);
  assign _zz_dataOut_payload_0_13397 = (_zz_dataOut_payload_0_13396 ? _zz_dataOut_payload_0_12966 : _zz_dataOut_payload_0_13014);
  assign _zz_dataOut_payload_0_13398 = (_zz_dataOut_payload_0_13396 ? _zz_dataOut_payload_0_13014 : _zz_dataOut_payload_0_12966);
  assign _zz_dataOut_payload_0_13399 = (_zz_dataOut_payload_0_12969 < _zz_dataOut_payload_0_13017);
  assign _zz_dataOut_payload_0_13400 = (_zz_dataOut_payload_0_13399 ? _zz_dataOut_payload_0_12969 : _zz_dataOut_payload_0_13017);
  assign _zz_dataOut_payload_0_13401 = (_zz_dataOut_payload_0_13399 ? _zz_dataOut_payload_0_13017 : _zz_dataOut_payload_0_12969);
  assign _zz_dataOut_payload_0_13402 = (_zz_dataOut_payload_0_12972 < _zz_dataOut_payload_0_13020);
  assign _zz_dataOut_payload_0_13403 = (_zz_dataOut_payload_0_13402 ? _zz_dataOut_payload_0_12972 : _zz_dataOut_payload_0_13020);
  assign _zz_dataOut_payload_0_13404 = (_zz_dataOut_payload_0_13402 ? _zz_dataOut_payload_0_13020 : _zz_dataOut_payload_0_12972);
  assign _zz_dataOut_payload_0_13405 = (_zz_dataOut_payload_0_12975 < _zz_dataOut_payload_0_13023);
  assign _zz_dataOut_payload_0_13406 = (_zz_dataOut_payload_0_13405 ? _zz_dataOut_payload_0_12975 : _zz_dataOut_payload_0_13023);
  assign _zz_dataOut_payload_0_13407 = (_zz_dataOut_payload_0_13405 ? _zz_dataOut_payload_0_13023 : _zz_dataOut_payload_0_12975);
  assign _zz_dataOut_payload_0_13408 = (_zz_dataOut_payload_0_13361 < _zz_dataOut_payload_0_13385);
  assign _zz_dataOut_payload_0_13409 = (_zz_dataOut_payload_0_13408 ? _zz_dataOut_payload_0_13361 : _zz_dataOut_payload_0_13385);
  assign _zz_dataOut_payload_0_13410 = (_zz_dataOut_payload_0_13408 ? _zz_dataOut_payload_0_13385 : _zz_dataOut_payload_0_13361);
  assign _zz_dataOut_payload_0_13411 = (_zz_dataOut_payload_0_13364 < _zz_dataOut_payload_0_13388);
  assign _zz_dataOut_payload_0_13412 = (_zz_dataOut_payload_0_13411 ? _zz_dataOut_payload_0_13364 : _zz_dataOut_payload_0_13388);
  assign _zz_dataOut_payload_0_13413 = (_zz_dataOut_payload_0_13411 ? _zz_dataOut_payload_0_13388 : _zz_dataOut_payload_0_13364);
  assign _zz_dataOut_payload_0_13414 = (_zz_dataOut_payload_0_13367 < _zz_dataOut_payload_0_13391);
  assign _zz_dataOut_payload_0_13415 = (_zz_dataOut_payload_0_13414 ? _zz_dataOut_payload_0_13367 : _zz_dataOut_payload_0_13391);
  assign _zz_dataOut_payload_0_13416 = (_zz_dataOut_payload_0_13414 ? _zz_dataOut_payload_0_13391 : _zz_dataOut_payload_0_13367);
  assign _zz_dataOut_payload_0_13417 = (_zz_dataOut_payload_0_13370 < _zz_dataOut_payload_0_13394);
  assign _zz_dataOut_payload_0_13418 = (_zz_dataOut_payload_0_13417 ? _zz_dataOut_payload_0_13370 : _zz_dataOut_payload_0_13394);
  assign _zz_dataOut_payload_0_13419 = (_zz_dataOut_payload_0_13417 ? _zz_dataOut_payload_0_13394 : _zz_dataOut_payload_0_13370);
  assign _zz_dataOut_payload_0_13420 = (_zz_dataOut_payload_0_13373 < _zz_dataOut_payload_0_13397);
  assign _zz_dataOut_payload_0_13421 = (_zz_dataOut_payload_0_13420 ? _zz_dataOut_payload_0_13373 : _zz_dataOut_payload_0_13397);
  assign _zz_dataOut_payload_0_13422 = (_zz_dataOut_payload_0_13420 ? _zz_dataOut_payload_0_13397 : _zz_dataOut_payload_0_13373);
  assign _zz_dataOut_payload_0_13423 = (_zz_dataOut_payload_0_13376 < _zz_dataOut_payload_0_13400);
  assign _zz_dataOut_payload_0_13424 = (_zz_dataOut_payload_0_13423 ? _zz_dataOut_payload_0_13376 : _zz_dataOut_payload_0_13400);
  assign _zz_dataOut_payload_0_13425 = (_zz_dataOut_payload_0_13423 ? _zz_dataOut_payload_0_13400 : _zz_dataOut_payload_0_13376);
  assign _zz_dataOut_payload_0_13426 = (_zz_dataOut_payload_0_13379 < _zz_dataOut_payload_0_13403);
  assign _zz_dataOut_payload_0_13427 = (_zz_dataOut_payload_0_13426 ? _zz_dataOut_payload_0_13379 : _zz_dataOut_payload_0_13403);
  assign _zz_dataOut_payload_0_13428 = (_zz_dataOut_payload_0_13426 ? _zz_dataOut_payload_0_13403 : _zz_dataOut_payload_0_13379);
  assign _zz_dataOut_payload_0_13429 = (_zz_dataOut_payload_0_13382 < _zz_dataOut_payload_0_13406);
  assign _zz_dataOut_payload_0_13430 = (_zz_dataOut_payload_0_13429 ? _zz_dataOut_payload_0_13382 : _zz_dataOut_payload_0_13406);
  assign _zz_dataOut_payload_0_13431 = (_zz_dataOut_payload_0_13429 ? _zz_dataOut_payload_0_13406 : _zz_dataOut_payload_0_13382);
  assign _zz_dataOut_payload_0_13432 = (_zz_dataOut_payload_0_13409 < _zz_dataOut_payload_0_13421);
  assign _zz_dataOut_payload_0_13433 = (_zz_dataOut_payload_0_13432 ? _zz_dataOut_payload_0_13409 : _zz_dataOut_payload_0_13421);
  assign _zz_dataOut_payload_0_13434 = (_zz_dataOut_payload_0_13432 ? _zz_dataOut_payload_0_13421 : _zz_dataOut_payload_0_13409);
  assign _zz_dataOut_payload_0_13435 = (_zz_dataOut_payload_0_13412 < _zz_dataOut_payload_0_13424);
  assign _zz_dataOut_payload_0_13436 = (_zz_dataOut_payload_0_13435 ? _zz_dataOut_payload_0_13412 : _zz_dataOut_payload_0_13424);
  assign _zz_dataOut_payload_0_13437 = (_zz_dataOut_payload_0_13435 ? _zz_dataOut_payload_0_13424 : _zz_dataOut_payload_0_13412);
  assign _zz_dataOut_payload_0_13438 = (_zz_dataOut_payload_0_13415 < _zz_dataOut_payload_0_13427);
  assign _zz_dataOut_payload_0_13439 = (_zz_dataOut_payload_0_13438 ? _zz_dataOut_payload_0_13415 : _zz_dataOut_payload_0_13427);
  assign _zz_dataOut_payload_0_13440 = (_zz_dataOut_payload_0_13438 ? _zz_dataOut_payload_0_13427 : _zz_dataOut_payload_0_13415);
  assign _zz_dataOut_payload_0_13441 = (_zz_dataOut_payload_0_13418 < _zz_dataOut_payload_0_13430);
  assign _zz_dataOut_payload_0_13442 = (_zz_dataOut_payload_0_13441 ? _zz_dataOut_payload_0_13418 : _zz_dataOut_payload_0_13430);
  assign _zz_dataOut_payload_0_13443 = (_zz_dataOut_payload_0_13441 ? _zz_dataOut_payload_0_13430 : _zz_dataOut_payload_0_13418);
  assign _zz_dataOut_payload_0_13444 = (_zz_dataOut_payload_0_13433 < _zz_dataOut_payload_0_13439);
  assign _zz_dataOut_payload_0_13445 = (_zz_dataOut_payload_0_13444 ? _zz_dataOut_payload_0_13433 : _zz_dataOut_payload_0_13439);
  assign _zz_dataOut_payload_0_13446 = (_zz_dataOut_payload_0_13444 ? _zz_dataOut_payload_0_13439 : _zz_dataOut_payload_0_13433);
  assign _zz_dataOut_payload_0_13447 = (_zz_dataOut_payload_0_13436 < _zz_dataOut_payload_0_13442);
  assign _zz_dataOut_payload_0_13448 = (_zz_dataOut_payload_0_13447 ? _zz_dataOut_payload_0_13436 : _zz_dataOut_payload_0_13442);
  assign _zz_dataOut_payload_0_13449 = (_zz_dataOut_payload_0_13447 ? _zz_dataOut_payload_0_13442 : _zz_dataOut_payload_0_13436);
  assign _zz_dataOut_payload_0_13450 = (_zz_dataOut_payload_0_13445 < _zz_dataOut_payload_0_13448);
  assign _zz_dataOut_payload_0_13451 = (_zz_dataOut_payload_0_13446 < _zz_dataOut_payload_0_13449);
  assign _zz_dataOut_payload_0_13456 = (_zz_dataOut_payload_0_13434 < _zz_dataOut_payload_0_13440);
  assign _zz_dataOut_payload_0_13457 = (_zz_dataOut_payload_0_13456 ? _zz_dataOut_payload_0_13434 : _zz_dataOut_payload_0_13440);
  assign _zz_dataOut_payload_0_13458 = (_zz_dataOut_payload_0_13456 ? _zz_dataOut_payload_0_13440 : _zz_dataOut_payload_0_13434);
  assign _zz_dataOut_payload_0_13459 = (_zz_dataOut_payload_0_13437 < _zz_dataOut_payload_0_13443);
  assign _zz_dataOut_payload_0_13460 = (_zz_dataOut_payload_0_13459 ? _zz_dataOut_payload_0_13437 : _zz_dataOut_payload_0_13443);
  assign _zz_dataOut_payload_0_13461 = (_zz_dataOut_payload_0_13459 ? _zz_dataOut_payload_0_13443 : _zz_dataOut_payload_0_13437);
  assign _zz_dataOut_payload_0_13462 = (_zz_dataOut_payload_0_13457 < _zz_dataOut_payload_0_13460);
  assign _zz_dataOut_payload_0_13463 = (_zz_dataOut_payload_0_13458 < _zz_dataOut_payload_0_13461);
  assign _zz_dataOut_payload_0_13476 = (_zz_dataOut_payload_0_13410 < _zz_dataOut_payload_0_13422);
  assign _zz_dataOut_payload_0_13477 = (_zz_dataOut_payload_0_13476 ? _zz_dataOut_payload_0_13410 : _zz_dataOut_payload_0_13422);
  assign _zz_dataOut_payload_0_13478 = (_zz_dataOut_payload_0_13476 ? _zz_dataOut_payload_0_13422 : _zz_dataOut_payload_0_13410);
  assign _zz_dataOut_payload_0_13479 = (_zz_dataOut_payload_0_13413 < _zz_dataOut_payload_0_13425);
  assign _zz_dataOut_payload_0_13480 = (_zz_dataOut_payload_0_13479 ? _zz_dataOut_payload_0_13413 : _zz_dataOut_payload_0_13425);
  assign _zz_dataOut_payload_0_13481 = (_zz_dataOut_payload_0_13479 ? _zz_dataOut_payload_0_13425 : _zz_dataOut_payload_0_13413);
  assign _zz_dataOut_payload_0_13482 = (_zz_dataOut_payload_0_13416 < _zz_dataOut_payload_0_13428);
  assign _zz_dataOut_payload_0_13483 = (_zz_dataOut_payload_0_13482 ? _zz_dataOut_payload_0_13416 : _zz_dataOut_payload_0_13428);
  assign _zz_dataOut_payload_0_13484 = (_zz_dataOut_payload_0_13482 ? _zz_dataOut_payload_0_13428 : _zz_dataOut_payload_0_13416);
  assign _zz_dataOut_payload_0_13485 = (_zz_dataOut_payload_0_13419 < _zz_dataOut_payload_0_13431);
  assign _zz_dataOut_payload_0_13486 = (_zz_dataOut_payload_0_13485 ? _zz_dataOut_payload_0_13419 : _zz_dataOut_payload_0_13431);
  assign _zz_dataOut_payload_0_13487 = (_zz_dataOut_payload_0_13485 ? _zz_dataOut_payload_0_13431 : _zz_dataOut_payload_0_13419);
  assign _zz_dataOut_payload_0_13488 = (_zz_dataOut_payload_0_13477 < _zz_dataOut_payload_0_13483);
  assign _zz_dataOut_payload_0_13489 = (_zz_dataOut_payload_0_13488 ? _zz_dataOut_payload_0_13477 : _zz_dataOut_payload_0_13483);
  assign _zz_dataOut_payload_0_13490 = (_zz_dataOut_payload_0_13488 ? _zz_dataOut_payload_0_13483 : _zz_dataOut_payload_0_13477);
  assign _zz_dataOut_payload_0_13491 = (_zz_dataOut_payload_0_13480 < _zz_dataOut_payload_0_13486);
  assign _zz_dataOut_payload_0_13492 = (_zz_dataOut_payload_0_13491 ? _zz_dataOut_payload_0_13480 : _zz_dataOut_payload_0_13486);
  assign _zz_dataOut_payload_0_13493 = (_zz_dataOut_payload_0_13491 ? _zz_dataOut_payload_0_13486 : _zz_dataOut_payload_0_13480);
  assign _zz_dataOut_payload_0_13494 = (_zz_dataOut_payload_0_13489 < _zz_dataOut_payload_0_13492);
  assign _zz_dataOut_payload_0_13495 = (_zz_dataOut_payload_0_13490 < _zz_dataOut_payload_0_13493);
  assign _zz_dataOut_payload_0_13500 = (_zz_dataOut_payload_0_13478 < _zz_dataOut_payload_0_13484);
  assign _zz_dataOut_payload_0_13501 = (_zz_dataOut_payload_0_13500 ? _zz_dataOut_payload_0_13478 : _zz_dataOut_payload_0_13484);
  assign _zz_dataOut_payload_0_13502 = (_zz_dataOut_payload_0_13500 ? _zz_dataOut_payload_0_13484 : _zz_dataOut_payload_0_13478);
  assign _zz_dataOut_payload_0_13503 = (_zz_dataOut_payload_0_13481 < _zz_dataOut_payload_0_13487);
  assign _zz_dataOut_payload_0_13504 = (_zz_dataOut_payload_0_13503 ? _zz_dataOut_payload_0_13481 : _zz_dataOut_payload_0_13487);
  assign _zz_dataOut_payload_0_13505 = (_zz_dataOut_payload_0_13503 ? _zz_dataOut_payload_0_13487 : _zz_dataOut_payload_0_13481);
  assign _zz_dataOut_payload_0_13506 = (_zz_dataOut_payload_0_13501 < _zz_dataOut_payload_0_13504);
  assign _zz_dataOut_payload_0_13507 = (_zz_dataOut_payload_0_13502 < _zz_dataOut_payload_0_13505);
  assign _zz_dataOut_payload_0_13536 = (_zz_dataOut_payload_0_13362 < _zz_dataOut_payload_0_13386);
  assign _zz_dataOut_payload_0_13537 = (_zz_dataOut_payload_0_13536 ? _zz_dataOut_payload_0_13362 : _zz_dataOut_payload_0_13386);
  assign _zz_dataOut_payload_0_13538 = (_zz_dataOut_payload_0_13536 ? _zz_dataOut_payload_0_13386 : _zz_dataOut_payload_0_13362);
  assign _zz_dataOut_payload_0_13539 = (_zz_dataOut_payload_0_13365 < _zz_dataOut_payload_0_13389);
  assign _zz_dataOut_payload_0_13540 = (_zz_dataOut_payload_0_13539 ? _zz_dataOut_payload_0_13365 : _zz_dataOut_payload_0_13389);
  assign _zz_dataOut_payload_0_13541 = (_zz_dataOut_payload_0_13539 ? _zz_dataOut_payload_0_13389 : _zz_dataOut_payload_0_13365);
  assign _zz_dataOut_payload_0_13542 = (_zz_dataOut_payload_0_13368 < _zz_dataOut_payload_0_13392);
  assign _zz_dataOut_payload_0_13543 = (_zz_dataOut_payload_0_13542 ? _zz_dataOut_payload_0_13368 : _zz_dataOut_payload_0_13392);
  assign _zz_dataOut_payload_0_13544 = (_zz_dataOut_payload_0_13542 ? _zz_dataOut_payload_0_13392 : _zz_dataOut_payload_0_13368);
  assign _zz_dataOut_payload_0_13545 = (_zz_dataOut_payload_0_13371 < _zz_dataOut_payload_0_13395);
  assign _zz_dataOut_payload_0_13546 = (_zz_dataOut_payload_0_13545 ? _zz_dataOut_payload_0_13371 : _zz_dataOut_payload_0_13395);
  assign _zz_dataOut_payload_0_13547 = (_zz_dataOut_payload_0_13545 ? _zz_dataOut_payload_0_13395 : _zz_dataOut_payload_0_13371);
  assign _zz_dataOut_payload_0_13548 = (_zz_dataOut_payload_0_13374 < _zz_dataOut_payload_0_13398);
  assign _zz_dataOut_payload_0_13549 = (_zz_dataOut_payload_0_13548 ? _zz_dataOut_payload_0_13374 : _zz_dataOut_payload_0_13398);
  assign _zz_dataOut_payload_0_13550 = (_zz_dataOut_payload_0_13548 ? _zz_dataOut_payload_0_13398 : _zz_dataOut_payload_0_13374);
  assign _zz_dataOut_payload_0_13551 = (_zz_dataOut_payload_0_13377 < _zz_dataOut_payload_0_13401);
  assign _zz_dataOut_payload_0_13552 = (_zz_dataOut_payload_0_13551 ? _zz_dataOut_payload_0_13377 : _zz_dataOut_payload_0_13401);
  assign _zz_dataOut_payload_0_13553 = (_zz_dataOut_payload_0_13551 ? _zz_dataOut_payload_0_13401 : _zz_dataOut_payload_0_13377);
  assign _zz_dataOut_payload_0_13554 = (_zz_dataOut_payload_0_13380 < _zz_dataOut_payload_0_13404);
  assign _zz_dataOut_payload_0_13555 = (_zz_dataOut_payload_0_13554 ? _zz_dataOut_payload_0_13380 : _zz_dataOut_payload_0_13404);
  assign _zz_dataOut_payload_0_13556 = (_zz_dataOut_payload_0_13554 ? _zz_dataOut_payload_0_13404 : _zz_dataOut_payload_0_13380);
  assign _zz_dataOut_payload_0_13557 = (_zz_dataOut_payload_0_13383 < _zz_dataOut_payload_0_13407);
  assign _zz_dataOut_payload_0_13558 = (_zz_dataOut_payload_0_13557 ? _zz_dataOut_payload_0_13383 : _zz_dataOut_payload_0_13407);
  assign _zz_dataOut_payload_0_13559 = (_zz_dataOut_payload_0_13557 ? _zz_dataOut_payload_0_13407 : _zz_dataOut_payload_0_13383);
  assign _zz_dataOut_payload_0_13560 = (_zz_dataOut_payload_0_13537 < _zz_dataOut_payload_0_13549);
  assign _zz_dataOut_payload_0_13561 = (_zz_dataOut_payload_0_13560 ? _zz_dataOut_payload_0_13537 : _zz_dataOut_payload_0_13549);
  assign _zz_dataOut_payload_0_13562 = (_zz_dataOut_payload_0_13560 ? _zz_dataOut_payload_0_13549 : _zz_dataOut_payload_0_13537);
  assign _zz_dataOut_payload_0_13563 = (_zz_dataOut_payload_0_13540 < _zz_dataOut_payload_0_13552);
  assign _zz_dataOut_payload_0_13564 = (_zz_dataOut_payload_0_13563 ? _zz_dataOut_payload_0_13540 : _zz_dataOut_payload_0_13552);
  assign _zz_dataOut_payload_0_13565 = (_zz_dataOut_payload_0_13563 ? _zz_dataOut_payload_0_13552 : _zz_dataOut_payload_0_13540);
  assign _zz_dataOut_payload_0_13566 = (_zz_dataOut_payload_0_13543 < _zz_dataOut_payload_0_13555);
  assign _zz_dataOut_payload_0_13567 = (_zz_dataOut_payload_0_13566 ? _zz_dataOut_payload_0_13543 : _zz_dataOut_payload_0_13555);
  assign _zz_dataOut_payload_0_13568 = (_zz_dataOut_payload_0_13566 ? _zz_dataOut_payload_0_13555 : _zz_dataOut_payload_0_13543);
  assign _zz_dataOut_payload_0_13569 = (_zz_dataOut_payload_0_13546 < _zz_dataOut_payload_0_13558);
  assign _zz_dataOut_payload_0_13570 = (_zz_dataOut_payload_0_13569 ? _zz_dataOut_payload_0_13546 : _zz_dataOut_payload_0_13558);
  assign _zz_dataOut_payload_0_13571 = (_zz_dataOut_payload_0_13569 ? _zz_dataOut_payload_0_13558 : _zz_dataOut_payload_0_13546);
  assign _zz_dataOut_payload_0_13572 = (_zz_dataOut_payload_0_13561 < _zz_dataOut_payload_0_13567);
  assign _zz_dataOut_payload_0_13573 = (_zz_dataOut_payload_0_13572 ? _zz_dataOut_payload_0_13561 : _zz_dataOut_payload_0_13567);
  assign _zz_dataOut_payload_0_13574 = (_zz_dataOut_payload_0_13572 ? _zz_dataOut_payload_0_13567 : _zz_dataOut_payload_0_13561);
  assign _zz_dataOut_payload_0_13575 = (_zz_dataOut_payload_0_13564 < _zz_dataOut_payload_0_13570);
  assign _zz_dataOut_payload_0_13576 = (_zz_dataOut_payload_0_13575 ? _zz_dataOut_payload_0_13564 : _zz_dataOut_payload_0_13570);
  assign _zz_dataOut_payload_0_13577 = (_zz_dataOut_payload_0_13575 ? _zz_dataOut_payload_0_13570 : _zz_dataOut_payload_0_13564);
  assign _zz_dataOut_payload_0_13578 = (_zz_dataOut_payload_0_13573 < _zz_dataOut_payload_0_13576);
  assign _zz_dataOut_payload_0_13579 = (_zz_dataOut_payload_0_13574 < _zz_dataOut_payload_0_13577);
  assign _zz_dataOut_payload_0_13584 = (_zz_dataOut_payload_0_13562 < _zz_dataOut_payload_0_13568);
  assign _zz_dataOut_payload_0_13585 = (_zz_dataOut_payload_0_13584 ? _zz_dataOut_payload_0_13562 : _zz_dataOut_payload_0_13568);
  assign _zz_dataOut_payload_0_13586 = (_zz_dataOut_payload_0_13584 ? _zz_dataOut_payload_0_13568 : _zz_dataOut_payload_0_13562);
  assign _zz_dataOut_payload_0_13587 = (_zz_dataOut_payload_0_13565 < _zz_dataOut_payload_0_13571);
  assign _zz_dataOut_payload_0_13588 = (_zz_dataOut_payload_0_13587 ? _zz_dataOut_payload_0_13565 : _zz_dataOut_payload_0_13571);
  assign _zz_dataOut_payload_0_13589 = (_zz_dataOut_payload_0_13587 ? _zz_dataOut_payload_0_13571 : _zz_dataOut_payload_0_13565);
  assign _zz_dataOut_payload_0_13590 = (_zz_dataOut_payload_0_13585 < _zz_dataOut_payload_0_13588);
  assign _zz_dataOut_payload_0_13591 = (_zz_dataOut_payload_0_13586 < _zz_dataOut_payload_0_13589);
  assign _zz_dataOut_payload_0_13604 = (_zz_dataOut_payload_0_13538 < _zz_dataOut_payload_0_13550);
  assign _zz_dataOut_payload_0_13605 = (_zz_dataOut_payload_0_13604 ? _zz_dataOut_payload_0_13538 : _zz_dataOut_payload_0_13550);
  assign _zz_dataOut_payload_0_13606 = (_zz_dataOut_payload_0_13604 ? _zz_dataOut_payload_0_13550 : _zz_dataOut_payload_0_13538);
  assign _zz_dataOut_payload_0_13607 = (_zz_dataOut_payload_0_13541 < _zz_dataOut_payload_0_13553);
  assign _zz_dataOut_payload_0_13608 = (_zz_dataOut_payload_0_13607 ? _zz_dataOut_payload_0_13541 : _zz_dataOut_payload_0_13553);
  assign _zz_dataOut_payload_0_13609 = (_zz_dataOut_payload_0_13607 ? _zz_dataOut_payload_0_13553 : _zz_dataOut_payload_0_13541);
  assign _zz_dataOut_payload_0_13610 = (_zz_dataOut_payload_0_13544 < _zz_dataOut_payload_0_13556);
  assign _zz_dataOut_payload_0_13611 = (_zz_dataOut_payload_0_13610 ? _zz_dataOut_payload_0_13544 : _zz_dataOut_payload_0_13556);
  assign _zz_dataOut_payload_0_13612 = (_zz_dataOut_payload_0_13610 ? _zz_dataOut_payload_0_13556 : _zz_dataOut_payload_0_13544);
  assign _zz_dataOut_payload_0_13613 = (_zz_dataOut_payload_0_13547 < _zz_dataOut_payload_0_13559);
  assign _zz_dataOut_payload_0_13614 = (_zz_dataOut_payload_0_13613 ? _zz_dataOut_payload_0_13547 : _zz_dataOut_payload_0_13559);
  assign _zz_dataOut_payload_0_13615 = (_zz_dataOut_payload_0_13613 ? _zz_dataOut_payload_0_13559 : _zz_dataOut_payload_0_13547);
  assign _zz_dataOut_payload_0_13616 = (_zz_dataOut_payload_0_13605 < _zz_dataOut_payload_0_13611);
  assign _zz_dataOut_payload_0_13617 = (_zz_dataOut_payload_0_13616 ? _zz_dataOut_payload_0_13605 : _zz_dataOut_payload_0_13611);
  assign _zz_dataOut_payload_0_13618 = (_zz_dataOut_payload_0_13616 ? _zz_dataOut_payload_0_13611 : _zz_dataOut_payload_0_13605);
  assign _zz_dataOut_payload_0_13619 = (_zz_dataOut_payload_0_13608 < _zz_dataOut_payload_0_13614);
  assign _zz_dataOut_payload_0_13620 = (_zz_dataOut_payload_0_13619 ? _zz_dataOut_payload_0_13608 : _zz_dataOut_payload_0_13614);
  assign _zz_dataOut_payload_0_13621 = (_zz_dataOut_payload_0_13619 ? _zz_dataOut_payload_0_13614 : _zz_dataOut_payload_0_13608);
  assign _zz_dataOut_payload_0_13622 = (_zz_dataOut_payload_0_13617 < _zz_dataOut_payload_0_13620);
  assign _zz_dataOut_payload_0_13623 = (_zz_dataOut_payload_0_13618 < _zz_dataOut_payload_0_13621);
  assign _zz_dataOut_payload_0_13628 = (_zz_dataOut_payload_0_13606 < _zz_dataOut_payload_0_13612);
  assign _zz_dataOut_payload_0_13629 = (_zz_dataOut_payload_0_13628 ? _zz_dataOut_payload_0_13606 : _zz_dataOut_payload_0_13612);
  assign _zz_dataOut_payload_0_13630 = (_zz_dataOut_payload_0_13628 ? _zz_dataOut_payload_0_13612 : _zz_dataOut_payload_0_13606);
  assign _zz_dataOut_payload_0_13631 = (_zz_dataOut_payload_0_13609 < _zz_dataOut_payload_0_13615);
  assign _zz_dataOut_payload_0_13632 = (_zz_dataOut_payload_0_13631 ? _zz_dataOut_payload_0_13609 : _zz_dataOut_payload_0_13615);
  assign _zz_dataOut_payload_0_13633 = (_zz_dataOut_payload_0_13631 ? _zz_dataOut_payload_0_13615 : _zz_dataOut_payload_0_13609);
  assign _zz_dataOut_payload_0_13634 = (_zz_dataOut_payload_0_13629 < _zz_dataOut_payload_0_13632);
  assign _zz_dataOut_payload_0_13635 = (_zz_dataOut_payload_0_13630 < _zz_dataOut_payload_0_13633);
  assign _zz_dataOut_payload_0_13888 = (_zz_dataOut_payload_0_11776 < _zz_dataOut_payload_0_11903);
  assign _zz_dataOut_payload_0_13889 = (_zz_dataOut_payload_0_13888 ? _zz_dataOut_payload_0_11776 : _zz_dataOut_payload_0_11903);
  assign _zz_dataOut_payload_0_13890 = (_zz_dataOut_payload_0_13888 ? _zz_dataOut_payload_0_11903 : _zz_dataOut_payload_0_11776);
  assign _zz_dataOut_payload_0_13891 = (_zz_dataOut_payload_0_11777 < _zz_dataOut_payload_0_11902);
  assign _zz_dataOut_payload_0_13892 = (_zz_dataOut_payload_0_13891 ? _zz_dataOut_payload_0_11777 : _zz_dataOut_payload_0_11902);
  assign _zz_dataOut_payload_0_13893 = (_zz_dataOut_payload_0_13891 ? _zz_dataOut_payload_0_11902 : _zz_dataOut_payload_0_11777);
  assign _zz_dataOut_payload_0_13894 = (_zz_dataOut_payload_0_11778 < _zz_dataOut_payload_0_11901);
  assign _zz_dataOut_payload_0_13895 = (_zz_dataOut_payload_0_13894 ? _zz_dataOut_payload_0_11778 : _zz_dataOut_payload_0_11901);
  assign _zz_dataOut_payload_0_13896 = (_zz_dataOut_payload_0_13894 ? _zz_dataOut_payload_0_11901 : _zz_dataOut_payload_0_11778);
  assign _zz_dataOut_payload_0_13897 = (_zz_dataOut_payload_0_11779 < _zz_dataOut_payload_0_11900);
  assign _zz_dataOut_payload_0_13898 = (_zz_dataOut_payload_0_13897 ? _zz_dataOut_payload_0_11779 : _zz_dataOut_payload_0_11900);
  assign _zz_dataOut_payload_0_13899 = (_zz_dataOut_payload_0_13897 ? _zz_dataOut_payload_0_11900 : _zz_dataOut_payload_0_11779);
  assign _zz_dataOut_payload_0_13900 = (_zz_dataOut_payload_0_11780 < _zz_dataOut_payload_0_11899);
  assign _zz_dataOut_payload_0_13901 = (_zz_dataOut_payload_0_13900 ? _zz_dataOut_payload_0_11780 : _zz_dataOut_payload_0_11899);
  assign _zz_dataOut_payload_0_13902 = (_zz_dataOut_payload_0_13900 ? _zz_dataOut_payload_0_11899 : _zz_dataOut_payload_0_11780);
  assign _zz_dataOut_payload_0_13903 = (_zz_dataOut_payload_0_11781 < _zz_dataOut_payload_0_11898);
  assign _zz_dataOut_payload_0_13904 = (_zz_dataOut_payload_0_13903 ? _zz_dataOut_payload_0_11781 : _zz_dataOut_payload_0_11898);
  assign _zz_dataOut_payload_0_13905 = (_zz_dataOut_payload_0_13903 ? _zz_dataOut_payload_0_11898 : _zz_dataOut_payload_0_11781);
  assign _zz_dataOut_payload_0_13906 = (_zz_dataOut_payload_0_11782 < _zz_dataOut_payload_0_11897);
  assign _zz_dataOut_payload_0_13907 = (_zz_dataOut_payload_0_13906 ? _zz_dataOut_payload_0_11782 : _zz_dataOut_payload_0_11897);
  assign _zz_dataOut_payload_0_13908 = (_zz_dataOut_payload_0_13906 ? _zz_dataOut_payload_0_11897 : _zz_dataOut_payload_0_11782);
  assign _zz_dataOut_payload_0_13909 = (_zz_dataOut_payload_0_11783 < _zz_dataOut_payload_0_11896);
  assign _zz_dataOut_payload_0_13910 = (_zz_dataOut_payload_0_13909 ? _zz_dataOut_payload_0_11783 : _zz_dataOut_payload_0_11896);
  assign _zz_dataOut_payload_0_13911 = (_zz_dataOut_payload_0_13909 ? _zz_dataOut_payload_0_11896 : _zz_dataOut_payload_0_11783);
  assign _zz_dataOut_payload_0_13912 = (_zz_dataOut_payload_0_11784 < _zz_dataOut_payload_0_11895);
  assign _zz_dataOut_payload_0_13913 = (_zz_dataOut_payload_0_13912 ? _zz_dataOut_payload_0_11784 : _zz_dataOut_payload_0_11895);
  assign _zz_dataOut_payload_0_13914 = (_zz_dataOut_payload_0_13912 ? _zz_dataOut_payload_0_11895 : _zz_dataOut_payload_0_11784);
  assign _zz_dataOut_payload_0_13915 = (_zz_dataOut_payload_0_11785 < _zz_dataOut_payload_0_11894);
  assign _zz_dataOut_payload_0_13916 = (_zz_dataOut_payload_0_13915 ? _zz_dataOut_payload_0_11785 : _zz_dataOut_payload_0_11894);
  assign _zz_dataOut_payload_0_13917 = (_zz_dataOut_payload_0_13915 ? _zz_dataOut_payload_0_11894 : _zz_dataOut_payload_0_11785);
  assign _zz_dataOut_payload_0_13918 = (_zz_dataOut_payload_0_11786 < _zz_dataOut_payload_0_11893);
  assign _zz_dataOut_payload_0_13919 = (_zz_dataOut_payload_0_13918 ? _zz_dataOut_payload_0_11786 : _zz_dataOut_payload_0_11893);
  assign _zz_dataOut_payload_0_13920 = (_zz_dataOut_payload_0_13918 ? _zz_dataOut_payload_0_11893 : _zz_dataOut_payload_0_11786);
  assign _zz_dataOut_payload_0_13921 = (_zz_dataOut_payload_0_11787 < _zz_dataOut_payload_0_11892);
  assign _zz_dataOut_payload_0_13922 = (_zz_dataOut_payload_0_13921 ? _zz_dataOut_payload_0_11787 : _zz_dataOut_payload_0_11892);
  assign _zz_dataOut_payload_0_13923 = (_zz_dataOut_payload_0_13921 ? _zz_dataOut_payload_0_11892 : _zz_dataOut_payload_0_11787);
  assign _zz_dataOut_payload_0_13924 = (_zz_dataOut_payload_0_11788 < _zz_dataOut_payload_0_11891);
  assign _zz_dataOut_payload_0_13925 = (_zz_dataOut_payload_0_13924 ? _zz_dataOut_payload_0_11788 : _zz_dataOut_payload_0_11891);
  assign _zz_dataOut_payload_0_13926 = (_zz_dataOut_payload_0_13924 ? _zz_dataOut_payload_0_11891 : _zz_dataOut_payload_0_11788);
  assign _zz_dataOut_payload_0_13927 = (_zz_dataOut_payload_0_11789 < _zz_dataOut_payload_0_11890);
  assign _zz_dataOut_payload_0_13928 = (_zz_dataOut_payload_0_13927 ? _zz_dataOut_payload_0_11789 : _zz_dataOut_payload_0_11890);
  assign _zz_dataOut_payload_0_13929 = (_zz_dataOut_payload_0_13927 ? _zz_dataOut_payload_0_11890 : _zz_dataOut_payload_0_11789);
  assign _zz_dataOut_payload_0_13930 = (_zz_dataOut_payload_0_11790 < _zz_dataOut_payload_0_11889);
  assign _zz_dataOut_payload_0_13931 = (_zz_dataOut_payload_0_13930 ? _zz_dataOut_payload_0_11790 : _zz_dataOut_payload_0_11889);
  assign _zz_dataOut_payload_0_13932 = (_zz_dataOut_payload_0_13930 ? _zz_dataOut_payload_0_11889 : _zz_dataOut_payload_0_11790);
  assign _zz_dataOut_payload_0_13933 = (_zz_dataOut_payload_0_11791 < _zz_dataOut_payload_0_11888);
  assign _zz_dataOut_payload_0_13934 = (_zz_dataOut_payload_0_13933 ? _zz_dataOut_payload_0_11791 : _zz_dataOut_payload_0_11888);
  assign _zz_dataOut_payload_0_13935 = (_zz_dataOut_payload_0_13933 ? _zz_dataOut_payload_0_11888 : _zz_dataOut_payload_0_11791);
  assign _zz_dataOut_payload_0_13936 = (_zz_dataOut_payload_0_11792 < _zz_dataOut_payload_0_11887);
  assign _zz_dataOut_payload_0_13937 = (_zz_dataOut_payload_0_13936 ? _zz_dataOut_payload_0_11792 : _zz_dataOut_payload_0_11887);
  assign _zz_dataOut_payload_0_13938 = (_zz_dataOut_payload_0_13936 ? _zz_dataOut_payload_0_11887 : _zz_dataOut_payload_0_11792);
  assign _zz_dataOut_payload_0_13939 = (_zz_dataOut_payload_0_11793 < _zz_dataOut_payload_0_11886);
  assign _zz_dataOut_payload_0_13940 = (_zz_dataOut_payload_0_13939 ? _zz_dataOut_payload_0_11793 : _zz_dataOut_payload_0_11886);
  assign _zz_dataOut_payload_0_13941 = (_zz_dataOut_payload_0_13939 ? _zz_dataOut_payload_0_11886 : _zz_dataOut_payload_0_11793);
  assign _zz_dataOut_payload_0_13942 = (_zz_dataOut_payload_0_11794 < _zz_dataOut_payload_0_11885);
  assign _zz_dataOut_payload_0_13943 = (_zz_dataOut_payload_0_13942 ? _zz_dataOut_payload_0_11794 : _zz_dataOut_payload_0_11885);
  assign _zz_dataOut_payload_0_13944 = (_zz_dataOut_payload_0_13942 ? _zz_dataOut_payload_0_11885 : _zz_dataOut_payload_0_11794);
  assign _zz_dataOut_payload_0_13945 = (_zz_dataOut_payload_0_11795 < _zz_dataOut_payload_0_11884);
  assign _zz_dataOut_payload_0_13946 = (_zz_dataOut_payload_0_13945 ? _zz_dataOut_payload_0_11795 : _zz_dataOut_payload_0_11884);
  assign _zz_dataOut_payload_0_13947 = (_zz_dataOut_payload_0_13945 ? _zz_dataOut_payload_0_11884 : _zz_dataOut_payload_0_11795);
  assign _zz_dataOut_payload_0_13948 = (_zz_dataOut_payload_0_11796 < _zz_dataOut_payload_0_11883);
  assign _zz_dataOut_payload_0_13949 = (_zz_dataOut_payload_0_13948 ? _zz_dataOut_payload_0_11796 : _zz_dataOut_payload_0_11883);
  assign _zz_dataOut_payload_0_13950 = (_zz_dataOut_payload_0_13948 ? _zz_dataOut_payload_0_11883 : _zz_dataOut_payload_0_11796);
  assign _zz_dataOut_payload_0_13951 = (_zz_dataOut_payload_0_11797 < _zz_dataOut_payload_0_11882);
  assign _zz_dataOut_payload_0_13952 = (_zz_dataOut_payload_0_13951 ? _zz_dataOut_payload_0_11797 : _zz_dataOut_payload_0_11882);
  assign _zz_dataOut_payload_0_13953 = (_zz_dataOut_payload_0_13951 ? _zz_dataOut_payload_0_11882 : _zz_dataOut_payload_0_11797);
  assign _zz_dataOut_payload_0_13954 = (_zz_dataOut_payload_0_11798 < _zz_dataOut_payload_0_11881);
  assign _zz_dataOut_payload_0_13955 = (_zz_dataOut_payload_0_13954 ? _zz_dataOut_payload_0_11798 : _zz_dataOut_payload_0_11881);
  assign _zz_dataOut_payload_0_13956 = (_zz_dataOut_payload_0_13954 ? _zz_dataOut_payload_0_11881 : _zz_dataOut_payload_0_11798);
  assign _zz_dataOut_payload_0_13957 = (_zz_dataOut_payload_0_11799 < _zz_dataOut_payload_0_11880);
  assign _zz_dataOut_payload_0_13958 = (_zz_dataOut_payload_0_13957 ? _zz_dataOut_payload_0_11799 : _zz_dataOut_payload_0_11880);
  assign _zz_dataOut_payload_0_13959 = (_zz_dataOut_payload_0_13957 ? _zz_dataOut_payload_0_11880 : _zz_dataOut_payload_0_11799);
  assign _zz_dataOut_payload_0_13960 = (_zz_dataOut_payload_0_11800 < _zz_dataOut_payload_0_11879);
  assign _zz_dataOut_payload_0_13961 = (_zz_dataOut_payload_0_13960 ? _zz_dataOut_payload_0_11800 : _zz_dataOut_payload_0_11879);
  assign _zz_dataOut_payload_0_13962 = (_zz_dataOut_payload_0_13960 ? _zz_dataOut_payload_0_11879 : _zz_dataOut_payload_0_11800);
  assign _zz_dataOut_payload_0_13963 = (_zz_dataOut_payload_0_11801 < _zz_dataOut_payload_0_11878);
  assign _zz_dataOut_payload_0_13964 = (_zz_dataOut_payload_0_13963 ? _zz_dataOut_payload_0_11801 : _zz_dataOut_payload_0_11878);
  assign _zz_dataOut_payload_0_13965 = (_zz_dataOut_payload_0_13963 ? _zz_dataOut_payload_0_11878 : _zz_dataOut_payload_0_11801);
  assign _zz_dataOut_payload_0_13966 = (_zz_dataOut_payload_0_11802 < _zz_dataOut_payload_0_11877);
  assign _zz_dataOut_payload_0_13967 = (_zz_dataOut_payload_0_13966 ? _zz_dataOut_payload_0_11802 : _zz_dataOut_payload_0_11877);
  assign _zz_dataOut_payload_0_13968 = (_zz_dataOut_payload_0_13966 ? _zz_dataOut_payload_0_11877 : _zz_dataOut_payload_0_11802);
  assign _zz_dataOut_payload_0_13969 = (_zz_dataOut_payload_0_11803 < _zz_dataOut_payload_0_11876);
  assign _zz_dataOut_payload_0_13970 = (_zz_dataOut_payload_0_13969 ? _zz_dataOut_payload_0_11803 : _zz_dataOut_payload_0_11876);
  assign _zz_dataOut_payload_0_13971 = (_zz_dataOut_payload_0_13969 ? _zz_dataOut_payload_0_11876 : _zz_dataOut_payload_0_11803);
  assign _zz_dataOut_payload_0_13972 = (_zz_dataOut_payload_0_11804 < _zz_dataOut_payload_0_11875);
  assign _zz_dataOut_payload_0_13973 = (_zz_dataOut_payload_0_13972 ? _zz_dataOut_payload_0_11804 : _zz_dataOut_payload_0_11875);
  assign _zz_dataOut_payload_0_13974 = (_zz_dataOut_payload_0_13972 ? _zz_dataOut_payload_0_11875 : _zz_dataOut_payload_0_11804);
  assign _zz_dataOut_payload_0_13975 = (_zz_dataOut_payload_0_11805 < _zz_dataOut_payload_0_11874);
  assign _zz_dataOut_payload_0_13976 = (_zz_dataOut_payload_0_13975 ? _zz_dataOut_payload_0_11805 : _zz_dataOut_payload_0_11874);
  assign _zz_dataOut_payload_0_13977 = (_zz_dataOut_payload_0_13975 ? _zz_dataOut_payload_0_11874 : _zz_dataOut_payload_0_11805);
  assign _zz_dataOut_payload_0_13978 = (_zz_dataOut_payload_0_11806 < _zz_dataOut_payload_0_11873);
  assign _zz_dataOut_payload_0_13979 = (_zz_dataOut_payload_0_13978 ? _zz_dataOut_payload_0_11806 : _zz_dataOut_payload_0_11873);
  assign _zz_dataOut_payload_0_13980 = (_zz_dataOut_payload_0_13978 ? _zz_dataOut_payload_0_11873 : _zz_dataOut_payload_0_11806);
  assign _zz_dataOut_payload_0_13981 = (_zz_dataOut_payload_0_11807 < _zz_dataOut_payload_0_11872);
  assign _zz_dataOut_payload_0_13982 = (_zz_dataOut_payload_0_13981 ? _zz_dataOut_payload_0_11807 : _zz_dataOut_payload_0_11872);
  assign _zz_dataOut_payload_0_13983 = (_zz_dataOut_payload_0_13981 ? _zz_dataOut_payload_0_11872 : _zz_dataOut_payload_0_11807);
  assign _zz_dataOut_payload_0_13984 = (_zz_dataOut_payload_0_11808 < _zz_dataOut_payload_0_11871);
  assign _zz_dataOut_payload_0_13985 = (_zz_dataOut_payload_0_13984 ? _zz_dataOut_payload_0_11808 : _zz_dataOut_payload_0_11871);
  assign _zz_dataOut_payload_0_13986 = (_zz_dataOut_payload_0_13984 ? _zz_dataOut_payload_0_11871 : _zz_dataOut_payload_0_11808);
  assign _zz_dataOut_payload_0_13987 = (_zz_dataOut_payload_0_11809 < _zz_dataOut_payload_0_11870);
  assign _zz_dataOut_payload_0_13988 = (_zz_dataOut_payload_0_13987 ? _zz_dataOut_payload_0_11809 : _zz_dataOut_payload_0_11870);
  assign _zz_dataOut_payload_0_13989 = (_zz_dataOut_payload_0_13987 ? _zz_dataOut_payload_0_11870 : _zz_dataOut_payload_0_11809);
  assign _zz_dataOut_payload_0_13990 = (_zz_dataOut_payload_0_11810 < _zz_dataOut_payload_0_11869);
  assign _zz_dataOut_payload_0_13991 = (_zz_dataOut_payload_0_13990 ? _zz_dataOut_payload_0_11810 : _zz_dataOut_payload_0_11869);
  assign _zz_dataOut_payload_0_13992 = (_zz_dataOut_payload_0_13990 ? _zz_dataOut_payload_0_11869 : _zz_dataOut_payload_0_11810);
  assign _zz_dataOut_payload_0_13993 = (_zz_dataOut_payload_0_11811 < _zz_dataOut_payload_0_11868);
  assign _zz_dataOut_payload_0_13994 = (_zz_dataOut_payload_0_13993 ? _zz_dataOut_payload_0_11811 : _zz_dataOut_payload_0_11868);
  assign _zz_dataOut_payload_0_13995 = (_zz_dataOut_payload_0_13993 ? _zz_dataOut_payload_0_11868 : _zz_dataOut_payload_0_11811);
  assign _zz_dataOut_payload_0_13996 = (_zz_dataOut_payload_0_11812 < _zz_dataOut_payload_0_11867);
  assign _zz_dataOut_payload_0_13997 = (_zz_dataOut_payload_0_13996 ? _zz_dataOut_payload_0_11812 : _zz_dataOut_payload_0_11867);
  assign _zz_dataOut_payload_0_13998 = (_zz_dataOut_payload_0_13996 ? _zz_dataOut_payload_0_11867 : _zz_dataOut_payload_0_11812);
  assign _zz_dataOut_payload_0_13999 = (_zz_dataOut_payload_0_11813 < _zz_dataOut_payload_0_11866);
  assign _zz_dataOut_payload_0_14000 = (_zz_dataOut_payload_0_13999 ? _zz_dataOut_payload_0_11813 : _zz_dataOut_payload_0_11866);
  assign _zz_dataOut_payload_0_14001 = (_zz_dataOut_payload_0_13999 ? _zz_dataOut_payload_0_11866 : _zz_dataOut_payload_0_11813);
  assign _zz_dataOut_payload_0_14002 = (_zz_dataOut_payload_0_11814 < _zz_dataOut_payload_0_11865);
  assign _zz_dataOut_payload_0_14003 = (_zz_dataOut_payload_0_14002 ? _zz_dataOut_payload_0_11814 : _zz_dataOut_payload_0_11865);
  assign _zz_dataOut_payload_0_14004 = (_zz_dataOut_payload_0_14002 ? _zz_dataOut_payload_0_11865 : _zz_dataOut_payload_0_11814);
  assign _zz_dataOut_payload_0_14005 = (_zz_dataOut_payload_0_11815 < _zz_dataOut_payload_0_11864);
  assign _zz_dataOut_payload_0_14006 = (_zz_dataOut_payload_0_14005 ? _zz_dataOut_payload_0_11815 : _zz_dataOut_payload_0_11864);
  assign _zz_dataOut_payload_0_14007 = (_zz_dataOut_payload_0_14005 ? _zz_dataOut_payload_0_11864 : _zz_dataOut_payload_0_11815);
  assign _zz_dataOut_payload_0_14008 = (_zz_dataOut_payload_0_11816 < _zz_dataOut_payload_0_11863);
  assign _zz_dataOut_payload_0_14009 = (_zz_dataOut_payload_0_14008 ? _zz_dataOut_payload_0_11816 : _zz_dataOut_payload_0_11863);
  assign _zz_dataOut_payload_0_14010 = (_zz_dataOut_payload_0_14008 ? _zz_dataOut_payload_0_11863 : _zz_dataOut_payload_0_11816);
  assign _zz_dataOut_payload_0_14011 = (_zz_dataOut_payload_0_11817 < _zz_dataOut_payload_0_11862);
  assign _zz_dataOut_payload_0_14012 = (_zz_dataOut_payload_0_14011 ? _zz_dataOut_payload_0_11817 : _zz_dataOut_payload_0_11862);
  assign _zz_dataOut_payload_0_14013 = (_zz_dataOut_payload_0_14011 ? _zz_dataOut_payload_0_11862 : _zz_dataOut_payload_0_11817);
  assign _zz_dataOut_payload_0_14014 = (_zz_dataOut_payload_0_11818 < _zz_dataOut_payload_0_11861);
  assign _zz_dataOut_payload_0_14015 = (_zz_dataOut_payload_0_14014 ? _zz_dataOut_payload_0_11818 : _zz_dataOut_payload_0_11861);
  assign _zz_dataOut_payload_0_14016 = (_zz_dataOut_payload_0_14014 ? _zz_dataOut_payload_0_11861 : _zz_dataOut_payload_0_11818);
  assign _zz_dataOut_payload_0_14017 = (_zz_dataOut_payload_0_11819 < _zz_dataOut_payload_0_11860);
  assign _zz_dataOut_payload_0_14018 = (_zz_dataOut_payload_0_14017 ? _zz_dataOut_payload_0_11819 : _zz_dataOut_payload_0_11860);
  assign _zz_dataOut_payload_0_14019 = (_zz_dataOut_payload_0_14017 ? _zz_dataOut_payload_0_11860 : _zz_dataOut_payload_0_11819);
  assign _zz_dataOut_payload_0_14020 = (_zz_dataOut_payload_0_11820 < _zz_dataOut_payload_0_11859);
  assign _zz_dataOut_payload_0_14021 = (_zz_dataOut_payload_0_14020 ? _zz_dataOut_payload_0_11820 : _zz_dataOut_payload_0_11859);
  assign _zz_dataOut_payload_0_14022 = (_zz_dataOut_payload_0_14020 ? _zz_dataOut_payload_0_11859 : _zz_dataOut_payload_0_11820);
  assign _zz_dataOut_payload_0_14023 = (_zz_dataOut_payload_0_11821 < _zz_dataOut_payload_0_11858);
  assign _zz_dataOut_payload_0_14024 = (_zz_dataOut_payload_0_14023 ? _zz_dataOut_payload_0_11821 : _zz_dataOut_payload_0_11858);
  assign _zz_dataOut_payload_0_14025 = (_zz_dataOut_payload_0_14023 ? _zz_dataOut_payload_0_11858 : _zz_dataOut_payload_0_11821);
  assign _zz_dataOut_payload_0_14026 = (_zz_dataOut_payload_0_11822 < _zz_dataOut_payload_0_11857);
  assign _zz_dataOut_payload_0_14027 = (_zz_dataOut_payload_0_14026 ? _zz_dataOut_payload_0_11822 : _zz_dataOut_payload_0_11857);
  assign _zz_dataOut_payload_0_14028 = (_zz_dataOut_payload_0_14026 ? _zz_dataOut_payload_0_11857 : _zz_dataOut_payload_0_11822);
  assign _zz_dataOut_payload_0_14029 = (_zz_dataOut_payload_0_11823 < _zz_dataOut_payload_0_11856);
  assign _zz_dataOut_payload_0_14030 = (_zz_dataOut_payload_0_14029 ? _zz_dataOut_payload_0_11823 : _zz_dataOut_payload_0_11856);
  assign _zz_dataOut_payload_0_14031 = (_zz_dataOut_payload_0_14029 ? _zz_dataOut_payload_0_11856 : _zz_dataOut_payload_0_11823);
  assign _zz_dataOut_payload_0_14032 = (_zz_dataOut_payload_0_11824 < _zz_dataOut_payload_0_11855);
  assign _zz_dataOut_payload_0_14033 = (_zz_dataOut_payload_0_14032 ? _zz_dataOut_payload_0_11824 : _zz_dataOut_payload_0_11855);
  assign _zz_dataOut_payload_0_14034 = (_zz_dataOut_payload_0_14032 ? _zz_dataOut_payload_0_11855 : _zz_dataOut_payload_0_11824);
  assign _zz_dataOut_payload_0_14035 = (_zz_dataOut_payload_0_11825 < _zz_dataOut_payload_0_11854);
  assign _zz_dataOut_payload_0_14036 = (_zz_dataOut_payload_0_14035 ? _zz_dataOut_payload_0_11825 : _zz_dataOut_payload_0_11854);
  assign _zz_dataOut_payload_0_14037 = (_zz_dataOut_payload_0_14035 ? _zz_dataOut_payload_0_11854 : _zz_dataOut_payload_0_11825);
  assign _zz_dataOut_payload_0_14038 = (_zz_dataOut_payload_0_11826 < _zz_dataOut_payload_0_11853);
  assign _zz_dataOut_payload_0_14039 = (_zz_dataOut_payload_0_14038 ? _zz_dataOut_payload_0_11826 : _zz_dataOut_payload_0_11853);
  assign _zz_dataOut_payload_0_14040 = (_zz_dataOut_payload_0_14038 ? _zz_dataOut_payload_0_11853 : _zz_dataOut_payload_0_11826);
  assign _zz_dataOut_payload_0_14041 = (_zz_dataOut_payload_0_11827 < _zz_dataOut_payload_0_11852);
  assign _zz_dataOut_payload_0_14042 = (_zz_dataOut_payload_0_14041 ? _zz_dataOut_payload_0_11827 : _zz_dataOut_payload_0_11852);
  assign _zz_dataOut_payload_0_14043 = (_zz_dataOut_payload_0_14041 ? _zz_dataOut_payload_0_11852 : _zz_dataOut_payload_0_11827);
  assign _zz_dataOut_payload_0_14044 = (_zz_dataOut_payload_0_11828 < _zz_dataOut_payload_0_11851);
  assign _zz_dataOut_payload_0_14045 = (_zz_dataOut_payload_0_14044 ? _zz_dataOut_payload_0_11828 : _zz_dataOut_payload_0_11851);
  assign _zz_dataOut_payload_0_14046 = (_zz_dataOut_payload_0_14044 ? _zz_dataOut_payload_0_11851 : _zz_dataOut_payload_0_11828);
  assign _zz_dataOut_payload_0_14047 = (_zz_dataOut_payload_0_11829 < _zz_dataOut_payload_0_11850);
  assign _zz_dataOut_payload_0_14048 = (_zz_dataOut_payload_0_14047 ? _zz_dataOut_payload_0_11829 : _zz_dataOut_payload_0_11850);
  assign _zz_dataOut_payload_0_14049 = (_zz_dataOut_payload_0_14047 ? _zz_dataOut_payload_0_11850 : _zz_dataOut_payload_0_11829);
  assign _zz_dataOut_payload_0_14050 = (_zz_dataOut_payload_0_11830 < _zz_dataOut_payload_0_11849);
  assign _zz_dataOut_payload_0_14051 = (_zz_dataOut_payload_0_14050 ? _zz_dataOut_payload_0_11830 : _zz_dataOut_payload_0_11849);
  assign _zz_dataOut_payload_0_14052 = (_zz_dataOut_payload_0_14050 ? _zz_dataOut_payload_0_11849 : _zz_dataOut_payload_0_11830);
  assign _zz_dataOut_payload_0_14053 = (_zz_dataOut_payload_0_11831 < _zz_dataOut_payload_0_11848);
  assign _zz_dataOut_payload_0_14054 = (_zz_dataOut_payload_0_14053 ? _zz_dataOut_payload_0_11831 : _zz_dataOut_payload_0_11848);
  assign _zz_dataOut_payload_0_14055 = (_zz_dataOut_payload_0_14053 ? _zz_dataOut_payload_0_11848 : _zz_dataOut_payload_0_11831);
  assign _zz_dataOut_payload_0_14056 = (_zz_dataOut_payload_0_11832 < _zz_dataOut_payload_0_11847);
  assign _zz_dataOut_payload_0_14057 = (_zz_dataOut_payload_0_14056 ? _zz_dataOut_payload_0_11832 : _zz_dataOut_payload_0_11847);
  assign _zz_dataOut_payload_0_14058 = (_zz_dataOut_payload_0_14056 ? _zz_dataOut_payload_0_11847 : _zz_dataOut_payload_0_11832);
  assign _zz_dataOut_payload_0_14059 = (_zz_dataOut_payload_0_11833 < _zz_dataOut_payload_0_11846);
  assign _zz_dataOut_payload_0_14060 = (_zz_dataOut_payload_0_14059 ? _zz_dataOut_payload_0_11833 : _zz_dataOut_payload_0_11846);
  assign _zz_dataOut_payload_0_14061 = (_zz_dataOut_payload_0_14059 ? _zz_dataOut_payload_0_11846 : _zz_dataOut_payload_0_11833);
  assign _zz_dataOut_payload_0_14062 = (_zz_dataOut_payload_0_11834 < _zz_dataOut_payload_0_11845);
  assign _zz_dataOut_payload_0_14063 = (_zz_dataOut_payload_0_14062 ? _zz_dataOut_payload_0_11834 : _zz_dataOut_payload_0_11845);
  assign _zz_dataOut_payload_0_14064 = (_zz_dataOut_payload_0_14062 ? _zz_dataOut_payload_0_11845 : _zz_dataOut_payload_0_11834);
  assign _zz_dataOut_payload_0_14065 = (_zz_dataOut_payload_0_11835 < _zz_dataOut_payload_0_11844);
  assign _zz_dataOut_payload_0_14066 = (_zz_dataOut_payload_0_14065 ? _zz_dataOut_payload_0_11835 : _zz_dataOut_payload_0_11844);
  assign _zz_dataOut_payload_0_14067 = (_zz_dataOut_payload_0_14065 ? _zz_dataOut_payload_0_11844 : _zz_dataOut_payload_0_11835);
  assign _zz_dataOut_payload_0_14068 = (_zz_dataOut_payload_0_11836 < _zz_dataOut_payload_0_11843);
  assign _zz_dataOut_payload_0_14069 = (_zz_dataOut_payload_0_14068 ? _zz_dataOut_payload_0_11836 : _zz_dataOut_payload_0_11843);
  assign _zz_dataOut_payload_0_14070 = (_zz_dataOut_payload_0_14068 ? _zz_dataOut_payload_0_11843 : _zz_dataOut_payload_0_11836);
  assign _zz_dataOut_payload_0_14071 = (_zz_dataOut_payload_0_11837 < _zz_dataOut_payload_0_11842);
  assign _zz_dataOut_payload_0_14072 = (_zz_dataOut_payload_0_14071 ? _zz_dataOut_payload_0_11837 : _zz_dataOut_payload_0_11842);
  assign _zz_dataOut_payload_0_14073 = (_zz_dataOut_payload_0_14071 ? _zz_dataOut_payload_0_11842 : _zz_dataOut_payload_0_11837);
  assign _zz_dataOut_payload_0_14074 = (_zz_dataOut_payload_0_11838 < _zz_dataOut_payload_0_11841);
  assign _zz_dataOut_payload_0_14075 = (_zz_dataOut_payload_0_14074 ? _zz_dataOut_payload_0_11838 : _zz_dataOut_payload_0_11841);
  assign _zz_dataOut_payload_0_14076 = (_zz_dataOut_payload_0_14074 ? _zz_dataOut_payload_0_11841 : _zz_dataOut_payload_0_11838);
  assign _zz_dataOut_payload_0_14077 = (_zz_dataOut_payload_0_11839 < _zz_dataOut_payload_0_11840);
  assign _zz_dataOut_payload_0_14078 = (_zz_dataOut_payload_0_14077 ? _zz_dataOut_payload_0_11839 : _zz_dataOut_payload_0_11840);
  assign _zz_dataOut_payload_0_14079 = (_zz_dataOut_payload_0_14077 ? _zz_dataOut_payload_0_11840 : _zz_dataOut_payload_0_11839);
  assign _zz_dataOut_payload_0_14080 = (_zz_dataOut_payload_0_13889 < _zz_dataOut_payload_0_13985);
  assign _zz_dataOut_payload_0_14081 = (_zz_dataOut_payload_0_14080 ? _zz_dataOut_payload_0_13889 : _zz_dataOut_payload_0_13985);
  assign _zz_dataOut_payload_0_14082 = (_zz_dataOut_payload_0_14080 ? _zz_dataOut_payload_0_13985 : _zz_dataOut_payload_0_13889);
  assign _zz_dataOut_payload_0_14083 = (_zz_dataOut_payload_0_13892 < _zz_dataOut_payload_0_13988);
  assign _zz_dataOut_payload_0_14084 = (_zz_dataOut_payload_0_14083 ? _zz_dataOut_payload_0_13892 : _zz_dataOut_payload_0_13988);
  assign _zz_dataOut_payload_0_14085 = (_zz_dataOut_payload_0_14083 ? _zz_dataOut_payload_0_13988 : _zz_dataOut_payload_0_13892);
  assign _zz_dataOut_payload_0_14086 = (_zz_dataOut_payload_0_13895 < _zz_dataOut_payload_0_13991);
  assign _zz_dataOut_payload_0_14087 = (_zz_dataOut_payload_0_14086 ? _zz_dataOut_payload_0_13895 : _zz_dataOut_payload_0_13991);
  assign _zz_dataOut_payload_0_14088 = (_zz_dataOut_payload_0_14086 ? _zz_dataOut_payload_0_13991 : _zz_dataOut_payload_0_13895);
  assign _zz_dataOut_payload_0_14089 = (_zz_dataOut_payload_0_13898 < _zz_dataOut_payload_0_13994);
  assign _zz_dataOut_payload_0_14090 = (_zz_dataOut_payload_0_14089 ? _zz_dataOut_payload_0_13898 : _zz_dataOut_payload_0_13994);
  assign _zz_dataOut_payload_0_14091 = (_zz_dataOut_payload_0_14089 ? _zz_dataOut_payload_0_13994 : _zz_dataOut_payload_0_13898);
  assign _zz_dataOut_payload_0_14092 = (_zz_dataOut_payload_0_13901 < _zz_dataOut_payload_0_13997);
  assign _zz_dataOut_payload_0_14093 = (_zz_dataOut_payload_0_14092 ? _zz_dataOut_payload_0_13901 : _zz_dataOut_payload_0_13997);
  assign _zz_dataOut_payload_0_14094 = (_zz_dataOut_payload_0_14092 ? _zz_dataOut_payload_0_13997 : _zz_dataOut_payload_0_13901);
  assign _zz_dataOut_payload_0_14095 = (_zz_dataOut_payload_0_13904 < _zz_dataOut_payload_0_14000);
  assign _zz_dataOut_payload_0_14096 = (_zz_dataOut_payload_0_14095 ? _zz_dataOut_payload_0_13904 : _zz_dataOut_payload_0_14000);
  assign _zz_dataOut_payload_0_14097 = (_zz_dataOut_payload_0_14095 ? _zz_dataOut_payload_0_14000 : _zz_dataOut_payload_0_13904);
  assign _zz_dataOut_payload_0_14098 = (_zz_dataOut_payload_0_13907 < _zz_dataOut_payload_0_14003);
  assign _zz_dataOut_payload_0_14099 = (_zz_dataOut_payload_0_14098 ? _zz_dataOut_payload_0_13907 : _zz_dataOut_payload_0_14003);
  assign _zz_dataOut_payload_0_14100 = (_zz_dataOut_payload_0_14098 ? _zz_dataOut_payload_0_14003 : _zz_dataOut_payload_0_13907);
  assign _zz_dataOut_payload_0_14101 = (_zz_dataOut_payload_0_13910 < _zz_dataOut_payload_0_14006);
  assign _zz_dataOut_payload_0_14102 = (_zz_dataOut_payload_0_14101 ? _zz_dataOut_payload_0_13910 : _zz_dataOut_payload_0_14006);
  assign _zz_dataOut_payload_0_14103 = (_zz_dataOut_payload_0_14101 ? _zz_dataOut_payload_0_14006 : _zz_dataOut_payload_0_13910);
  assign _zz_dataOut_payload_0_14104 = (_zz_dataOut_payload_0_13913 < _zz_dataOut_payload_0_14009);
  assign _zz_dataOut_payload_0_14105 = (_zz_dataOut_payload_0_14104 ? _zz_dataOut_payload_0_13913 : _zz_dataOut_payload_0_14009);
  assign _zz_dataOut_payload_0_14106 = (_zz_dataOut_payload_0_14104 ? _zz_dataOut_payload_0_14009 : _zz_dataOut_payload_0_13913);
  assign _zz_dataOut_payload_0_14107 = (_zz_dataOut_payload_0_13916 < _zz_dataOut_payload_0_14012);
  assign _zz_dataOut_payload_0_14108 = (_zz_dataOut_payload_0_14107 ? _zz_dataOut_payload_0_13916 : _zz_dataOut_payload_0_14012);
  assign _zz_dataOut_payload_0_14109 = (_zz_dataOut_payload_0_14107 ? _zz_dataOut_payload_0_14012 : _zz_dataOut_payload_0_13916);
  assign _zz_dataOut_payload_0_14110 = (_zz_dataOut_payload_0_13919 < _zz_dataOut_payload_0_14015);
  assign _zz_dataOut_payload_0_14111 = (_zz_dataOut_payload_0_14110 ? _zz_dataOut_payload_0_13919 : _zz_dataOut_payload_0_14015);
  assign _zz_dataOut_payload_0_14112 = (_zz_dataOut_payload_0_14110 ? _zz_dataOut_payload_0_14015 : _zz_dataOut_payload_0_13919);
  assign _zz_dataOut_payload_0_14113 = (_zz_dataOut_payload_0_13922 < _zz_dataOut_payload_0_14018);
  assign _zz_dataOut_payload_0_14114 = (_zz_dataOut_payload_0_14113 ? _zz_dataOut_payload_0_13922 : _zz_dataOut_payload_0_14018);
  assign _zz_dataOut_payload_0_14115 = (_zz_dataOut_payload_0_14113 ? _zz_dataOut_payload_0_14018 : _zz_dataOut_payload_0_13922);
  assign _zz_dataOut_payload_0_14116 = (_zz_dataOut_payload_0_13925 < _zz_dataOut_payload_0_14021);
  assign _zz_dataOut_payload_0_14117 = (_zz_dataOut_payload_0_14116 ? _zz_dataOut_payload_0_13925 : _zz_dataOut_payload_0_14021);
  assign _zz_dataOut_payload_0_14118 = (_zz_dataOut_payload_0_14116 ? _zz_dataOut_payload_0_14021 : _zz_dataOut_payload_0_13925);
  assign _zz_dataOut_payload_0_14119 = (_zz_dataOut_payload_0_13928 < _zz_dataOut_payload_0_14024);
  assign _zz_dataOut_payload_0_14120 = (_zz_dataOut_payload_0_14119 ? _zz_dataOut_payload_0_13928 : _zz_dataOut_payload_0_14024);
  assign _zz_dataOut_payload_0_14121 = (_zz_dataOut_payload_0_14119 ? _zz_dataOut_payload_0_14024 : _zz_dataOut_payload_0_13928);
  assign _zz_dataOut_payload_0_14122 = (_zz_dataOut_payload_0_13931 < _zz_dataOut_payload_0_14027);
  assign _zz_dataOut_payload_0_14123 = (_zz_dataOut_payload_0_14122 ? _zz_dataOut_payload_0_13931 : _zz_dataOut_payload_0_14027);
  assign _zz_dataOut_payload_0_14124 = (_zz_dataOut_payload_0_14122 ? _zz_dataOut_payload_0_14027 : _zz_dataOut_payload_0_13931);
  assign _zz_dataOut_payload_0_14125 = (_zz_dataOut_payload_0_13934 < _zz_dataOut_payload_0_14030);
  assign _zz_dataOut_payload_0_14126 = (_zz_dataOut_payload_0_14125 ? _zz_dataOut_payload_0_13934 : _zz_dataOut_payload_0_14030);
  assign _zz_dataOut_payload_0_14127 = (_zz_dataOut_payload_0_14125 ? _zz_dataOut_payload_0_14030 : _zz_dataOut_payload_0_13934);
  assign _zz_dataOut_payload_0_14128 = (_zz_dataOut_payload_0_13937 < _zz_dataOut_payload_0_14033);
  assign _zz_dataOut_payload_0_14129 = (_zz_dataOut_payload_0_14128 ? _zz_dataOut_payload_0_13937 : _zz_dataOut_payload_0_14033);
  assign _zz_dataOut_payload_0_14130 = (_zz_dataOut_payload_0_14128 ? _zz_dataOut_payload_0_14033 : _zz_dataOut_payload_0_13937);
  assign _zz_dataOut_payload_0_14131 = (_zz_dataOut_payload_0_13940 < _zz_dataOut_payload_0_14036);
  assign _zz_dataOut_payload_0_14132 = (_zz_dataOut_payload_0_14131 ? _zz_dataOut_payload_0_13940 : _zz_dataOut_payload_0_14036);
  assign _zz_dataOut_payload_0_14133 = (_zz_dataOut_payload_0_14131 ? _zz_dataOut_payload_0_14036 : _zz_dataOut_payload_0_13940);
  assign _zz_dataOut_payload_0_14134 = (_zz_dataOut_payload_0_13943 < _zz_dataOut_payload_0_14039);
  assign _zz_dataOut_payload_0_14135 = (_zz_dataOut_payload_0_14134 ? _zz_dataOut_payload_0_13943 : _zz_dataOut_payload_0_14039);
  assign _zz_dataOut_payload_0_14136 = (_zz_dataOut_payload_0_14134 ? _zz_dataOut_payload_0_14039 : _zz_dataOut_payload_0_13943);
  assign _zz_dataOut_payload_0_14137 = (_zz_dataOut_payload_0_13946 < _zz_dataOut_payload_0_14042);
  assign _zz_dataOut_payload_0_14138 = (_zz_dataOut_payload_0_14137 ? _zz_dataOut_payload_0_13946 : _zz_dataOut_payload_0_14042);
  assign _zz_dataOut_payload_0_14139 = (_zz_dataOut_payload_0_14137 ? _zz_dataOut_payload_0_14042 : _zz_dataOut_payload_0_13946);
  assign _zz_dataOut_payload_0_14140 = (_zz_dataOut_payload_0_13949 < _zz_dataOut_payload_0_14045);
  assign _zz_dataOut_payload_0_14141 = (_zz_dataOut_payload_0_14140 ? _zz_dataOut_payload_0_13949 : _zz_dataOut_payload_0_14045);
  assign _zz_dataOut_payload_0_14142 = (_zz_dataOut_payload_0_14140 ? _zz_dataOut_payload_0_14045 : _zz_dataOut_payload_0_13949);
  assign _zz_dataOut_payload_0_14143 = (_zz_dataOut_payload_0_13952 < _zz_dataOut_payload_0_14048);
  assign _zz_dataOut_payload_0_14144 = (_zz_dataOut_payload_0_14143 ? _zz_dataOut_payload_0_13952 : _zz_dataOut_payload_0_14048);
  assign _zz_dataOut_payload_0_14145 = (_zz_dataOut_payload_0_14143 ? _zz_dataOut_payload_0_14048 : _zz_dataOut_payload_0_13952);
  assign _zz_dataOut_payload_0_14146 = (_zz_dataOut_payload_0_13955 < _zz_dataOut_payload_0_14051);
  assign _zz_dataOut_payload_0_14147 = (_zz_dataOut_payload_0_14146 ? _zz_dataOut_payload_0_13955 : _zz_dataOut_payload_0_14051);
  assign _zz_dataOut_payload_0_14148 = (_zz_dataOut_payload_0_14146 ? _zz_dataOut_payload_0_14051 : _zz_dataOut_payload_0_13955);
  assign _zz_dataOut_payload_0_14149 = (_zz_dataOut_payload_0_13958 < _zz_dataOut_payload_0_14054);
  assign _zz_dataOut_payload_0_14150 = (_zz_dataOut_payload_0_14149 ? _zz_dataOut_payload_0_13958 : _zz_dataOut_payload_0_14054);
  assign _zz_dataOut_payload_0_14151 = (_zz_dataOut_payload_0_14149 ? _zz_dataOut_payload_0_14054 : _zz_dataOut_payload_0_13958);
  assign _zz_dataOut_payload_0_14152 = (_zz_dataOut_payload_0_13961 < _zz_dataOut_payload_0_14057);
  assign _zz_dataOut_payload_0_14153 = (_zz_dataOut_payload_0_14152 ? _zz_dataOut_payload_0_13961 : _zz_dataOut_payload_0_14057);
  assign _zz_dataOut_payload_0_14154 = (_zz_dataOut_payload_0_14152 ? _zz_dataOut_payload_0_14057 : _zz_dataOut_payload_0_13961);
  assign _zz_dataOut_payload_0_14155 = (_zz_dataOut_payload_0_13964 < _zz_dataOut_payload_0_14060);
  assign _zz_dataOut_payload_0_14156 = (_zz_dataOut_payload_0_14155 ? _zz_dataOut_payload_0_13964 : _zz_dataOut_payload_0_14060);
  assign _zz_dataOut_payload_0_14157 = (_zz_dataOut_payload_0_14155 ? _zz_dataOut_payload_0_14060 : _zz_dataOut_payload_0_13964);
  assign _zz_dataOut_payload_0_14158 = (_zz_dataOut_payload_0_13967 < _zz_dataOut_payload_0_14063);
  assign _zz_dataOut_payload_0_14159 = (_zz_dataOut_payload_0_14158 ? _zz_dataOut_payload_0_13967 : _zz_dataOut_payload_0_14063);
  assign _zz_dataOut_payload_0_14160 = (_zz_dataOut_payload_0_14158 ? _zz_dataOut_payload_0_14063 : _zz_dataOut_payload_0_13967);
  assign _zz_dataOut_payload_0_14161 = (_zz_dataOut_payload_0_13970 < _zz_dataOut_payload_0_14066);
  assign _zz_dataOut_payload_0_14162 = (_zz_dataOut_payload_0_14161 ? _zz_dataOut_payload_0_13970 : _zz_dataOut_payload_0_14066);
  assign _zz_dataOut_payload_0_14163 = (_zz_dataOut_payload_0_14161 ? _zz_dataOut_payload_0_14066 : _zz_dataOut_payload_0_13970);
  assign _zz_dataOut_payload_0_14164 = (_zz_dataOut_payload_0_13973 < _zz_dataOut_payload_0_14069);
  assign _zz_dataOut_payload_0_14165 = (_zz_dataOut_payload_0_14164 ? _zz_dataOut_payload_0_13973 : _zz_dataOut_payload_0_14069);
  assign _zz_dataOut_payload_0_14166 = (_zz_dataOut_payload_0_14164 ? _zz_dataOut_payload_0_14069 : _zz_dataOut_payload_0_13973);
  assign _zz_dataOut_payload_0_14167 = (_zz_dataOut_payload_0_13976 < _zz_dataOut_payload_0_14072);
  assign _zz_dataOut_payload_0_14168 = (_zz_dataOut_payload_0_14167 ? _zz_dataOut_payload_0_13976 : _zz_dataOut_payload_0_14072);
  assign _zz_dataOut_payload_0_14169 = (_zz_dataOut_payload_0_14167 ? _zz_dataOut_payload_0_14072 : _zz_dataOut_payload_0_13976);
  assign _zz_dataOut_payload_0_14170 = (_zz_dataOut_payload_0_13979 < _zz_dataOut_payload_0_14075);
  assign _zz_dataOut_payload_0_14171 = (_zz_dataOut_payload_0_14170 ? _zz_dataOut_payload_0_13979 : _zz_dataOut_payload_0_14075);
  assign _zz_dataOut_payload_0_14172 = (_zz_dataOut_payload_0_14170 ? _zz_dataOut_payload_0_14075 : _zz_dataOut_payload_0_13979);
  assign _zz_dataOut_payload_0_14173 = (_zz_dataOut_payload_0_13982 < _zz_dataOut_payload_0_14078);
  assign _zz_dataOut_payload_0_14174 = (_zz_dataOut_payload_0_14173 ? _zz_dataOut_payload_0_13982 : _zz_dataOut_payload_0_14078);
  assign _zz_dataOut_payload_0_14175 = (_zz_dataOut_payload_0_14173 ? _zz_dataOut_payload_0_14078 : _zz_dataOut_payload_0_13982);
  assign _zz_dataOut_payload_0_14176 = (_zz_dataOut_payload_0_14081 < _zz_dataOut_payload_0_14129);
  assign _zz_dataOut_payload_0_14177 = (_zz_dataOut_payload_0_14176 ? _zz_dataOut_payload_0_14081 : _zz_dataOut_payload_0_14129);
  assign _zz_dataOut_payload_0_14178 = (_zz_dataOut_payload_0_14176 ? _zz_dataOut_payload_0_14129 : _zz_dataOut_payload_0_14081);
  assign _zz_dataOut_payload_0_14179 = (_zz_dataOut_payload_0_14084 < _zz_dataOut_payload_0_14132);
  assign _zz_dataOut_payload_0_14180 = (_zz_dataOut_payload_0_14179 ? _zz_dataOut_payload_0_14084 : _zz_dataOut_payload_0_14132);
  assign _zz_dataOut_payload_0_14181 = (_zz_dataOut_payload_0_14179 ? _zz_dataOut_payload_0_14132 : _zz_dataOut_payload_0_14084);
  assign _zz_dataOut_payload_0_14182 = (_zz_dataOut_payload_0_14087 < _zz_dataOut_payload_0_14135);
  assign _zz_dataOut_payload_0_14183 = (_zz_dataOut_payload_0_14182 ? _zz_dataOut_payload_0_14087 : _zz_dataOut_payload_0_14135);
  assign _zz_dataOut_payload_0_14184 = (_zz_dataOut_payload_0_14182 ? _zz_dataOut_payload_0_14135 : _zz_dataOut_payload_0_14087);
  assign _zz_dataOut_payload_0_14185 = (_zz_dataOut_payload_0_14090 < _zz_dataOut_payload_0_14138);
  assign _zz_dataOut_payload_0_14186 = (_zz_dataOut_payload_0_14185 ? _zz_dataOut_payload_0_14090 : _zz_dataOut_payload_0_14138);
  assign _zz_dataOut_payload_0_14187 = (_zz_dataOut_payload_0_14185 ? _zz_dataOut_payload_0_14138 : _zz_dataOut_payload_0_14090);
  assign _zz_dataOut_payload_0_14188 = (_zz_dataOut_payload_0_14093 < _zz_dataOut_payload_0_14141);
  assign _zz_dataOut_payload_0_14189 = (_zz_dataOut_payload_0_14188 ? _zz_dataOut_payload_0_14093 : _zz_dataOut_payload_0_14141);
  assign _zz_dataOut_payload_0_14190 = (_zz_dataOut_payload_0_14188 ? _zz_dataOut_payload_0_14141 : _zz_dataOut_payload_0_14093);
  assign _zz_dataOut_payload_0_14191 = (_zz_dataOut_payload_0_14096 < _zz_dataOut_payload_0_14144);
  assign _zz_dataOut_payload_0_14192 = (_zz_dataOut_payload_0_14191 ? _zz_dataOut_payload_0_14096 : _zz_dataOut_payload_0_14144);
  assign _zz_dataOut_payload_0_14193 = (_zz_dataOut_payload_0_14191 ? _zz_dataOut_payload_0_14144 : _zz_dataOut_payload_0_14096);
  assign _zz_dataOut_payload_0_14194 = (_zz_dataOut_payload_0_14099 < _zz_dataOut_payload_0_14147);
  assign _zz_dataOut_payload_0_14195 = (_zz_dataOut_payload_0_14194 ? _zz_dataOut_payload_0_14099 : _zz_dataOut_payload_0_14147);
  assign _zz_dataOut_payload_0_14196 = (_zz_dataOut_payload_0_14194 ? _zz_dataOut_payload_0_14147 : _zz_dataOut_payload_0_14099);
  assign _zz_dataOut_payload_0_14197 = (_zz_dataOut_payload_0_14102 < _zz_dataOut_payload_0_14150);
  assign _zz_dataOut_payload_0_14198 = (_zz_dataOut_payload_0_14197 ? _zz_dataOut_payload_0_14102 : _zz_dataOut_payload_0_14150);
  assign _zz_dataOut_payload_0_14199 = (_zz_dataOut_payload_0_14197 ? _zz_dataOut_payload_0_14150 : _zz_dataOut_payload_0_14102);
  assign _zz_dataOut_payload_0_14200 = (_zz_dataOut_payload_0_14105 < _zz_dataOut_payload_0_14153);
  assign _zz_dataOut_payload_0_14201 = (_zz_dataOut_payload_0_14200 ? _zz_dataOut_payload_0_14105 : _zz_dataOut_payload_0_14153);
  assign _zz_dataOut_payload_0_14202 = (_zz_dataOut_payload_0_14200 ? _zz_dataOut_payload_0_14153 : _zz_dataOut_payload_0_14105);
  assign _zz_dataOut_payload_0_14203 = (_zz_dataOut_payload_0_14108 < _zz_dataOut_payload_0_14156);
  assign _zz_dataOut_payload_0_14204 = (_zz_dataOut_payload_0_14203 ? _zz_dataOut_payload_0_14108 : _zz_dataOut_payload_0_14156);
  assign _zz_dataOut_payload_0_14205 = (_zz_dataOut_payload_0_14203 ? _zz_dataOut_payload_0_14156 : _zz_dataOut_payload_0_14108);
  assign _zz_dataOut_payload_0_14206 = (_zz_dataOut_payload_0_14111 < _zz_dataOut_payload_0_14159);
  assign _zz_dataOut_payload_0_14207 = (_zz_dataOut_payload_0_14206 ? _zz_dataOut_payload_0_14111 : _zz_dataOut_payload_0_14159);
  assign _zz_dataOut_payload_0_14208 = (_zz_dataOut_payload_0_14206 ? _zz_dataOut_payload_0_14159 : _zz_dataOut_payload_0_14111);
  assign _zz_dataOut_payload_0_14209 = (_zz_dataOut_payload_0_14114 < _zz_dataOut_payload_0_14162);
  assign _zz_dataOut_payload_0_14210 = (_zz_dataOut_payload_0_14209 ? _zz_dataOut_payload_0_14114 : _zz_dataOut_payload_0_14162);
  assign _zz_dataOut_payload_0_14211 = (_zz_dataOut_payload_0_14209 ? _zz_dataOut_payload_0_14162 : _zz_dataOut_payload_0_14114);
  assign _zz_dataOut_payload_0_14212 = (_zz_dataOut_payload_0_14117 < _zz_dataOut_payload_0_14165);
  assign _zz_dataOut_payload_0_14213 = (_zz_dataOut_payload_0_14212 ? _zz_dataOut_payload_0_14117 : _zz_dataOut_payload_0_14165);
  assign _zz_dataOut_payload_0_14214 = (_zz_dataOut_payload_0_14212 ? _zz_dataOut_payload_0_14165 : _zz_dataOut_payload_0_14117);
  assign _zz_dataOut_payload_0_14215 = (_zz_dataOut_payload_0_14120 < _zz_dataOut_payload_0_14168);
  assign _zz_dataOut_payload_0_14216 = (_zz_dataOut_payload_0_14215 ? _zz_dataOut_payload_0_14120 : _zz_dataOut_payload_0_14168);
  assign _zz_dataOut_payload_0_14217 = (_zz_dataOut_payload_0_14215 ? _zz_dataOut_payload_0_14168 : _zz_dataOut_payload_0_14120);
  assign _zz_dataOut_payload_0_14218 = (_zz_dataOut_payload_0_14123 < _zz_dataOut_payload_0_14171);
  assign _zz_dataOut_payload_0_14219 = (_zz_dataOut_payload_0_14218 ? _zz_dataOut_payload_0_14123 : _zz_dataOut_payload_0_14171);
  assign _zz_dataOut_payload_0_14220 = (_zz_dataOut_payload_0_14218 ? _zz_dataOut_payload_0_14171 : _zz_dataOut_payload_0_14123);
  assign _zz_dataOut_payload_0_14221 = (_zz_dataOut_payload_0_14126 < _zz_dataOut_payload_0_14174);
  assign _zz_dataOut_payload_0_14222 = (_zz_dataOut_payload_0_14221 ? _zz_dataOut_payload_0_14126 : _zz_dataOut_payload_0_14174);
  assign _zz_dataOut_payload_0_14223 = (_zz_dataOut_payload_0_14221 ? _zz_dataOut_payload_0_14174 : _zz_dataOut_payload_0_14126);
  assign _zz_dataOut_payload_0_14224 = (_zz_dataOut_payload_0_14177 < _zz_dataOut_payload_0_14201);
  assign _zz_dataOut_payload_0_14225 = (_zz_dataOut_payload_0_14224 ? _zz_dataOut_payload_0_14177 : _zz_dataOut_payload_0_14201);
  assign _zz_dataOut_payload_0_14226 = (_zz_dataOut_payload_0_14224 ? _zz_dataOut_payload_0_14201 : _zz_dataOut_payload_0_14177);
  assign _zz_dataOut_payload_0_14227 = (_zz_dataOut_payload_0_14180 < _zz_dataOut_payload_0_14204);
  assign _zz_dataOut_payload_0_14228 = (_zz_dataOut_payload_0_14227 ? _zz_dataOut_payload_0_14180 : _zz_dataOut_payload_0_14204);
  assign _zz_dataOut_payload_0_14229 = (_zz_dataOut_payload_0_14227 ? _zz_dataOut_payload_0_14204 : _zz_dataOut_payload_0_14180);
  assign _zz_dataOut_payload_0_14230 = (_zz_dataOut_payload_0_14183 < _zz_dataOut_payload_0_14207);
  assign _zz_dataOut_payload_0_14231 = (_zz_dataOut_payload_0_14230 ? _zz_dataOut_payload_0_14183 : _zz_dataOut_payload_0_14207);
  assign _zz_dataOut_payload_0_14232 = (_zz_dataOut_payload_0_14230 ? _zz_dataOut_payload_0_14207 : _zz_dataOut_payload_0_14183);
  assign _zz_dataOut_payload_0_14233 = (_zz_dataOut_payload_0_14186 < _zz_dataOut_payload_0_14210);
  assign _zz_dataOut_payload_0_14234 = (_zz_dataOut_payload_0_14233 ? _zz_dataOut_payload_0_14186 : _zz_dataOut_payload_0_14210);
  assign _zz_dataOut_payload_0_14235 = (_zz_dataOut_payload_0_14233 ? _zz_dataOut_payload_0_14210 : _zz_dataOut_payload_0_14186);
  assign _zz_dataOut_payload_0_14236 = (_zz_dataOut_payload_0_14189 < _zz_dataOut_payload_0_14213);
  assign _zz_dataOut_payload_0_14237 = (_zz_dataOut_payload_0_14236 ? _zz_dataOut_payload_0_14189 : _zz_dataOut_payload_0_14213);
  assign _zz_dataOut_payload_0_14238 = (_zz_dataOut_payload_0_14236 ? _zz_dataOut_payload_0_14213 : _zz_dataOut_payload_0_14189);
  assign _zz_dataOut_payload_0_14239 = (_zz_dataOut_payload_0_14192 < _zz_dataOut_payload_0_14216);
  assign _zz_dataOut_payload_0_14240 = (_zz_dataOut_payload_0_14239 ? _zz_dataOut_payload_0_14192 : _zz_dataOut_payload_0_14216);
  assign _zz_dataOut_payload_0_14241 = (_zz_dataOut_payload_0_14239 ? _zz_dataOut_payload_0_14216 : _zz_dataOut_payload_0_14192);
  assign _zz_dataOut_payload_0_14242 = (_zz_dataOut_payload_0_14195 < _zz_dataOut_payload_0_14219);
  assign _zz_dataOut_payload_0_14243 = (_zz_dataOut_payload_0_14242 ? _zz_dataOut_payload_0_14195 : _zz_dataOut_payload_0_14219);
  assign _zz_dataOut_payload_0_14244 = (_zz_dataOut_payload_0_14242 ? _zz_dataOut_payload_0_14219 : _zz_dataOut_payload_0_14195);
  assign _zz_dataOut_payload_0_14245 = (_zz_dataOut_payload_0_14198 < _zz_dataOut_payload_0_14222);
  assign _zz_dataOut_payload_0_14246 = (_zz_dataOut_payload_0_14245 ? _zz_dataOut_payload_0_14198 : _zz_dataOut_payload_0_14222);
  assign _zz_dataOut_payload_0_14247 = (_zz_dataOut_payload_0_14245 ? _zz_dataOut_payload_0_14222 : _zz_dataOut_payload_0_14198);
  assign _zz_dataOut_payload_0_14248 = (_zz_dataOut_payload_0_14225 < _zz_dataOut_payload_0_14237);
  assign _zz_dataOut_payload_0_14249 = (_zz_dataOut_payload_0_14248 ? _zz_dataOut_payload_0_14225 : _zz_dataOut_payload_0_14237);
  assign _zz_dataOut_payload_0_14250 = (_zz_dataOut_payload_0_14248 ? _zz_dataOut_payload_0_14237 : _zz_dataOut_payload_0_14225);
  assign _zz_dataOut_payload_0_14251 = (_zz_dataOut_payload_0_14228 < _zz_dataOut_payload_0_14240);
  assign _zz_dataOut_payload_0_14252 = (_zz_dataOut_payload_0_14251 ? _zz_dataOut_payload_0_14228 : _zz_dataOut_payload_0_14240);
  assign _zz_dataOut_payload_0_14253 = (_zz_dataOut_payload_0_14251 ? _zz_dataOut_payload_0_14240 : _zz_dataOut_payload_0_14228);
  assign _zz_dataOut_payload_0_14254 = (_zz_dataOut_payload_0_14231 < _zz_dataOut_payload_0_14243);
  assign _zz_dataOut_payload_0_14255 = (_zz_dataOut_payload_0_14254 ? _zz_dataOut_payload_0_14231 : _zz_dataOut_payload_0_14243);
  assign _zz_dataOut_payload_0_14256 = (_zz_dataOut_payload_0_14254 ? _zz_dataOut_payload_0_14243 : _zz_dataOut_payload_0_14231);
  assign _zz_dataOut_payload_0_14257 = (_zz_dataOut_payload_0_14234 < _zz_dataOut_payload_0_14246);
  assign _zz_dataOut_payload_0_14258 = (_zz_dataOut_payload_0_14257 ? _zz_dataOut_payload_0_14234 : _zz_dataOut_payload_0_14246);
  assign _zz_dataOut_payload_0_14259 = (_zz_dataOut_payload_0_14257 ? _zz_dataOut_payload_0_14246 : _zz_dataOut_payload_0_14234);
  assign _zz_dataOut_payload_0_14260 = (_zz_dataOut_payload_0_14249 < _zz_dataOut_payload_0_14255);
  assign _zz_dataOut_payload_0_14261 = (_zz_dataOut_payload_0_14260 ? _zz_dataOut_payload_0_14249 : _zz_dataOut_payload_0_14255);
  assign _zz_dataOut_payload_0_14262 = (_zz_dataOut_payload_0_14260 ? _zz_dataOut_payload_0_14255 : _zz_dataOut_payload_0_14249);
  assign _zz_dataOut_payload_0_14263 = (_zz_dataOut_payload_0_14252 < _zz_dataOut_payload_0_14258);
  assign _zz_dataOut_payload_0_14264 = (_zz_dataOut_payload_0_14263 ? _zz_dataOut_payload_0_14252 : _zz_dataOut_payload_0_14258);
  assign _zz_dataOut_payload_0_14265 = (_zz_dataOut_payload_0_14263 ? _zz_dataOut_payload_0_14258 : _zz_dataOut_payload_0_14252);
  assign _zz_dataOut_payload_0_14266 = (_zz_dataOut_payload_0_14261 < _zz_dataOut_payload_0_14264);
  assign _zz_dataOut_payload_0_14267 = (_zz_dataOut_payload_0_14262 < _zz_dataOut_payload_0_14265);
  assign _zz_dataOut_payload_0_14272 = (_zz_dataOut_payload_0_14250 < _zz_dataOut_payload_0_14256);
  assign _zz_dataOut_payload_0_14273 = (_zz_dataOut_payload_0_14272 ? _zz_dataOut_payload_0_14250 : _zz_dataOut_payload_0_14256);
  assign _zz_dataOut_payload_0_14274 = (_zz_dataOut_payload_0_14272 ? _zz_dataOut_payload_0_14256 : _zz_dataOut_payload_0_14250);
  assign _zz_dataOut_payload_0_14275 = (_zz_dataOut_payload_0_14253 < _zz_dataOut_payload_0_14259);
  assign _zz_dataOut_payload_0_14276 = (_zz_dataOut_payload_0_14275 ? _zz_dataOut_payload_0_14253 : _zz_dataOut_payload_0_14259);
  assign _zz_dataOut_payload_0_14277 = (_zz_dataOut_payload_0_14275 ? _zz_dataOut_payload_0_14259 : _zz_dataOut_payload_0_14253);
  assign _zz_dataOut_payload_0_14278 = (_zz_dataOut_payload_0_14273 < _zz_dataOut_payload_0_14276);
  assign _zz_dataOut_payload_0_14279 = (_zz_dataOut_payload_0_14274 < _zz_dataOut_payload_0_14277);
  assign _zz_dataOut_payload_0_14292 = (_zz_dataOut_payload_0_14226 < _zz_dataOut_payload_0_14238);
  assign _zz_dataOut_payload_0_14293 = (_zz_dataOut_payload_0_14292 ? _zz_dataOut_payload_0_14226 : _zz_dataOut_payload_0_14238);
  assign _zz_dataOut_payload_0_14294 = (_zz_dataOut_payload_0_14292 ? _zz_dataOut_payload_0_14238 : _zz_dataOut_payload_0_14226);
  assign _zz_dataOut_payload_0_14295 = (_zz_dataOut_payload_0_14229 < _zz_dataOut_payload_0_14241);
  assign _zz_dataOut_payload_0_14296 = (_zz_dataOut_payload_0_14295 ? _zz_dataOut_payload_0_14229 : _zz_dataOut_payload_0_14241);
  assign _zz_dataOut_payload_0_14297 = (_zz_dataOut_payload_0_14295 ? _zz_dataOut_payload_0_14241 : _zz_dataOut_payload_0_14229);
  assign _zz_dataOut_payload_0_14298 = (_zz_dataOut_payload_0_14232 < _zz_dataOut_payload_0_14244);
  assign _zz_dataOut_payload_0_14299 = (_zz_dataOut_payload_0_14298 ? _zz_dataOut_payload_0_14232 : _zz_dataOut_payload_0_14244);
  assign _zz_dataOut_payload_0_14300 = (_zz_dataOut_payload_0_14298 ? _zz_dataOut_payload_0_14244 : _zz_dataOut_payload_0_14232);
  assign _zz_dataOut_payload_0_14301 = (_zz_dataOut_payload_0_14235 < _zz_dataOut_payload_0_14247);
  assign _zz_dataOut_payload_0_14302 = (_zz_dataOut_payload_0_14301 ? _zz_dataOut_payload_0_14235 : _zz_dataOut_payload_0_14247);
  assign _zz_dataOut_payload_0_14303 = (_zz_dataOut_payload_0_14301 ? _zz_dataOut_payload_0_14247 : _zz_dataOut_payload_0_14235);
  assign _zz_dataOut_payload_0_14304 = (_zz_dataOut_payload_0_14293 < _zz_dataOut_payload_0_14299);
  assign _zz_dataOut_payload_0_14305 = (_zz_dataOut_payload_0_14304 ? _zz_dataOut_payload_0_14293 : _zz_dataOut_payload_0_14299);
  assign _zz_dataOut_payload_0_14306 = (_zz_dataOut_payload_0_14304 ? _zz_dataOut_payload_0_14299 : _zz_dataOut_payload_0_14293);
  assign _zz_dataOut_payload_0_14307 = (_zz_dataOut_payload_0_14296 < _zz_dataOut_payload_0_14302);
  assign _zz_dataOut_payload_0_14308 = (_zz_dataOut_payload_0_14307 ? _zz_dataOut_payload_0_14296 : _zz_dataOut_payload_0_14302);
  assign _zz_dataOut_payload_0_14309 = (_zz_dataOut_payload_0_14307 ? _zz_dataOut_payload_0_14302 : _zz_dataOut_payload_0_14296);
  assign _zz_dataOut_payload_0_14310 = (_zz_dataOut_payload_0_14305 < _zz_dataOut_payload_0_14308);
  assign _zz_dataOut_payload_0_14311 = (_zz_dataOut_payload_0_14306 < _zz_dataOut_payload_0_14309);
  assign _zz_dataOut_payload_0_14316 = (_zz_dataOut_payload_0_14294 < _zz_dataOut_payload_0_14300);
  assign _zz_dataOut_payload_0_14317 = (_zz_dataOut_payload_0_14316 ? _zz_dataOut_payload_0_14294 : _zz_dataOut_payload_0_14300);
  assign _zz_dataOut_payload_0_14318 = (_zz_dataOut_payload_0_14316 ? _zz_dataOut_payload_0_14300 : _zz_dataOut_payload_0_14294);
  assign _zz_dataOut_payload_0_14319 = (_zz_dataOut_payload_0_14297 < _zz_dataOut_payload_0_14303);
  assign _zz_dataOut_payload_0_14320 = (_zz_dataOut_payload_0_14319 ? _zz_dataOut_payload_0_14297 : _zz_dataOut_payload_0_14303);
  assign _zz_dataOut_payload_0_14321 = (_zz_dataOut_payload_0_14319 ? _zz_dataOut_payload_0_14303 : _zz_dataOut_payload_0_14297);
  assign _zz_dataOut_payload_0_14322 = (_zz_dataOut_payload_0_14317 < _zz_dataOut_payload_0_14320);
  assign _zz_dataOut_payload_0_14323 = (_zz_dataOut_payload_0_14318 < _zz_dataOut_payload_0_14321);
  assign _zz_dataOut_payload_0_14352 = (_zz_dataOut_payload_0_14178 < _zz_dataOut_payload_0_14202);
  assign _zz_dataOut_payload_0_14353 = (_zz_dataOut_payload_0_14352 ? _zz_dataOut_payload_0_14178 : _zz_dataOut_payload_0_14202);
  assign _zz_dataOut_payload_0_14354 = (_zz_dataOut_payload_0_14352 ? _zz_dataOut_payload_0_14202 : _zz_dataOut_payload_0_14178);
  assign _zz_dataOut_payload_0_14355 = (_zz_dataOut_payload_0_14181 < _zz_dataOut_payload_0_14205);
  assign _zz_dataOut_payload_0_14356 = (_zz_dataOut_payload_0_14355 ? _zz_dataOut_payload_0_14181 : _zz_dataOut_payload_0_14205);
  assign _zz_dataOut_payload_0_14357 = (_zz_dataOut_payload_0_14355 ? _zz_dataOut_payload_0_14205 : _zz_dataOut_payload_0_14181);
  assign _zz_dataOut_payload_0_14358 = (_zz_dataOut_payload_0_14184 < _zz_dataOut_payload_0_14208);
  assign _zz_dataOut_payload_0_14359 = (_zz_dataOut_payload_0_14358 ? _zz_dataOut_payload_0_14184 : _zz_dataOut_payload_0_14208);
  assign _zz_dataOut_payload_0_14360 = (_zz_dataOut_payload_0_14358 ? _zz_dataOut_payload_0_14208 : _zz_dataOut_payload_0_14184);
  assign _zz_dataOut_payload_0_14361 = (_zz_dataOut_payload_0_14187 < _zz_dataOut_payload_0_14211);
  assign _zz_dataOut_payload_0_14362 = (_zz_dataOut_payload_0_14361 ? _zz_dataOut_payload_0_14187 : _zz_dataOut_payload_0_14211);
  assign _zz_dataOut_payload_0_14363 = (_zz_dataOut_payload_0_14361 ? _zz_dataOut_payload_0_14211 : _zz_dataOut_payload_0_14187);
  assign _zz_dataOut_payload_0_14364 = (_zz_dataOut_payload_0_14190 < _zz_dataOut_payload_0_14214);
  assign _zz_dataOut_payload_0_14365 = (_zz_dataOut_payload_0_14364 ? _zz_dataOut_payload_0_14190 : _zz_dataOut_payload_0_14214);
  assign _zz_dataOut_payload_0_14366 = (_zz_dataOut_payload_0_14364 ? _zz_dataOut_payload_0_14214 : _zz_dataOut_payload_0_14190);
  assign _zz_dataOut_payload_0_14367 = (_zz_dataOut_payload_0_14193 < _zz_dataOut_payload_0_14217);
  assign _zz_dataOut_payload_0_14368 = (_zz_dataOut_payload_0_14367 ? _zz_dataOut_payload_0_14193 : _zz_dataOut_payload_0_14217);
  assign _zz_dataOut_payload_0_14369 = (_zz_dataOut_payload_0_14367 ? _zz_dataOut_payload_0_14217 : _zz_dataOut_payload_0_14193);
  assign _zz_dataOut_payload_0_14370 = (_zz_dataOut_payload_0_14196 < _zz_dataOut_payload_0_14220);
  assign _zz_dataOut_payload_0_14371 = (_zz_dataOut_payload_0_14370 ? _zz_dataOut_payload_0_14196 : _zz_dataOut_payload_0_14220);
  assign _zz_dataOut_payload_0_14372 = (_zz_dataOut_payload_0_14370 ? _zz_dataOut_payload_0_14220 : _zz_dataOut_payload_0_14196);
  assign _zz_dataOut_payload_0_14373 = (_zz_dataOut_payload_0_14199 < _zz_dataOut_payload_0_14223);
  assign _zz_dataOut_payload_0_14374 = (_zz_dataOut_payload_0_14373 ? _zz_dataOut_payload_0_14199 : _zz_dataOut_payload_0_14223);
  assign _zz_dataOut_payload_0_14375 = (_zz_dataOut_payload_0_14373 ? _zz_dataOut_payload_0_14223 : _zz_dataOut_payload_0_14199);
  assign _zz_dataOut_payload_0_14376 = (_zz_dataOut_payload_0_14353 < _zz_dataOut_payload_0_14365);
  assign _zz_dataOut_payload_0_14377 = (_zz_dataOut_payload_0_14376 ? _zz_dataOut_payload_0_14353 : _zz_dataOut_payload_0_14365);
  assign _zz_dataOut_payload_0_14378 = (_zz_dataOut_payload_0_14376 ? _zz_dataOut_payload_0_14365 : _zz_dataOut_payload_0_14353);
  assign _zz_dataOut_payload_0_14379 = (_zz_dataOut_payload_0_14356 < _zz_dataOut_payload_0_14368);
  assign _zz_dataOut_payload_0_14380 = (_zz_dataOut_payload_0_14379 ? _zz_dataOut_payload_0_14356 : _zz_dataOut_payload_0_14368);
  assign _zz_dataOut_payload_0_14381 = (_zz_dataOut_payload_0_14379 ? _zz_dataOut_payload_0_14368 : _zz_dataOut_payload_0_14356);
  assign _zz_dataOut_payload_0_14382 = (_zz_dataOut_payload_0_14359 < _zz_dataOut_payload_0_14371);
  assign _zz_dataOut_payload_0_14383 = (_zz_dataOut_payload_0_14382 ? _zz_dataOut_payload_0_14359 : _zz_dataOut_payload_0_14371);
  assign _zz_dataOut_payload_0_14384 = (_zz_dataOut_payload_0_14382 ? _zz_dataOut_payload_0_14371 : _zz_dataOut_payload_0_14359);
  assign _zz_dataOut_payload_0_14385 = (_zz_dataOut_payload_0_14362 < _zz_dataOut_payload_0_14374);
  assign _zz_dataOut_payload_0_14386 = (_zz_dataOut_payload_0_14385 ? _zz_dataOut_payload_0_14362 : _zz_dataOut_payload_0_14374);
  assign _zz_dataOut_payload_0_14387 = (_zz_dataOut_payload_0_14385 ? _zz_dataOut_payload_0_14374 : _zz_dataOut_payload_0_14362);
  assign _zz_dataOut_payload_0_14388 = (_zz_dataOut_payload_0_14377 < _zz_dataOut_payload_0_14383);
  assign _zz_dataOut_payload_0_14389 = (_zz_dataOut_payload_0_14388 ? _zz_dataOut_payload_0_14377 : _zz_dataOut_payload_0_14383);
  assign _zz_dataOut_payload_0_14390 = (_zz_dataOut_payload_0_14388 ? _zz_dataOut_payload_0_14383 : _zz_dataOut_payload_0_14377);
  assign _zz_dataOut_payload_0_14391 = (_zz_dataOut_payload_0_14380 < _zz_dataOut_payload_0_14386);
  assign _zz_dataOut_payload_0_14392 = (_zz_dataOut_payload_0_14391 ? _zz_dataOut_payload_0_14380 : _zz_dataOut_payload_0_14386);
  assign _zz_dataOut_payload_0_14393 = (_zz_dataOut_payload_0_14391 ? _zz_dataOut_payload_0_14386 : _zz_dataOut_payload_0_14380);
  assign _zz_dataOut_payload_0_14394 = (_zz_dataOut_payload_0_14389 < _zz_dataOut_payload_0_14392);
  assign _zz_dataOut_payload_0_14395 = (_zz_dataOut_payload_0_14390 < _zz_dataOut_payload_0_14393);
  assign _zz_dataOut_payload_0_14400 = (_zz_dataOut_payload_0_14378 < _zz_dataOut_payload_0_14384);
  assign _zz_dataOut_payload_0_14401 = (_zz_dataOut_payload_0_14400 ? _zz_dataOut_payload_0_14378 : _zz_dataOut_payload_0_14384);
  assign _zz_dataOut_payload_0_14402 = (_zz_dataOut_payload_0_14400 ? _zz_dataOut_payload_0_14384 : _zz_dataOut_payload_0_14378);
  assign _zz_dataOut_payload_0_14403 = (_zz_dataOut_payload_0_14381 < _zz_dataOut_payload_0_14387);
  assign _zz_dataOut_payload_0_14404 = (_zz_dataOut_payload_0_14403 ? _zz_dataOut_payload_0_14381 : _zz_dataOut_payload_0_14387);
  assign _zz_dataOut_payload_0_14405 = (_zz_dataOut_payload_0_14403 ? _zz_dataOut_payload_0_14387 : _zz_dataOut_payload_0_14381);
  assign _zz_dataOut_payload_0_14406 = (_zz_dataOut_payload_0_14401 < _zz_dataOut_payload_0_14404);
  assign _zz_dataOut_payload_0_14407 = (_zz_dataOut_payload_0_14402 < _zz_dataOut_payload_0_14405);
  assign _zz_dataOut_payload_0_14420 = (_zz_dataOut_payload_0_14354 < _zz_dataOut_payload_0_14366);
  assign _zz_dataOut_payload_0_14421 = (_zz_dataOut_payload_0_14420 ? _zz_dataOut_payload_0_14354 : _zz_dataOut_payload_0_14366);
  assign _zz_dataOut_payload_0_14422 = (_zz_dataOut_payload_0_14420 ? _zz_dataOut_payload_0_14366 : _zz_dataOut_payload_0_14354);
  assign _zz_dataOut_payload_0_14423 = (_zz_dataOut_payload_0_14357 < _zz_dataOut_payload_0_14369);
  assign _zz_dataOut_payload_0_14424 = (_zz_dataOut_payload_0_14423 ? _zz_dataOut_payload_0_14357 : _zz_dataOut_payload_0_14369);
  assign _zz_dataOut_payload_0_14425 = (_zz_dataOut_payload_0_14423 ? _zz_dataOut_payload_0_14369 : _zz_dataOut_payload_0_14357);
  assign _zz_dataOut_payload_0_14426 = (_zz_dataOut_payload_0_14360 < _zz_dataOut_payload_0_14372);
  assign _zz_dataOut_payload_0_14427 = (_zz_dataOut_payload_0_14426 ? _zz_dataOut_payload_0_14360 : _zz_dataOut_payload_0_14372);
  assign _zz_dataOut_payload_0_14428 = (_zz_dataOut_payload_0_14426 ? _zz_dataOut_payload_0_14372 : _zz_dataOut_payload_0_14360);
  assign _zz_dataOut_payload_0_14429 = (_zz_dataOut_payload_0_14363 < _zz_dataOut_payload_0_14375);
  assign _zz_dataOut_payload_0_14430 = (_zz_dataOut_payload_0_14429 ? _zz_dataOut_payload_0_14363 : _zz_dataOut_payload_0_14375);
  assign _zz_dataOut_payload_0_14431 = (_zz_dataOut_payload_0_14429 ? _zz_dataOut_payload_0_14375 : _zz_dataOut_payload_0_14363);
  assign _zz_dataOut_payload_0_14432 = (_zz_dataOut_payload_0_14421 < _zz_dataOut_payload_0_14427);
  assign _zz_dataOut_payload_0_14433 = (_zz_dataOut_payload_0_14432 ? _zz_dataOut_payload_0_14421 : _zz_dataOut_payload_0_14427);
  assign _zz_dataOut_payload_0_14434 = (_zz_dataOut_payload_0_14432 ? _zz_dataOut_payload_0_14427 : _zz_dataOut_payload_0_14421);
  assign _zz_dataOut_payload_0_14435 = (_zz_dataOut_payload_0_14424 < _zz_dataOut_payload_0_14430);
  assign _zz_dataOut_payload_0_14436 = (_zz_dataOut_payload_0_14435 ? _zz_dataOut_payload_0_14424 : _zz_dataOut_payload_0_14430);
  assign _zz_dataOut_payload_0_14437 = (_zz_dataOut_payload_0_14435 ? _zz_dataOut_payload_0_14430 : _zz_dataOut_payload_0_14424);
  assign _zz_dataOut_payload_0_14438 = (_zz_dataOut_payload_0_14433 < _zz_dataOut_payload_0_14436);
  assign _zz_dataOut_payload_0_14439 = (_zz_dataOut_payload_0_14434 < _zz_dataOut_payload_0_14437);
  assign _zz_dataOut_payload_0_14444 = (_zz_dataOut_payload_0_14422 < _zz_dataOut_payload_0_14428);
  assign _zz_dataOut_payload_0_14445 = (_zz_dataOut_payload_0_14444 ? _zz_dataOut_payload_0_14422 : _zz_dataOut_payload_0_14428);
  assign _zz_dataOut_payload_0_14446 = (_zz_dataOut_payload_0_14444 ? _zz_dataOut_payload_0_14428 : _zz_dataOut_payload_0_14422);
  assign _zz_dataOut_payload_0_14447 = (_zz_dataOut_payload_0_14425 < _zz_dataOut_payload_0_14431);
  assign _zz_dataOut_payload_0_14448 = (_zz_dataOut_payload_0_14447 ? _zz_dataOut_payload_0_14425 : _zz_dataOut_payload_0_14431);
  assign _zz_dataOut_payload_0_14449 = (_zz_dataOut_payload_0_14447 ? _zz_dataOut_payload_0_14431 : _zz_dataOut_payload_0_14425);
  assign _zz_dataOut_payload_0_14450 = (_zz_dataOut_payload_0_14445 < _zz_dataOut_payload_0_14448);
  assign _zz_dataOut_payload_0_14451 = (_zz_dataOut_payload_0_14446 < _zz_dataOut_payload_0_14449);
  assign _zz_dataOut_payload_0_14512 = (_zz_dataOut_payload_0_14082 < _zz_dataOut_payload_0_14130);
  assign _zz_dataOut_payload_0_14513 = (_zz_dataOut_payload_0_14512 ? _zz_dataOut_payload_0_14082 : _zz_dataOut_payload_0_14130);
  assign _zz_dataOut_payload_0_14514 = (_zz_dataOut_payload_0_14512 ? _zz_dataOut_payload_0_14130 : _zz_dataOut_payload_0_14082);
  assign _zz_dataOut_payload_0_14515 = (_zz_dataOut_payload_0_14085 < _zz_dataOut_payload_0_14133);
  assign _zz_dataOut_payload_0_14516 = (_zz_dataOut_payload_0_14515 ? _zz_dataOut_payload_0_14085 : _zz_dataOut_payload_0_14133);
  assign _zz_dataOut_payload_0_14517 = (_zz_dataOut_payload_0_14515 ? _zz_dataOut_payload_0_14133 : _zz_dataOut_payload_0_14085);
  assign _zz_dataOut_payload_0_14518 = (_zz_dataOut_payload_0_14088 < _zz_dataOut_payload_0_14136);
  assign _zz_dataOut_payload_0_14519 = (_zz_dataOut_payload_0_14518 ? _zz_dataOut_payload_0_14088 : _zz_dataOut_payload_0_14136);
  assign _zz_dataOut_payload_0_14520 = (_zz_dataOut_payload_0_14518 ? _zz_dataOut_payload_0_14136 : _zz_dataOut_payload_0_14088);
  assign _zz_dataOut_payload_0_14521 = (_zz_dataOut_payload_0_14091 < _zz_dataOut_payload_0_14139);
  assign _zz_dataOut_payload_0_14522 = (_zz_dataOut_payload_0_14521 ? _zz_dataOut_payload_0_14091 : _zz_dataOut_payload_0_14139);
  assign _zz_dataOut_payload_0_14523 = (_zz_dataOut_payload_0_14521 ? _zz_dataOut_payload_0_14139 : _zz_dataOut_payload_0_14091);
  assign _zz_dataOut_payload_0_14524 = (_zz_dataOut_payload_0_14094 < _zz_dataOut_payload_0_14142);
  assign _zz_dataOut_payload_0_14525 = (_zz_dataOut_payload_0_14524 ? _zz_dataOut_payload_0_14094 : _zz_dataOut_payload_0_14142);
  assign _zz_dataOut_payload_0_14526 = (_zz_dataOut_payload_0_14524 ? _zz_dataOut_payload_0_14142 : _zz_dataOut_payload_0_14094);
  assign _zz_dataOut_payload_0_14527 = (_zz_dataOut_payload_0_14097 < _zz_dataOut_payload_0_14145);
  assign _zz_dataOut_payload_0_14528 = (_zz_dataOut_payload_0_14527 ? _zz_dataOut_payload_0_14097 : _zz_dataOut_payload_0_14145);
  assign _zz_dataOut_payload_0_14529 = (_zz_dataOut_payload_0_14527 ? _zz_dataOut_payload_0_14145 : _zz_dataOut_payload_0_14097);
  assign _zz_dataOut_payload_0_14530 = (_zz_dataOut_payload_0_14100 < _zz_dataOut_payload_0_14148);
  assign _zz_dataOut_payload_0_14531 = (_zz_dataOut_payload_0_14530 ? _zz_dataOut_payload_0_14100 : _zz_dataOut_payload_0_14148);
  assign _zz_dataOut_payload_0_14532 = (_zz_dataOut_payload_0_14530 ? _zz_dataOut_payload_0_14148 : _zz_dataOut_payload_0_14100);
  assign _zz_dataOut_payload_0_14533 = (_zz_dataOut_payload_0_14103 < _zz_dataOut_payload_0_14151);
  assign _zz_dataOut_payload_0_14534 = (_zz_dataOut_payload_0_14533 ? _zz_dataOut_payload_0_14103 : _zz_dataOut_payload_0_14151);
  assign _zz_dataOut_payload_0_14535 = (_zz_dataOut_payload_0_14533 ? _zz_dataOut_payload_0_14151 : _zz_dataOut_payload_0_14103);
  assign _zz_dataOut_payload_0_14536 = (_zz_dataOut_payload_0_14106 < _zz_dataOut_payload_0_14154);
  assign _zz_dataOut_payload_0_14537 = (_zz_dataOut_payload_0_14536 ? _zz_dataOut_payload_0_14106 : _zz_dataOut_payload_0_14154);
  assign _zz_dataOut_payload_0_14538 = (_zz_dataOut_payload_0_14536 ? _zz_dataOut_payload_0_14154 : _zz_dataOut_payload_0_14106);
  assign _zz_dataOut_payload_0_14539 = (_zz_dataOut_payload_0_14109 < _zz_dataOut_payload_0_14157);
  assign _zz_dataOut_payload_0_14540 = (_zz_dataOut_payload_0_14539 ? _zz_dataOut_payload_0_14109 : _zz_dataOut_payload_0_14157);
  assign _zz_dataOut_payload_0_14541 = (_zz_dataOut_payload_0_14539 ? _zz_dataOut_payload_0_14157 : _zz_dataOut_payload_0_14109);
  assign _zz_dataOut_payload_0_14542 = (_zz_dataOut_payload_0_14112 < _zz_dataOut_payload_0_14160);
  assign _zz_dataOut_payload_0_14543 = (_zz_dataOut_payload_0_14542 ? _zz_dataOut_payload_0_14112 : _zz_dataOut_payload_0_14160);
  assign _zz_dataOut_payload_0_14544 = (_zz_dataOut_payload_0_14542 ? _zz_dataOut_payload_0_14160 : _zz_dataOut_payload_0_14112);
  assign _zz_dataOut_payload_0_14545 = (_zz_dataOut_payload_0_14115 < _zz_dataOut_payload_0_14163);
  assign _zz_dataOut_payload_0_14546 = (_zz_dataOut_payload_0_14545 ? _zz_dataOut_payload_0_14115 : _zz_dataOut_payload_0_14163);
  assign _zz_dataOut_payload_0_14547 = (_zz_dataOut_payload_0_14545 ? _zz_dataOut_payload_0_14163 : _zz_dataOut_payload_0_14115);
  assign _zz_dataOut_payload_0_14548 = (_zz_dataOut_payload_0_14118 < _zz_dataOut_payload_0_14166);
  assign _zz_dataOut_payload_0_14549 = (_zz_dataOut_payload_0_14548 ? _zz_dataOut_payload_0_14118 : _zz_dataOut_payload_0_14166);
  assign _zz_dataOut_payload_0_14550 = (_zz_dataOut_payload_0_14548 ? _zz_dataOut_payload_0_14166 : _zz_dataOut_payload_0_14118);
  assign _zz_dataOut_payload_0_14551 = (_zz_dataOut_payload_0_14121 < _zz_dataOut_payload_0_14169);
  assign _zz_dataOut_payload_0_14552 = (_zz_dataOut_payload_0_14551 ? _zz_dataOut_payload_0_14121 : _zz_dataOut_payload_0_14169);
  assign _zz_dataOut_payload_0_14553 = (_zz_dataOut_payload_0_14551 ? _zz_dataOut_payload_0_14169 : _zz_dataOut_payload_0_14121);
  assign _zz_dataOut_payload_0_14554 = (_zz_dataOut_payload_0_14124 < _zz_dataOut_payload_0_14172);
  assign _zz_dataOut_payload_0_14555 = (_zz_dataOut_payload_0_14554 ? _zz_dataOut_payload_0_14124 : _zz_dataOut_payload_0_14172);
  assign _zz_dataOut_payload_0_14556 = (_zz_dataOut_payload_0_14554 ? _zz_dataOut_payload_0_14172 : _zz_dataOut_payload_0_14124);
  assign _zz_dataOut_payload_0_14557 = (_zz_dataOut_payload_0_14127 < _zz_dataOut_payload_0_14175);
  assign _zz_dataOut_payload_0_14558 = (_zz_dataOut_payload_0_14557 ? _zz_dataOut_payload_0_14127 : _zz_dataOut_payload_0_14175);
  assign _zz_dataOut_payload_0_14559 = (_zz_dataOut_payload_0_14557 ? _zz_dataOut_payload_0_14175 : _zz_dataOut_payload_0_14127);
  assign _zz_dataOut_payload_0_14560 = (_zz_dataOut_payload_0_14513 < _zz_dataOut_payload_0_14537);
  assign _zz_dataOut_payload_0_14561 = (_zz_dataOut_payload_0_14560 ? _zz_dataOut_payload_0_14513 : _zz_dataOut_payload_0_14537);
  assign _zz_dataOut_payload_0_14562 = (_zz_dataOut_payload_0_14560 ? _zz_dataOut_payload_0_14537 : _zz_dataOut_payload_0_14513);
  assign _zz_dataOut_payload_0_14563 = (_zz_dataOut_payload_0_14516 < _zz_dataOut_payload_0_14540);
  assign _zz_dataOut_payload_0_14564 = (_zz_dataOut_payload_0_14563 ? _zz_dataOut_payload_0_14516 : _zz_dataOut_payload_0_14540);
  assign _zz_dataOut_payload_0_14565 = (_zz_dataOut_payload_0_14563 ? _zz_dataOut_payload_0_14540 : _zz_dataOut_payload_0_14516);
  assign _zz_dataOut_payload_0_14566 = (_zz_dataOut_payload_0_14519 < _zz_dataOut_payload_0_14543);
  assign _zz_dataOut_payload_0_14567 = (_zz_dataOut_payload_0_14566 ? _zz_dataOut_payload_0_14519 : _zz_dataOut_payload_0_14543);
  assign _zz_dataOut_payload_0_14568 = (_zz_dataOut_payload_0_14566 ? _zz_dataOut_payload_0_14543 : _zz_dataOut_payload_0_14519);
  assign _zz_dataOut_payload_0_14569 = (_zz_dataOut_payload_0_14522 < _zz_dataOut_payload_0_14546);
  assign _zz_dataOut_payload_0_14570 = (_zz_dataOut_payload_0_14569 ? _zz_dataOut_payload_0_14522 : _zz_dataOut_payload_0_14546);
  assign _zz_dataOut_payload_0_14571 = (_zz_dataOut_payload_0_14569 ? _zz_dataOut_payload_0_14546 : _zz_dataOut_payload_0_14522);
  assign _zz_dataOut_payload_0_14572 = (_zz_dataOut_payload_0_14525 < _zz_dataOut_payload_0_14549);
  assign _zz_dataOut_payload_0_14573 = (_zz_dataOut_payload_0_14572 ? _zz_dataOut_payload_0_14525 : _zz_dataOut_payload_0_14549);
  assign _zz_dataOut_payload_0_14574 = (_zz_dataOut_payload_0_14572 ? _zz_dataOut_payload_0_14549 : _zz_dataOut_payload_0_14525);
  assign _zz_dataOut_payload_0_14575 = (_zz_dataOut_payload_0_14528 < _zz_dataOut_payload_0_14552);
  assign _zz_dataOut_payload_0_14576 = (_zz_dataOut_payload_0_14575 ? _zz_dataOut_payload_0_14528 : _zz_dataOut_payload_0_14552);
  assign _zz_dataOut_payload_0_14577 = (_zz_dataOut_payload_0_14575 ? _zz_dataOut_payload_0_14552 : _zz_dataOut_payload_0_14528);
  assign _zz_dataOut_payload_0_14578 = (_zz_dataOut_payload_0_14531 < _zz_dataOut_payload_0_14555);
  assign _zz_dataOut_payload_0_14579 = (_zz_dataOut_payload_0_14578 ? _zz_dataOut_payload_0_14531 : _zz_dataOut_payload_0_14555);
  assign _zz_dataOut_payload_0_14580 = (_zz_dataOut_payload_0_14578 ? _zz_dataOut_payload_0_14555 : _zz_dataOut_payload_0_14531);
  assign _zz_dataOut_payload_0_14581 = (_zz_dataOut_payload_0_14534 < _zz_dataOut_payload_0_14558);
  assign _zz_dataOut_payload_0_14582 = (_zz_dataOut_payload_0_14581 ? _zz_dataOut_payload_0_14534 : _zz_dataOut_payload_0_14558);
  assign _zz_dataOut_payload_0_14583 = (_zz_dataOut_payload_0_14581 ? _zz_dataOut_payload_0_14558 : _zz_dataOut_payload_0_14534);
  assign _zz_dataOut_payload_0_14584 = (_zz_dataOut_payload_0_14561 < _zz_dataOut_payload_0_14573);
  assign _zz_dataOut_payload_0_14585 = (_zz_dataOut_payload_0_14584 ? _zz_dataOut_payload_0_14561 : _zz_dataOut_payload_0_14573);
  assign _zz_dataOut_payload_0_14586 = (_zz_dataOut_payload_0_14584 ? _zz_dataOut_payload_0_14573 : _zz_dataOut_payload_0_14561);
  assign _zz_dataOut_payload_0_14587 = (_zz_dataOut_payload_0_14564 < _zz_dataOut_payload_0_14576);
  assign _zz_dataOut_payload_0_14588 = (_zz_dataOut_payload_0_14587 ? _zz_dataOut_payload_0_14564 : _zz_dataOut_payload_0_14576);
  assign _zz_dataOut_payload_0_14589 = (_zz_dataOut_payload_0_14587 ? _zz_dataOut_payload_0_14576 : _zz_dataOut_payload_0_14564);
  assign _zz_dataOut_payload_0_14590 = (_zz_dataOut_payload_0_14567 < _zz_dataOut_payload_0_14579);
  assign _zz_dataOut_payload_0_14591 = (_zz_dataOut_payload_0_14590 ? _zz_dataOut_payload_0_14567 : _zz_dataOut_payload_0_14579);
  assign _zz_dataOut_payload_0_14592 = (_zz_dataOut_payload_0_14590 ? _zz_dataOut_payload_0_14579 : _zz_dataOut_payload_0_14567);
  assign _zz_dataOut_payload_0_14593 = (_zz_dataOut_payload_0_14570 < _zz_dataOut_payload_0_14582);
  assign _zz_dataOut_payload_0_14594 = (_zz_dataOut_payload_0_14593 ? _zz_dataOut_payload_0_14570 : _zz_dataOut_payload_0_14582);
  assign _zz_dataOut_payload_0_14595 = (_zz_dataOut_payload_0_14593 ? _zz_dataOut_payload_0_14582 : _zz_dataOut_payload_0_14570);
  assign _zz_dataOut_payload_0_14596 = (_zz_dataOut_payload_0_14585 < _zz_dataOut_payload_0_14591);
  assign _zz_dataOut_payload_0_14597 = (_zz_dataOut_payload_0_14596 ? _zz_dataOut_payload_0_14585 : _zz_dataOut_payload_0_14591);
  assign _zz_dataOut_payload_0_14598 = (_zz_dataOut_payload_0_14596 ? _zz_dataOut_payload_0_14591 : _zz_dataOut_payload_0_14585);
  assign _zz_dataOut_payload_0_14599 = (_zz_dataOut_payload_0_14588 < _zz_dataOut_payload_0_14594);
  assign _zz_dataOut_payload_0_14600 = (_zz_dataOut_payload_0_14599 ? _zz_dataOut_payload_0_14588 : _zz_dataOut_payload_0_14594);
  assign _zz_dataOut_payload_0_14601 = (_zz_dataOut_payload_0_14599 ? _zz_dataOut_payload_0_14594 : _zz_dataOut_payload_0_14588);
  assign _zz_dataOut_payload_0_14602 = (_zz_dataOut_payload_0_14597 < _zz_dataOut_payload_0_14600);
  assign _zz_dataOut_payload_0_14603 = (_zz_dataOut_payload_0_14598 < _zz_dataOut_payload_0_14601);
  assign _zz_dataOut_payload_0_14608 = (_zz_dataOut_payload_0_14586 < _zz_dataOut_payload_0_14592);
  assign _zz_dataOut_payload_0_14609 = (_zz_dataOut_payload_0_14608 ? _zz_dataOut_payload_0_14586 : _zz_dataOut_payload_0_14592);
  assign _zz_dataOut_payload_0_14610 = (_zz_dataOut_payload_0_14608 ? _zz_dataOut_payload_0_14592 : _zz_dataOut_payload_0_14586);
  assign _zz_dataOut_payload_0_14611 = (_zz_dataOut_payload_0_14589 < _zz_dataOut_payload_0_14595);
  assign _zz_dataOut_payload_0_14612 = (_zz_dataOut_payload_0_14611 ? _zz_dataOut_payload_0_14589 : _zz_dataOut_payload_0_14595);
  assign _zz_dataOut_payload_0_14613 = (_zz_dataOut_payload_0_14611 ? _zz_dataOut_payload_0_14595 : _zz_dataOut_payload_0_14589);
  assign _zz_dataOut_payload_0_14614 = (_zz_dataOut_payload_0_14609 < _zz_dataOut_payload_0_14612);
  assign _zz_dataOut_payload_0_14615 = (_zz_dataOut_payload_0_14610 < _zz_dataOut_payload_0_14613);
  assign _zz_dataOut_payload_0_14628 = (_zz_dataOut_payload_0_14562 < _zz_dataOut_payload_0_14574);
  assign _zz_dataOut_payload_0_14629 = (_zz_dataOut_payload_0_14628 ? _zz_dataOut_payload_0_14562 : _zz_dataOut_payload_0_14574);
  assign _zz_dataOut_payload_0_14630 = (_zz_dataOut_payload_0_14628 ? _zz_dataOut_payload_0_14574 : _zz_dataOut_payload_0_14562);
  assign _zz_dataOut_payload_0_14631 = (_zz_dataOut_payload_0_14565 < _zz_dataOut_payload_0_14577);
  assign _zz_dataOut_payload_0_14632 = (_zz_dataOut_payload_0_14631 ? _zz_dataOut_payload_0_14565 : _zz_dataOut_payload_0_14577);
  assign _zz_dataOut_payload_0_14633 = (_zz_dataOut_payload_0_14631 ? _zz_dataOut_payload_0_14577 : _zz_dataOut_payload_0_14565);
  assign _zz_dataOut_payload_0_14634 = (_zz_dataOut_payload_0_14568 < _zz_dataOut_payload_0_14580);
  assign _zz_dataOut_payload_0_14635 = (_zz_dataOut_payload_0_14634 ? _zz_dataOut_payload_0_14568 : _zz_dataOut_payload_0_14580);
  assign _zz_dataOut_payload_0_14636 = (_zz_dataOut_payload_0_14634 ? _zz_dataOut_payload_0_14580 : _zz_dataOut_payload_0_14568);
  assign _zz_dataOut_payload_0_14637 = (_zz_dataOut_payload_0_14571 < _zz_dataOut_payload_0_14583);
  assign _zz_dataOut_payload_0_14638 = (_zz_dataOut_payload_0_14637 ? _zz_dataOut_payload_0_14571 : _zz_dataOut_payload_0_14583);
  assign _zz_dataOut_payload_0_14639 = (_zz_dataOut_payload_0_14637 ? _zz_dataOut_payload_0_14583 : _zz_dataOut_payload_0_14571);
  assign _zz_dataOut_payload_0_14640 = (_zz_dataOut_payload_0_14629 < _zz_dataOut_payload_0_14635);
  assign _zz_dataOut_payload_0_14641 = (_zz_dataOut_payload_0_14640 ? _zz_dataOut_payload_0_14629 : _zz_dataOut_payload_0_14635);
  assign _zz_dataOut_payload_0_14642 = (_zz_dataOut_payload_0_14640 ? _zz_dataOut_payload_0_14635 : _zz_dataOut_payload_0_14629);
  assign _zz_dataOut_payload_0_14643 = (_zz_dataOut_payload_0_14632 < _zz_dataOut_payload_0_14638);
  assign _zz_dataOut_payload_0_14644 = (_zz_dataOut_payload_0_14643 ? _zz_dataOut_payload_0_14632 : _zz_dataOut_payload_0_14638);
  assign _zz_dataOut_payload_0_14645 = (_zz_dataOut_payload_0_14643 ? _zz_dataOut_payload_0_14638 : _zz_dataOut_payload_0_14632);
  assign _zz_dataOut_payload_0_14646 = (_zz_dataOut_payload_0_14641 < _zz_dataOut_payload_0_14644);
  assign _zz_dataOut_payload_0_14647 = (_zz_dataOut_payload_0_14642 < _zz_dataOut_payload_0_14645);
  assign _zz_dataOut_payload_0_14652 = (_zz_dataOut_payload_0_14630 < _zz_dataOut_payload_0_14636);
  assign _zz_dataOut_payload_0_14653 = (_zz_dataOut_payload_0_14652 ? _zz_dataOut_payload_0_14630 : _zz_dataOut_payload_0_14636);
  assign _zz_dataOut_payload_0_14654 = (_zz_dataOut_payload_0_14652 ? _zz_dataOut_payload_0_14636 : _zz_dataOut_payload_0_14630);
  assign _zz_dataOut_payload_0_14655 = (_zz_dataOut_payload_0_14633 < _zz_dataOut_payload_0_14639);
  assign _zz_dataOut_payload_0_14656 = (_zz_dataOut_payload_0_14655 ? _zz_dataOut_payload_0_14633 : _zz_dataOut_payload_0_14639);
  assign _zz_dataOut_payload_0_14657 = (_zz_dataOut_payload_0_14655 ? _zz_dataOut_payload_0_14639 : _zz_dataOut_payload_0_14633);
  assign _zz_dataOut_payload_0_14658 = (_zz_dataOut_payload_0_14653 < _zz_dataOut_payload_0_14656);
  assign _zz_dataOut_payload_0_14659 = (_zz_dataOut_payload_0_14654 < _zz_dataOut_payload_0_14657);
  assign _zz_dataOut_payload_0_14688 = (_zz_dataOut_payload_0_14514 < _zz_dataOut_payload_0_14538);
  assign _zz_dataOut_payload_0_14689 = (_zz_dataOut_payload_0_14688 ? _zz_dataOut_payload_0_14514 : _zz_dataOut_payload_0_14538);
  assign _zz_dataOut_payload_0_14690 = (_zz_dataOut_payload_0_14688 ? _zz_dataOut_payload_0_14538 : _zz_dataOut_payload_0_14514);
  assign _zz_dataOut_payload_0_14691 = (_zz_dataOut_payload_0_14517 < _zz_dataOut_payload_0_14541);
  assign _zz_dataOut_payload_0_14692 = (_zz_dataOut_payload_0_14691 ? _zz_dataOut_payload_0_14517 : _zz_dataOut_payload_0_14541);
  assign _zz_dataOut_payload_0_14693 = (_zz_dataOut_payload_0_14691 ? _zz_dataOut_payload_0_14541 : _zz_dataOut_payload_0_14517);
  assign _zz_dataOut_payload_0_14694 = (_zz_dataOut_payload_0_14520 < _zz_dataOut_payload_0_14544);
  assign _zz_dataOut_payload_0_14695 = (_zz_dataOut_payload_0_14694 ? _zz_dataOut_payload_0_14520 : _zz_dataOut_payload_0_14544);
  assign _zz_dataOut_payload_0_14696 = (_zz_dataOut_payload_0_14694 ? _zz_dataOut_payload_0_14544 : _zz_dataOut_payload_0_14520);
  assign _zz_dataOut_payload_0_14697 = (_zz_dataOut_payload_0_14523 < _zz_dataOut_payload_0_14547);
  assign _zz_dataOut_payload_0_14698 = (_zz_dataOut_payload_0_14697 ? _zz_dataOut_payload_0_14523 : _zz_dataOut_payload_0_14547);
  assign _zz_dataOut_payload_0_14699 = (_zz_dataOut_payload_0_14697 ? _zz_dataOut_payload_0_14547 : _zz_dataOut_payload_0_14523);
  assign _zz_dataOut_payload_0_14700 = (_zz_dataOut_payload_0_14526 < _zz_dataOut_payload_0_14550);
  assign _zz_dataOut_payload_0_14701 = (_zz_dataOut_payload_0_14700 ? _zz_dataOut_payload_0_14526 : _zz_dataOut_payload_0_14550);
  assign _zz_dataOut_payload_0_14702 = (_zz_dataOut_payload_0_14700 ? _zz_dataOut_payload_0_14550 : _zz_dataOut_payload_0_14526);
  assign _zz_dataOut_payload_0_14703 = (_zz_dataOut_payload_0_14529 < _zz_dataOut_payload_0_14553);
  assign _zz_dataOut_payload_0_14704 = (_zz_dataOut_payload_0_14703 ? _zz_dataOut_payload_0_14529 : _zz_dataOut_payload_0_14553);
  assign _zz_dataOut_payload_0_14705 = (_zz_dataOut_payload_0_14703 ? _zz_dataOut_payload_0_14553 : _zz_dataOut_payload_0_14529);
  assign _zz_dataOut_payload_0_14706 = (_zz_dataOut_payload_0_14532 < _zz_dataOut_payload_0_14556);
  assign _zz_dataOut_payload_0_14707 = (_zz_dataOut_payload_0_14706 ? _zz_dataOut_payload_0_14532 : _zz_dataOut_payload_0_14556);
  assign _zz_dataOut_payload_0_14708 = (_zz_dataOut_payload_0_14706 ? _zz_dataOut_payload_0_14556 : _zz_dataOut_payload_0_14532);
  assign _zz_dataOut_payload_0_14709 = (_zz_dataOut_payload_0_14535 < _zz_dataOut_payload_0_14559);
  assign _zz_dataOut_payload_0_14710 = (_zz_dataOut_payload_0_14709 ? _zz_dataOut_payload_0_14535 : _zz_dataOut_payload_0_14559);
  assign _zz_dataOut_payload_0_14711 = (_zz_dataOut_payload_0_14709 ? _zz_dataOut_payload_0_14559 : _zz_dataOut_payload_0_14535);
  assign _zz_dataOut_payload_0_14712 = (_zz_dataOut_payload_0_14689 < _zz_dataOut_payload_0_14701);
  assign _zz_dataOut_payload_0_14713 = (_zz_dataOut_payload_0_14712 ? _zz_dataOut_payload_0_14689 : _zz_dataOut_payload_0_14701);
  assign _zz_dataOut_payload_0_14714 = (_zz_dataOut_payload_0_14712 ? _zz_dataOut_payload_0_14701 : _zz_dataOut_payload_0_14689);
  assign _zz_dataOut_payload_0_14715 = (_zz_dataOut_payload_0_14692 < _zz_dataOut_payload_0_14704);
  assign _zz_dataOut_payload_0_14716 = (_zz_dataOut_payload_0_14715 ? _zz_dataOut_payload_0_14692 : _zz_dataOut_payload_0_14704);
  assign _zz_dataOut_payload_0_14717 = (_zz_dataOut_payload_0_14715 ? _zz_dataOut_payload_0_14704 : _zz_dataOut_payload_0_14692);
  assign _zz_dataOut_payload_0_14718 = (_zz_dataOut_payload_0_14695 < _zz_dataOut_payload_0_14707);
  assign _zz_dataOut_payload_0_14719 = (_zz_dataOut_payload_0_14718 ? _zz_dataOut_payload_0_14695 : _zz_dataOut_payload_0_14707);
  assign _zz_dataOut_payload_0_14720 = (_zz_dataOut_payload_0_14718 ? _zz_dataOut_payload_0_14707 : _zz_dataOut_payload_0_14695);
  assign _zz_dataOut_payload_0_14721 = (_zz_dataOut_payload_0_14698 < _zz_dataOut_payload_0_14710);
  assign _zz_dataOut_payload_0_14722 = (_zz_dataOut_payload_0_14721 ? _zz_dataOut_payload_0_14698 : _zz_dataOut_payload_0_14710);
  assign _zz_dataOut_payload_0_14723 = (_zz_dataOut_payload_0_14721 ? _zz_dataOut_payload_0_14710 : _zz_dataOut_payload_0_14698);
  assign _zz_dataOut_payload_0_14724 = (_zz_dataOut_payload_0_14713 < _zz_dataOut_payload_0_14719);
  assign _zz_dataOut_payload_0_14725 = (_zz_dataOut_payload_0_14724 ? _zz_dataOut_payload_0_14713 : _zz_dataOut_payload_0_14719);
  assign _zz_dataOut_payload_0_14726 = (_zz_dataOut_payload_0_14724 ? _zz_dataOut_payload_0_14719 : _zz_dataOut_payload_0_14713);
  assign _zz_dataOut_payload_0_14727 = (_zz_dataOut_payload_0_14716 < _zz_dataOut_payload_0_14722);
  assign _zz_dataOut_payload_0_14728 = (_zz_dataOut_payload_0_14727 ? _zz_dataOut_payload_0_14716 : _zz_dataOut_payload_0_14722);
  assign _zz_dataOut_payload_0_14729 = (_zz_dataOut_payload_0_14727 ? _zz_dataOut_payload_0_14722 : _zz_dataOut_payload_0_14716);
  assign _zz_dataOut_payload_0_14730 = (_zz_dataOut_payload_0_14725 < _zz_dataOut_payload_0_14728);
  assign _zz_dataOut_payload_0_14731 = (_zz_dataOut_payload_0_14726 < _zz_dataOut_payload_0_14729);
  assign _zz_dataOut_payload_0_14736 = (_zz_dataOut_payload_0_14714 < _zz_dataOut_payload_0_14720);
  assign _zz_dataOut_payload_0_14737 = (_zz_dataOut_payload_0_14736 ? _zz_dataOut_payload_0_14714 : _zz_dataOut_payload_0_14720);
  assign _zz_dataOut_payload_0_14738 = (_zz_dataOut_payload_0_14736 ? _zz_dataOut_payload_0_14720 : _zz_dataOut_payload_0_14714);
  assign _zz_dataOut_payload_0_14739 = (_zz_dataOut_payload_0_14717 < _zz_dataOut_payload_0_14723);
  assign _zz_dataOut_payload_0_14740 = (_zz_dataOut_payload_0_14739 ? _zz_dataOut_payload_0_14717 : _zz_dataOut_payload_0_14723);
  assign _zz_dataOut_payload_0_14741 = (_zz_dataOut_payload_0_14739 ? _zz_dataOut_payload_0_14723 : _zz_dataOut_payload_0_14717);
  assign _zz_dataOut_payload_0_14742 = (_zz_dataOut_payload_0_14737 < _zz_dataOut_payload_0_14740);
  assign _zz_dataOut_payload_0_14743 = (_zz_dataOut_payload_0_14738 < _zz_dataOut_payload_0_14741);
  assign _zz_dataOut_payload_0_14756 = (_zz_dataOut_payload_0_14690 < _zz_dataOut_payload_0_14702);
  assign _zz_dataOut_payload_0_14757 = (_zz_dataOut_payload_0_14756 ? _zz_dataOut_payload_0_14690 : _zz_dataOut_payload_0_14702);
  assign _zz_dataOut_payload_0_14758 = (_zz_dataOut_payload_0_14756 ? _zz_dataOut_payload_0_14702 : _zz_dataOut_payload_0_14690);
  assign _zz_dataOut_payload_0_14759 = (_zz_dataOut_payload_0_14693 < _zz_dataOut_payload_0_14705);
  assign _zz_dataOut_payload_0_14760 = (_zz_dataOut_payload_0_14759 ? _zz_dataOut_payload_0_14693 : _zz_dataOut_payload_0_14705);
  assign _zz_dataOut_payload_0_14761 = (_zz_dataOut_payload_0_14759 ? _zz_dataOut_payload_0_14705 : _zz_dataOut_payload_0_14693);
  assign _zz_dataOut_payload_0_14762 = (_zz_dataOut_payload_0_14696 < _zz_dataOut_payload_0_14708);
  assign _zz_dataOut_payload_0_14763 = (_zz_dataOut_payload_0_14762 ? _zz_dataOut_payload_0_14696 : _zz_dataOut_payload_0_14708);
  assign _zz_dataOut_payload_0_14764 = (_zz_dataOut_payload_0_14762 ? _zz_dataOut_payload_0_14708 : _zz_dataOut_payload_0_14696);
  assign _zz_dataOut_payload_0_14765 = (_zz_dataOut_payload_0_14699 < _zz_dataOut_payload_0_14711);
  assign _zz_dataOut_payload_0_14766 = (_zz_dataOut_payload_0_14765 ? _zz_dataOut_payload_0_14699 : _zz_dataOut_payload_0_14711);
  assign _zz_dataOut_payload_0_14767 = (_zz_dataOut_payload_0_14765 ? _zz_dataOut_payload_0_14711 : _zz_dataOut_payload_0_14699);
  assign _zz_dataOut_payload_0_14768 = (_zz_dataOut_payload_0_14757 < _zz_dataOut_payload_0_14763);
  assign _zz_dataOut_payload_0_14769 = (_zz_dataOut_payload_0_14768 ? _zz_dataOut_payload_0_14757 : _zz_dataOut_payload_0_14763);
  assign _zz_dataOut_payload_0_14770 = (_zz_dataOut_payload_0_14768 ? _zz_dataOut_payload_0_14763 : _zz_dataOut_payload_0_14757);
  assign _zz_dataOut_payload_0_14771 = (_zz_dataOut_payload_0_14760 < _zz_dataOut_payload_0_14766);
  assign _zz_dataOut_payload_0_14772 = (_zz_dataOut_payload_0_14771 ? _zz_dataOut_payload_0_14760 : _zz_dataOut_payload_0_14766);
  assign _zz_dataOut_payload_0_14773 = (_zz_dataOut_payload_0_14771 ? _zz_dataOut_payload_0_14766 : _zz_dataOut_payload_0_14760);
  assign _zz_dataOut_payload_0_14774 = (_zz_dataOut_payload_0_14769 < _zz_dataOut_payload_0_14772);
  assign _zz_dataOut_payload_0_14775 = (_zz_dataOut_payload_0_14770 < _zz_dataOut_payload_0_14773);
  assign _zz_dataOut_payload_0_14780 = (_zz_dataOut_payload_0_14758 < _zz_dataOut_payload_0_14764);
  assign _zz_dataOut_payload_0_14781 = (_zz_dataOut_payload_0_14780 ? _zz_dataOut_payload_0_14758 : _zz_dataOut_payload_0_14764);
  assign _zz_dataOut_payload_0_14782 = (_zz_dataOut_payload_0_14780 ? _zz_dataOut_payload_0_14764 : _zz_dataOut_payload_0_14758);
  assign _zz_dataOut_payload_0_14783 = (_zz_dataOut_payload_0_14761 < _zz_dataOut_payload_0_14767);
  assign _zz_dataOut_payload_0_14784 = (_zz_dataOut_payload_0_14783 ? _zz_dataOut_payload_0_14761 : _zz_dataOut_payload_0_14767);
  assign _zz_dataOut_payload_0_14785 = (_zz_dataOut_payload_0_14783 ? _zz_dataOut_payload_0_14767 : _zz_dataOut_payload_0_14761);
  assign _zz_dataOut_payload_0_14786 = (_zz_dataOut_payload_0_14781 < _zz_dataOut_payload_0_14784);
  assign _zz_dataOut_payload_0_14787 = (_zz_dataOut_payload_0_14782 < _zz_dataOut_payload_0_14785);
  assign _zz_dataOut_payload_0_14912 = (_zz_dataOut_payload_0_14079 < _zz_dataOut_payload_0_13983);
  assign _zz_dataOut_payload_0_14913 = (_zz_dataOut_payload_0_14912 ? _zz_dataOut_payload_0_14079 : _zz_dataOut_payload_0_13983);
  assign _zz_dataOut_payload_0_14914 = (_zz_dataOut_payload_0_14912 ? _zz_dataOut_payload_0_13983 : _zz_dataOut_payload_0_14079);
  assign _zz_dataOut_payload_0_14915 = (_zz_dataOut_payload_0_14076 < _zz_dataOut_payload_0_13980);
  assign _zz_dataOut_payload_0_14916 = (_zz_dataOut_payload_0_14915 ? _zz_dataOut_payload_0_14076 : _zz_dataOut_payload_0_13980);
  assign _zz_dataOut_payload_0_14917 = (_zz_dataOut_payload_0_14915 ? _zz_dataOut_payload_0_13980 : _zz_dataOut_payload_0_14076);
  assign _zz_dataOut_payload_0_14918 = (_zz_dataOut_payload_0_14073 < _zz_dataOut_payload_0_13977);
  assign _zz_dataOut_payload_0_14919 = (_zz_dataOut_payload_0_14918 ? _zz_dataOut_payload_0_14073 : _zz_dataOut_payload_0_13977);
  assign _zz_dataOut_payload_0_14920 = (_zz_dataOut_payload_0_14918 ? _zz_dataOut_payload_0_13977 : _zz_dataOut_payload_0_14073);
  assign _zz_dataOut_payload_0_14921 = (_zz_dataOut_payload_0_14070 < _zz_dataOut_payload_0_13974);
  assign _zz_dataOut_payload_0_14922 = (_zz_dataOut_payload_0_14921 ? _zz_dataOut_payload_0_14070 : _zz_dataOut_payload_0_13974);
  assign _zz_dataOut_payload_0_14923 = (_zz_dataOut_payload_0_14921 ? _zz_dataOut_payload_0_13974 : _zz_dataOut_payload_0_14070);
  assign _zz_dataOut_payload_0_14924 = (_zz_dataOut_payload_0_14067 < _zz_dataOut_payload_0_13971);
  assign _zz_dataOut_payload_0_14925 = (_zz_dataOut_payload_0_14924 ? _zz_dataOut_payload_0_14067 : _zz_dataOut_payload_0_13971);
  assign _zz_dataOut_payload_0_14926 = (_zz_dataOut_payload_0_14924 ? _zz_dataOut_payload_0_13971 : _zz_dataOut_payload_0_14067);
  assign _zz_dataOut_payload_0_14927 = (_zz_dataOut_payload_0_14064 < _zz_dataOut_payload_0_13968);
  assign _zz_dataOut_payload_0_14928 = (_zz_dataOut_payload_0_14927 ? _zz_dataOut_payload_0_14064 : _zz_dataOut_payload_0_13968);
  assign _zz_dataOut_payload_0_14929 = (_zz_dataOut_payload_0_14927 ? _zz_dataOut_payload_0_13968 : _zz_dataOut_payload_0_14064);
  assign _zz_dataOut_payload_0_14930 = (_zz_dataOut_payload_0_14061 < _zz_dataOut_payload_0_13965);
  assign _zz_dataOut_payload_0_14931 = (_zz_dataOut_payload_0_14930 ? _zz_dataOut_payload_0_14061 : _zz_dataOut_payload_0_13965);
  assign _zz_dataOut_payload_0_14932 = (_zz_dataOut_payload_0_14930 ? _zz_dataOut_payload_0_13965 : _zz_dataOut_payload_0_14061);
  assign _zz_dataOut_payload_0_14933 = (_zz_dataOut_payload_0_14058 < _zz_dataOut_payload_0_13962);
  assign _zz_dataOut_payload_0_14934 = (_zz_dataOut_payload_0_14933 ? _zz_dataOut_payload_0_14058 : _zz_dataOut_payload_0_13962);
  assign _zz_dataOut_payload_0_14935 = (_zz_dataOut_payload_0_14933 ? _zz_dataOut_payload_0_13962 : _zz_dataOut_payload_0_14058);
  assign _zz_dataOut_payload_0_14936 = (_zz_dataOut_payload_0_14055 < _zz_dataOut_payload_0_13959);
  assign _zz_dataOut_payload_0_14937 = (_zz_dataOut_payload_0_14936 ? _zz_dataOut_payload_0_14055 : _zz_dataOut_payload_0_13959);
  assign _zz_dataOut_payload_0_14938 = (_zz_dataOut_payload_0_14936 ? _zz_dataOut_payload_0_13959 : _zz_dataOut_payload_0_14055);
  assign _zz_dataOut_payload_0_14939 = (_zz_dataOut_payload_0_14052 < _zz_dataOut_payload_0_13956);
  assign _zz_dataOut_payload_0_14940 = (_zz_dataOut_payload_0_14939 ? _zz_dataOut_payload_0_14052 : _zz_dataOut_payload_0_13956);
  assign _zz_dataOut_payload_0_14941 = (_zz_dataOut_payload_0_14939 ? _zz_dataOut_payload_0_13956 : _zz_dataOut_payload_0_14052);
  assign _zz_dataOut_payload_0_14942 = (_zz_dataOut_payload_0_14049 < _zz_dataOut_payload_0_13953);
  assign _zz_dataOut_payload_0_14943 = (_zz_dataOut_payload_0_14942 ? _zz_dataOut_payload_0_14049 : _zz_dataOut_payload_0_13953);
  assign _zz_dataOut_payload_0_14944 = (_zz_dataOut_payload_0_14942 ? _zz_dataOut_payload_0_13953 : _zz_dataOut_payload_0_14049);
  assign _zz_dataOut_payload_0_14945 = (_zz_dataOut_payload_0_14046 < _zz_dataOut_payload_0_13950);
  assign _zz_dataOut_payload_0_14946 = (_zz_dataOut_payload_0_14945 ? _zz_dataOut_payload_0_14046 : _zz_dataOut_payload_0_13950);
  assign _zz_dataOut_payload_0_14947 = (_zz_dataOut_payload_0_14945 ? _zz_dataOut_payload_0_13950 : _zz_dataOut_payload_0_14046);
  assign _zz_dataOut_payload_0_14948 = (_zz_dataOut_payload_0_14043 < _zz_dataOut_payload_0_13947);
  assign _zz_dataOut_payload_0_14949 = (_zz_dataOut_payload_0_14948 ? _zz_dataOut_payload_0_14043 : _zz_dataOut_payload_0_13947);
  assign _zz_dataOut_payload_0_14950 = (_zz_dataOut_payload_0_14948 ? _zz_dataOut_payload_0_13947 : _zz_dataOut_payload_0_14043);
  assign _zz_dataOut_payload_0_14951 = (_zz_dataOut_payload_0_14040 < _zz_dataOut_payload_0_13944);
  assign _zz_dataOut_payload_0_14952 = (_zz_dataOut_payload_0_14951 ? _zz_dataOut_payload_0_14040 : _zz_dataOut_payload_0_13944);
  assign _zz_dataOut_payload_0_14953 = (_zz_dataOut_payload_0_14951 ? _zz_dataOut_payload_0_13944 : _zz_dataOut_payload_0_14040);
  assign _zz_dataOut_payload_0_14954 = (_zz_dataOut_payload_0_14037 < _zz_dataOut_payload_0_13941);
  assign _zz_dataOut_payload_0_14955 = (_zz_dataOut_payload_0_14954 ? _zz_dataOut_payload_0_14037 : _zz_dataOut_payload_0_13941);
  assign _zz_dataOut_payload_0_14956 = (_zz_dataOut_payload_0_14954 ? _zz_dataOut_payload_0_13941 : _zz_dataOut_payload_0_14037);
  assign _zz_dataOut_payload_0_14957 = (_zz_dataOut_payload_0_14034 < _zz_dataOut_payload_0_13938);
  assign _zz_dataOut_payload_0_14958 = (_zz_dataOut_payload_0_14957 ? _zz_dataOut_payload_0_14034 : _zz_dataOut_payload_0_13938);
  assign _zz_dataOut_payload_0_14959 = (_zz_dataOut_payload_0_14957 ? _zz_dataOut_payload_0_13938 : _zz_dataOut_payload_0_14034);
  assign _zz_dataOut_payload_0_14960 = (_zz_dataOut_payload_0_14031 < _zz_dataOut_payload_0_13935);
  assign _zz_dataOut_payload_0_14961 = (_zz_dataOut_payload_0_14960 ? _zz_dataOut_payload_0_14031 : _zz_dataOut_payload_0_13935);
  assign _zz_dataOut_payload_0_14962 = (_zz_dataOut_payload_0_14960 ? _zz_dataOut_payload_0_13935 : _zz_dataOut_payload_0_14031);
  assign _zz_dataOut_payload_0_14963 = (_zz_dataOut_payload_0_14028 < _zz_dataOut_payload_0_13932);
  assign _zz_dataOut_payload_0_14964 = (_zz_dataOut_payload_0_14963 ? _zz_dataOut_payload_0_14028 : _zz_dataOut_payload_0_13932);
  assign _zz_dataOut_payload_0_14965 = (_zz_dataOut_payload_0_14963 ? _zz_dataOut_payload_0_13932 : _zz_dataOut_payload_0_14028);
  assign _zz_dataOut_payload_0_14966 = (_zz_dataOut_payload_0_14025 < _zz_dataOut_payload_0_13929);
  assign _zz_dataOut_payload_0_14967 = (_zz_dataOut_payload_0_14966 ? _zz_dataOut_payload_0_14025 : _zz_dataOut_payload_0_13929);
  assign _zz_dataOut_payload_0_14968 = (_zz_dataOut_payload_0_14966 ? _zz_dataOut_payload_0_13929 : _zz_dataOut_payload_0_14025);
  assign _zz_dataOut_payload_0_14969 = (_zz_dataOut_payload_0_14022 < _zz_dataOut_payload_0_13926);
  assign _zz_dataOut_payload_0_14970 = (_zz_dataOut_payload_0_14969 ? _zz_dataOut_payload_0_14022 : _zz_dataOut_payload_0_13926);
  assign _zz_dataOut_payload_0_14971 = (_zz_dataOut_payload_0_14969 ? _zz_dataOut_payload_0_13926 : _zz_dataOut_payload_0_14022);
  assign _zz_dataOut_payload_0_14972 = (_zz_dataOut_payload_0_14019 < _zz_dataOut_payload_0_13923);
  assign _zz_dataOut_payload_0_14973 = (_zz_dataOut_payload_0_14972 ? _zz_dataOut_payload_0_14019 : _zz_dataOut_payload_0_13923);
  assign _zz_dataOut_payload_0_14974 = (_zz_dataOut_payload_0_14972 ? _zz_dataOut_payload_0_13923 : _zz_dataOut_payload_0_14019);
  assign _zz_dataOut_payload_0_14975 = (_zz_dataOut_payload_0_14016 < _zz_dataOut_payload_0_13920);
  assign _zz_dataOut_payload_0_14976 = (_zz_dataOut_payload_0_14975 ? _zz_dataOut_payload_0_14016 : _zz_dataOut_payload_0_13920);
  assign _zz_dataOut_payload_0_14977 = (_zz_dataOut_payload_0_14975 ? _zz_dataOut_payload_0_13920 : _zz_dataOut_payload_0_14016);
  assign _zz_dataOut_payload_0_14978 = (_zz_dataOut_payload_0_14013 < _zz_dataOut_payload_0_13917);
  assign _zz_dataOut_payload_0_14979 = (_zz_dataOut_payload_0_14978 ? _zz_dataOut_payload_0_14013 : _zz_dataOut_payload_0_13917);
  assign _zz_dataOut_payload_0_14980 = (_zz_dataOut_payload_0_14978 ? _zz_dataOut_payload_0_13917 : _zz_dataOut_payload_0_14013);
  assign _zz_dataOut_payload_0_14981 = (_zz_dataOut_payload_0_14010 < _zz_dataOut_payload_0_13914);
  assign _zz_dataOut_payload_0_14982 = (_zz_dataOut_payload_0_14981 ? _zz_dataOut_payload_0_14010 : _zz_dataOut_payload_0_13914);
  assign _zz_dataOut_payload_0_14983 = (_zz_dataOut_payload_0_14981 ? _zz_dataOut_payload_0_13914 : _zz_dataOut_payload_0_14010);
  assign _zz_dataOut_payload_0_14984 = (_zz_dataOut_payload_0_14007 < _zz_dataOut_payload_0_13911);
  assign _zz_dataOut_payload_0_14985 = (_zz_dataOut_payload_0_14984 ? _zz_dataOut_payload_0_14007 : _zz_dataOut_payload_0_13911);
  assign _zz_dataOut_payload_0_14986 = (_zz_dataOut_payload_0_14984 ? _zz_dataOut_payload_0_13911 : _zz_dataOut_payload_0_14007);
  assign _zz_dataOut_payload_0_14987 = (_zz_dataOut_payload_0_14004 < _zz_dataOut_payload_0_13908);
  assign _zz_dataOut_payload_0_14988 = (_zz_dataOut_payload_0_14987 ? _zz_dataOut_payload_0_14004 : _zz_dataOut_payload_0_13908);
  assign _zz_dataOut_payload_0_14989 = (_zz_dataOut_payload_0_14987 ? _zz_dataOut_payload_0_13908 : _zz_dataOut_payload_0_14004);
  assign _zz_dataOut_payload_0_14990 = (_zz_dataOut_payload_0_14001 < _zz_dataOut_payload_0_13905);
  assign _zz_dataOut_payload_0_14991 = (_zz_dataOut_payload_0_14990 ? _zz_dataOut_payload_0_14001 : _zz_dataOut_payload_0_13905);
  assign _zz_dataOut_payload_0_14992 = (_zz_dataOut_payload_0_14990 ? _zz_dataOut_payload_0_13905 : _zz_dataOut_payload_0_14001);
  assign _zz_dataOut_payload_0_14993 = (_zz_dataOut_payload_0_13998 < _zz_dataOut_payload_0_13902);
  assign _zz_dataOut_payload_0_14994 = (_zz_dataOut_payload_0_14993 ? _zz_dataOut_payload_0_13998 : _zz_dataOut_payload_0_13902);
  assign _zz_dataOut_payload_0_14995 = (_zz_dataOut_payload_0_14993 ? _zz_dataOut_payload_0_13902 : _zz_dataOut_payload_0_13998);
  assign _zz_dataOut_payload_0_14996 = (_zz_dataOut_payload_0_13995 < _zz_dataOut_payload_0_13899);
  assign _zz_dataOut_payload_0_14997 = (_zz_dataOut_payload_0_14996 ? _zz_dataOut_payload_0_13995 : _zz_dataOut_payload_0_13899);
  assign _zz_dataOut_payload_0_14998 = (_zz_dataOut_payload_0_14996 ? _zz_dataOut_payload_0_13899 : _zz_dataOut_payload_0_13995);
  assign _zz_dataOut_payload_0_14999 = (_zz_dataOut_payload_0_13992 < _zz_dataOut_payload_0_13896);
  assign _zz_dataOut_payload_0_15000 = (_zz_dataOut_payload_0_14999 ? _zz_dataOut_payload_0_13992 : _zz_dataOut_payload_0_13896);
  assign _zz_dataOut_payload_0_15001 = (_zz_dataOut_payload_0_14999 ? _zz_dataOut_payload_0_13896 : _zz_dataOut_payload_0_13992);
  assign _zz_dataOut_payload_0_15002 = (_zz_dataOut_payload_0_13989 < _zz_dataOut_payload_0_13893);
  assign _zz_dataOut_payload_0_15003 = (_zz_dataOut_payload_0_15002 ? _zz_dataOut_payload_0_13989 : _zz_dataOut_payload_0_13893);
  assign _zz_dataOut_payload_0_15004 = (_zz_dataOut_payload_0_15002 ? _zz_dataOut_payload_0_13893 : _zz_dataOut_payload_0_13989);
  assign _zz_dataOut_payload_0_15005 = (_zz_dataOut_payload_0_13986 < _zz_dataOut_payload_0_13890);
  assign _zz_dataOut_payload_0_15006 = (_zz_dataOut_payload_0_15005 ? _zz_dataOut_payload_0_13986 : _zz_dataOut_payload_0_13890);
  assign _zz_dataOut_payload_0_15007 = (_zz_dataOut_payload_0_15005 ? _zz_dataOut_payload_0_13890 : _zz_dataOut_payload_0_13986);
  assign _zz_dataOut_payload_0_15008 = (_zz_dataOut_payload_0_14913 < _zz_dataOut_payload_0_14961);
  assign _zz_dataOut_payload_0_15009 = (_zz_dataOut_payload_0_15008 ? _zz_dataOut_payload_0_14913 : _zz_dataOut_payload_0_14961);
  assign _zz_dataOut_payload_0_15010 = (_zz_dataOut_payload_0_15008 ? _zz_dataOut_payload_0_14961 : _zz_dataOut_payload_0_14913);
  assign _zz_dataOut_payload_0_15011 = (_zz_dataOut_payload_0_14916 < _zz_dataOut_payload_0_14964);
  assign _zz_dataOut_payload_0_15012 = (_zz_dataOut_payload_0_15011 ? _zz_dataOut_payload_0_14916 : _zz_dataOut_payload_0_14964);
  assign _zz_dataOut_payload_0_15013 = (_zz_dataOut_payload_0_15011 ? _zz_dataOut_payload_0_14964 : _zz_dataOut_payload_0_14916);
  assign _zz_dataOut_payload_0_15014 = (_zz_dataOut_payload_0_14919 < _zz_dataOut_payload_0_14967);
  assign _zz_dataOut_payload_0_15015 = (_zz_dataOut_payload_0_15014 ? _zz_dataOut_payload_0_14919 : _zz_dataOut_payload_0_14967);
  assign _zz_dataOut_payload_0_15016 = (_zz_dataOut_payload_0_15014 ? _zz_dataOut_payload_0_14967 : _zz_dataOut_payload_0_14919);
  assign _zz_dataOut_payload_0_15017 = (_zz_dataOut_payload_0_14922 < _zz_dataOut_payload_0_14970);
  assign _zz_dataOut_payload_0_15018 = (_zz_dataOut_payload_0_15017 ? _zz_dataOut_payload_0_14922 : _zz_dataOut_payload_0_14970);
  assign _zz_dataOut_payload_0_15019 = (_zz_dataOut_payload_0_15017 ? _zz_dataOut_payload_0_14970 : _zz_dataOut_payload_0_14922);
  assign _zz_dataOut_payload_0_15020 = (_zz_dataOut_payload_0_14925 < _zz_dataOut_payload_0_14973);
  assign _zz_dataOut_payload_0_15021 = (_zz_dataOut_payload_0_15020 ? _zz_dataOut_payload_0_14925 : _zz_dataOut_payload_0_14973);
  assign _zz_dataOut_payload_0_15022 = (_zz_dataOut_payload_0_15020 ? _zz_dataOut_payload_0_14973 : _zz_dataOut_payload_0_14925);
  assign _zz_dataOut_payload_0_15023 = (_zz_dataOut_payload_0_14928 < _zz_dataOut_payload_0_14976);
  assign _zz_dataOut_payload_0_15024 = (_zz_dataOut_payload_0_15023 ? _zz_dataOut_payload_0_14928 : _zz_dataOut_payload_0_14976);
  assign _zz_dataOut_payload_0_15025 = (_zz_dataOut_payload_0_15023 ? _zz_dataOut_payload_0_14976 : _zz_dataOut_payload_0_14928);
  assign _zz_dataOut_payload_0_15026 = (_zz_dataOut_payload_0_14931 < _zz_dataOut_payload_0_14979);
  assign _zz_dataOut_payload_0_15027 = (_zz_dataOut_payload_0_15026 ? _zz_dataOut_payload_0_14931 : _zz_dataOut_payload_0_14979);
  assign _zz_dataOut_payload_0_15028 = (_zz_dataOut_payload_0_15026 ? _zz_dataOut_payload_0_14979 : _zz_dataOut_payload_0_14931);
  assign _zz_dataOut_payload_0_15029 = (_zz_dataOut_payload_0_14934 < _zz_dataOut_payload_0_14982);
  assign _zz_dataOut_payload_0_15030 = (_zz_dataOut_payload_0_15029 ? _zz_dataOut_payload_0_14934 : _zz_dataOut_payload_0_14982);
  assign _zz_dataOut_payload_0_15031 = (_zz_dataOut_payload_0_15029 ? _zz_dataOut_payload_0_14982 : _zz_dataOut_payload_0_14934);
  assign _zz_dataOut_payload_0_15032 = (_zz_dataOut_payload_0_14937 < _zz_dataOut_payload_0_14985);
  assign _zz_dataOut_payload_0_15033 = (_zz_dataOut_payload_0_15032 ? _zz_dataOut_payload_0_14937 : _zz_dataOut_payload_0_14985);
  assign _zz_dataOut_payload_0_15034 = (_zz_dataOut_payload_0_15032 ? _zz_dataOut_payload_0_14985 : _zz_dataOut_payload_0_14937);
  assign _zz_dataOut_payload_0_15035 = (_zz_dataOut_payload_0_14940 < _zz_dataOut_payload_0_14988);
  assign _zz_dataOut_payload_0_15036 = (_zz_dataOut_payload_0_15035 ? _zz_dataOut_payload_0_14940 : _zz_dataOut_payload_0_14988);
  assign _zz_dataOut_payload_0_15037 = (_zz_dataOut_payload_0_15035 ? _zz_dataOut_payload_0_14988 : _zz_dataOut_payload_0_14940);
  assign _zz_dataOut_payload_0_15038 = (_zz_dataOut_payload_0_14943 < _zz_dataOut_payload_0_14991);
  assign _zz_dataOut_payload_0_15039 = (_zz_dataOut_payload_0_15038 ? _zz_dataOut_payload_0_14943 : _zz_dataOut_payload_0_14991);
  assign _zz_dataOut_payload_0_15040 = (_zz_dataOut_payload_0_15038 ? _zz_dataOut_payload_0_14991 : _zz_dataOut_payload_0_14943);
  assign _zz_dataOut_payload_0_15041 = (_zz_dataOut_payload_0_14946 < _zz_dataOut_payload_0_14994);
  assign _zz_dataOut_payload_0_15042 = (_zz_dataOut_payload_0_15041 ? _zz_dataOut_payload_0_14946 : _zz_dataOut_payload_0_14994);
  assign _zz_dataOut_payload_0_15043 = (_zz_dataOut_payload_0_15041 ? _zz_dataOut_payload_0_14994 : _zz_dataOut_payload_0_14946);
  assign _zz_dataOut_payload_0_15044 = (_zz_dataOut_payload_0_14949 < _zz_dataOut_payload_0_14997);
  assign _zz_dataOut_payload_0_15045 = (_zz_dataOut_payload_0_15044 ? _zz_dataOut_payload_0_14949 : _zz_dataOut_payload_0_14997);
  assign _zz_dataOut_payload_0_15046 = (_zz_dataOut_payload_0_15044 ? _zz_dataOut_payload_0_14997 : _zz_dataOut_payload_0_14949);
  assign _zz_dataOut_payload_0_15047 = (_zz_dataOut_payload_0_14952 < _zz_dataOut_payload_0_15000);
  assign _zz_dataOut_payload_0_15048 = (_zz_dataOut_payload_0_15047 ? _zz_dataOut_payload_0_14952 : _zz_dataOut_payload_0_15000);
  assign _zz_dataOut_payload_0_15049 = (_zz_dataOut_payload_0_15047 ? _zz_dataOut_payload_0_15000 : _zz_dataOut_payload_0_14952);
  assign _zz_dataOut_payload_0_15050 = (_zz_dataOut_payload_0_14955 < _zz_dataOut_payload_0_15003);
  assign _zz_dataOut_payload_0_15051 = (_zz_dataOut_payload_0_15050 ? _zz_dataOut_payload_0_14955 : _zz_dataOut_payload_0_15003);
  assign _zz_dataOut_payload_0_15052 = (_zz_dataOut_payload_0_15050 ? _zz_dataOut_payload_0_15003 : _zz_dataOut_payload_0_14955);
  assign _zz_dataOut_payload_0_15053 = (_zz_dataOut_payload_0_14958 < _zz_dataOut_payload_0_15006);
  assign _zz_dataOut_payload_0_15054 = (_zz_dataOut_payload_0_15053 ? _zz_dataOut_payload_0_14958 : _zz_dataOut_payload_0_15006);
  assign _zz_dataOut_payload_0_15055 = (_zz_dataOut_payload_0_15053 ? _zz_dataOut_payload_0_15006 : _zz_dataOut_payload_0_14958);
  assign _zz_dataOut_payload_0_15056 = (_zz_dataOut_payload_0_15009 < _zz_dataOut_payload_0_15033);
  assign _zz_dataOut_payload_0_15057 = (_zz_dataOut_payload_0_15056 ? _zz_dataOut_payload_0_15009 : _zz_dataOut_payload_0_15033);
  assign _zz_dataOut_payload_0_15058 = (_zz_dataOut_payload_0_15056 ? _zz_dataOut_payload_0_15033 : _zz_dataOut_payload_0_15009);
  assign _zz_dataOut_payload_0_15059 = (_zz_dataOut_payload_0_15012 < _zz_dataOut_payload_0_15036);
  assign _zz_dataOut_payload_0_15060 = (_zz_dataOut_payload_0_15059 ? _zz_dataOut_payload_0_15012 : _zz_dataOut_payload_0_15036);
  assign _zz_dataOut_payload_0_15061 = (_zz_dataOut_payload_0_15059 ? _zz_dataOut_payload_0_15036 : _zz_dataOut_payload_0_15012);
  assign _zz_dataOut_payload_0_15062 = (_zz_dataOut_payload_0_15015 < _zz_dataOut_payload_0_15039);
  assign _zz_dataOut_payload_0_15063 = (_zz_dataOut_payload_0_15062 ? _zz_dataOut_payload_0_15015 : _zz_dataOut_payload_0_15039);
  assign _zz_dataOut_payload_0_15064 = (_zz_dataOut_payload_0_15062 ? _zz_dataOut_payload_0_15039 : _zz_dataOut_payload_0_15015);
  assign _zz_dataOut_payload_0_15065 = (_zz_dataOut_payload_0_15018 < _zz_dataOut_payload_0_15042);
  assign _zz_dataOut_payload_0_15066 = (_zz_dataOut_payload_0_15065 ? _zz_dataOut_payload_0_15018 : _zz_dataOut_payload_0_15042);
  assign _zz_dataOut_payload_0_15067 = (_zz_dataOut_payload_0_15065 ? _zz_dataOut_payload_0_15042 : _zz_dataOut_payload_0_15018);
  assign _zz_dataOut_payload_0_15068 = (_zz_dataOut_payload_0_15021 < _zz_dataOut_payload_0_15045);
  assign _zz_dataOut_payload_0_15069 = (_zz_dataOut_payload_0_15068 ? _zz_dataOut_payload_0_15021 : _zz_dataOut_payload_0_15045);
  assign _zz_dataOut_payload_0_15070 = (_zz_dataOut_payload_0_15068 ? _zz_dataOut_payload_0_15045 : _zz_dataOut_payload_0_15021);
  assign _zz_dataOut_payload_0_15071 = (_zz_dataOut_payload_0_15024 < _zz_dataOut_payload_0_15048);
  assign _zz_dataOut_payload_0_15072 = (_zz_dataOut_payload_0_15071 ? _zz_dataOut_payload_0_15024 : _zz_dataOut_payload_0_15048);
  assign _zz_dataOut_payload_0_15073 = (_zz_dataOut_payload_0_15071 ? _zz_dataOut_payload_0_15048 : _zz_dataOut_payload_0_15024);
  assign _zz_dataOut_payload_0_15074 = (_zz_dataOut_payload_0_15027 < _zz_dataOut_payload_0_15051);
  assign _zz_dataOut_payload_0_15075 = (_zz_dataOut_payload_0_15074 ? _zz_dataOut_payload_0_15027 : _zz_dataOut_payload_0_15051);
  assign _zz_dataOut_payload_0_15076 = (_zz_dataOut_payload_0_15074 ? _zz_dataOut_payload_0_15051 : _zz_dataOut_payload_0_15027);
  assign _zz_dataOut_payload_0_15077 = (_zz_dataOut_payload_0_15030 < _zz_dataOut_payload_0_15054);
  assign _zz_dataOut_payload_0_15078 = (_zz_dataOut_payload_0_15077 ? _zz_dataOut_payload_0_15030 : _zz_dataOut_payload_0_15054);
  assign _zz_dataOut_payload_0_15079 = (_zz_dataOut_payload_0_15077 ? _zz_dataOut_payload_0_15054 : _zz_dataOut_payload_0_15030);
  assign _zz_dataOut_payload_0_15080 = (_zz_dataOut_payload_0_15057 < _zz_dataOut_payload_0_15069);
  assign _zz_dataOut_payload_0_15081 = (_zz_dataOut_payload_0_15080 ? _zz_dataOut_payload_0_15057 : _zz_dataOut_payload_0_15069);
  assign _zz_dataOut_payload_0_15082 = (_zz_dataOut_payload_0_15080 ? _zz_dataOut_payload_0_15069 : _zz_dataOut_payload_0_15057);
  assign _zz_dataOut_payload_0_15083 = (_zz_dataOut_payload_0_15060 < _zz_dataOut_payload_0_15072);
  assign _zz_dataOut_payload_0_15084 = (_zz_dataOut_payload_0_15083 ? _zz_dataOut_payload_0_15060 : _zz_dataOut_payload_0_15072);
  assign _zz_dataOut_payload_0_15085 = (_zz_dataOut_payload_0_15083 ? _zz_dataOut_payload_0_15072 : _zz_dataOut_payload_0_15060);
  assign _zz_dataOut_payload_0_15086 = (_zz_dataOut_payload_0_15063 < _zz_dataOut_payload_0_15075);
  assign _zz_dataOut_payload_0_15087 = (_zz_dataOut_payload_0_15086 ? _zz_dataOut_payload_0_15063 : _zz_dataOut_payload_0_15075);
  assign _zz_dataOut_payload_0_15088 = (_zz_dataOut_payload_0_15086 ? _zz_dataOut_payload_0_15075 : _zz_dataOut_payload_0_15063);
  assign _zz_dataOut_payload_0_15089 = (_zz_dataOut_payload_0_15066 < _zz_dataOut_payload_0_15078);
  assign _zz_dataOut_payload_0_15090 = (_zz_dataOut_payload_0_15089 ? _zz_dataOut_payload_0_15066 : _zz_dataOut_payload_0_15078);
  assign _zz_dataOut_payload_0_15091 = (_zz_dataOut_payload_0_15089 ? _zz_dataOut_payload_0_15078 : _zz_dataOut_payload_0_15066);
  assign _zz_dataOut_payload_0_15092 = (_zz_dataOut_payload_0_15081 < _zz_dataOut_payload_0_15087);
  assign _zz_dataOut_payload_0_15093 = (_zz_dataOut_payload_0_15092 ? _zz_dataOut_payload_0_15081 : _zz_dataOut_payload_0_15087);
  assign _zz_dataOut_payload_0_15094 = (_zz_dataOut_payload_0_15092 ? _zz_dataOut_payload_0_15087 : _zz_dataOut_payload_0_15081);
  assign _zz_dataOut_payload_0_15095 = (_zz_dataOut_payload_0_15084 < _zz_dataOut_payload_0_15090);
  assign _zz_dataOut_payload_0_15096 = (_zz_dataOut_payload_0_15095 ? _zz_dataOut_payload_0_15084 : _zz_dataOut_payload_0_15090);
  assign _zz_dataOut_payload_0_15097 = (_zz_dataOut_payload_0_15095 ? _zz_dataOut_payload_0_15090 : _zz_dataOut_payload_0_15084);
  assign _zz_dataOut_payload_0_15098 = (_zz_dataOut_payload_0_15093 < _zz_dataOut_payload_0_15096);
  assign _zz_dataOut_payload_0_15099 = (_zz_dataOut_payload_0_15094 < _zz_dataOut_payload_0_15097);
  assign _zz_dataOut_payload_0_15104 = (_zz_dataOut_payload_0_15082 < _zz_dataOut_payload_0_15088);
  assign _zz_dataOut_payload_0_15105 = (_zz_dataOut_payload_0_15104 ? _zz_dataOut_payload_0_15082 : _zz_dataOut_payload_0_15088);
  assign _zz_dataOut_payload_0_15106 = (_zz_dataOut_payload_0_15104 ? _zz_dataOut_payload_0_15088 : _zz_dataOut_payload_0_15082);
  assign _zz_dataOut_payload_0_15107 = (_zz_dataOut_payload_0_15085 < _zz_dataOut_payload_0_15091);
  assign _zz_dataOut_payload_0_15108 = (_zz_dataOut_payload_0_15107 ? _zz_dataOut_payload_0_15085 : _zz_dataOut_payload_0_15091);
  assign _zz_dataOut_payload_0_15109 = (_zz_dataOut_payload_0_15107 ? _zz_dataOut_payload_0_15091 : _zz_dataOut_payload_0_15085);
  assign _zz_dataOut_payload_0_15110 = (_zz_dataOut_payload_0_15105 < _zz_dataOut_payload_0_15108);
  assign _zz_dataOut_payload_0_15111 = (_zz_dataOut_payload_0_15106 < _zz_dataOut_payload_0_15109);
  assign _zz_dataOut_payload_0_15124 = (_zz_dataOut_payload_0_15058 < _zz_dataOut_payload_0_15070);
  assign _zz_dataOut_payload_0_15125 = (_zz_dataOut_payload_0_15124 ? _zz_dataOut_payload_0_15058 : _zz_dataOut_payload_0_15070);
  assign _zz_dataOut_payload_0_15126 = (_zz_dataOut_payload_0_15124 ? _zz_dataOut_payload_0_15070 : _zz_dataOut_payload_0_15058);
  assign _zz_dataOut_payload_0_15127 = (_zz_dataOut_payload_0_15061 < _zz_dataOut_payload_0_15073);
  assign _zz_dataOut_payload_0_15128 = (_zz_dataOut_payload_0_15127 ? _zz_dataOut_payload_0_15061 : _zz_dataOut_payload_0_15073);
  assign _zz_dataOut_payload_0_15129 = (_zz_dataOut_payload_0_15127 ? _zz_dataOut_payload_0_15073 : _zz_dataOut_payload_0_15061);
  assign _zz_dataOut_payload_0_15130 = (_zz_dataOut_payload_0_15064 < _zz_dataOut_payload_0_15076);
  assign _zz_dataOut_payload_0_15131 = (_zz_dataOut_payload_0_15130 ? _zz_dataOut_payload_0_15064 : _zz_dataOut_payload_0_15076);
  assign _zz_dataOut_payload_0_15132 = (_zz_dataOut_payload_0_15130 ? _zz_dataOut_payload_0_15076 : _zz_dataOut_payload_0_15064);
  assign _zz_dataOut_payload_0_15133 = (_zz_dataOut_payload_0_15067 < _zz_dataOut_payload_0_15079);
  assign _zz_dataOut_payload_0_15134 = (_zz_dataOut_payload_0_15133 ? _zz_dataOut_payload_0_15067 : _zz_dataOut_payload_0_15079);
  assign _zz_dataOut_payload_0_15135 = (_zz_dataOut_payload_0_15133 ? _zz_dataOut_payload_0_15079 : _zz_dataOut_payload_0_15067);
  assign _zz_dataOut_payload_0_15136 = (_zz_dataOut_payload_0_15125 < _zz_dataOut_payload_0_15131);
  assign _zz_dataOut_payload_0_15137 = (_zz_dataOut_payload_0_15136 ? _zz_dataOut_payload_0_15125 : _zz_dataOut_payload_0_15131);
  assign _zz_dataOut_payload_0_15138 = (_zz_dataOut_payload_0_15136 ? _zz_dataOut_payload_0_15131 : _zz_dataOut_payload_0_15125);
  assign _zz_dataOut_payload_0_15139 = (_zz_dataOut_payload_0_15128 < _zz_dataOut_payload_0_15134);
  assign _zz_dataOut_payload_0_15140 = (_zz_dataOut_payload_0_15139 ? _zz_dataOut_payload_0_15128 : _zz_dataOut_payload_0_15134);
  assign _zz_dataOut_payload_0_15141 = (_zz_dataOut_payload_0_15139 ? _zz_dataOut_payload_0_15134 : _zz_dataOut_payload_0_15128);
  assign _zz_dataOut_payload_0_15142 = (_zz_dataOut_payload_0_15137 < _zz_dataOut_payload_0_15140);
  assign _zz_dataOut_payload_0_15143 = (_zz_dataOut_payload_0_15138 < _zz_dataOut_payload_0_15141);
  assign _zz_dataOut_payload_0_15148 = (_zz_dataOut_payload_0_15126 < _zz_dataOut_payload_0_15132);
  assign _zz_dataOut_payload_0_15149 = (_zz_dataOut_payload_0_15148 ? _zz_dataOut_payload_0_15126 : _zz_dataOut_payload_0_15132);
  assign _zz_dataOut_payload_0_15150 = (_zz_dataOut_payload_0_15148 ? _zz_dataOut_payload_0_15132 : _zz_dataOut_payload_0_15126);
  assign _zz_dataOut_payload_0_15151 = (_zz_dataOut_payload_0_15129 < _zz_dataOut_payload_0_15135);
  assign _zz_dataOut_payload_0_15152 = (_zz_dataOut_payload_0_15151 ? _zz_dataOut_payload_0_15129 : _zz_dataOut_payload_0_15135);
  assign _zz_dataOut_payload_0_15153 = (_zz_dataOut_payload_0_15151 ? _zz_dataOut_payload_0_15135 : _zz_dataOut_payload_0_15129);
  assign _zz_dataOut_payload_0_15154 = (_zz_dataOut_payload_0_15149 < _zz_dataOut_payload_0_15152);
  assign _zz_dataOut_payload_0_15155 = (_zz_dataOut_payload_0_15150 < _zz_dataOut_payload_0_15153);
  assign _zz_dataOut_payload_0_15184 = (_zz_dataOut_payload_0_15010 < _zz_dataOut_payload_0_15034);
  assign _zz_dataOut_payload_0_15185 = (_zz_dataOut_payload_0_15184 ? _zz_dataOut_payload_0_15010 : _zz_dataOut_payload_0_15034);
  assign _zz_dataOut_payload_0_15186 = (_zz_dataOut_payload_0_15184 ? _zz_dataOut_payload_0_15034 : _zz_dataOut_payload_0_15010);
  assign _zz_dataOut_payload_0_15187 = (_zz_dataOut_payload_0_15013 < _zz_dataOut_payload_0_15037);
  assign _zz_dataOut_payload_0_15188 = (_zz_dataOut_payload_0_15187 ? _zz_dataOut_payload_0_15013 : _zz_dataOut_payload_0_15037);
  assign _zz_dataOut_payload_0_15189 = (_zz_dataOut_payload_0_15187 ? _zz_dataOut_payload_0_15037 : _zz_dataOut_payload_0_15013);
  assign _zz_dataOut_payload_0_15190 = (_zz_dataOut_payload_0_15016 < _zz_dataOut_payload_0_15040);
  assign _zz_dataOut_payload_0_15191 = (_zz_dataOut_payload_0_15190 ? _zz_dataOut_payload_0_15016 : _zz_dataOut_payload_0_15040);
  assign _zz_dataOut_payload_0_15192 = (_zz_dataOut_payload_0_15190 ? _zz_dataOut_payload_0_15040 : _zz_dataOut_payload_0_15016);
  assign _zz_dataOut_payload_0_15193 = (_zz_dataOut_payload_0_15019 < _zz_dataOut_payload_0_15043);
  assign _zz_dataOut_payload_0_15194 = (_zz_dataOut_payload_0_15193 ? _zz_dataOut_payload_0_15019 : _zz_dataOut_payload_0_15043);
  assign _zz_dataOut_payload_0_15195 = (_zz_dataOut_payload_0_15193 ? _zz_dataOut_payload_0_15043 : _zz_dataOut_payload_0_15019);
  assign _zz_dataOut_payload_0_15196 = (_zz_dataOut_payload_0_15022 < _zz_dataOut_payload_0_15046);
  assign _zz_dataOut_payload_0_15197 = (_zz_dataOut_payload_0_15196 ? _zz_dataOut_payload_0_15022 : _zz_dataOut_payload_0_15046);
  assign _zz_dataOut_payload_0_15198 = (_zz_dataOut_payload_0_15196 ? _zz_dataOut_payload_0_15046 : _zz_dataOut_payload_0_15022);
  assign _zz_dataOut_payload_0_15199 = (_zz_dataOut_payload_0_15025 < _zz_dataOut_payload_0_15049);
  assign _zz_dataOut_payload_0_15200 = (_zz_dataOut_payload_0_15199 ? _zz_dataOut_payload_0_15025 : _zz_dataOut_payload_0_15049);
  assign _zz_dataOut_payload_0_15201 = (_zz_dataOut_payload_0_15199 ? _zz_dataOut_payload_0_15049 : _zz_dataOut_payload_0_15025);
  assign _zz_dataOut_payload_0_15202 = (_zz_dataOut_payload_0_15028 < _zz_dataOut_payload_0_15052);
  assign _zz_dataOut_payload_0_15203 = (_zz_dataOut_payload_0_15202 ? _zz_dataOut_payload_0_15028 : _zz_dataOut_payload_0_15052);
  assign _zz_dataOut_payload_0_15204 = (_zz_dataOut_payload_0_15202 ? _zz_dataOut_payload_0_15052 : _zz_dataOut_payload_0_15028);
  assign _zz_dataOut_payload_0_15205 = (_zz_dataOut_payload_0_15031 < _zz_dataOut_payload_0_15055);
  assign _zz_dataOut_payload_0_15206 = (_zz_dataOut_payload_0_15205 ? _zz_dataOut_payload_0_15031 : _zz_dataOut_payload_0_15055);
  assign _zz_dataOut_payload_0_15207 = (_zz_dataOut_payload_0_15205 ? _zz_dataOut_payload_0_15055 : _zz_dataOut_payload_0_15031);
  assign _zz_dataOut_payload_0_15208 = (_zz_dataOut_payload_0_15185 < _zz_dataOut_payload_0_15197);
  assign _zz_dataOut_payload_0_15209 = (_zz_dataOut_payload_0_15208 ? _zz_dataOut_payload_0_15185 : _zz_dataOut_payload_0_15197);
  assign _zz_dataOut_payload_0_15210 = (_zz_dataOut_payload_0_15208 ? _zz_dataOut_payload_0_15197 : _zz_dataOut_payload_0_15185);
  assign _zz_dataOut_payload_0_15211 = (_zz_dataOut_payload_0_15188 < _zz_dataOut_payload_0_15200);
  assign _zz_dataOut_payload_0_15212 = (_zz_dataOut_payload_0_15211 ? _zz_dataOut_payload_0_15188 : _zz_dataOut_payload_0_15200);
  assign _zz_dataOut_payload_0_15213 = (_zz_dataOut_payload_0_15211 ? _zz_dataOut_payload_0_15200 : _zz_dataOut_payload_0_15188);
  assign _zz_dataOut_payload_0_15214 = (_zz_dataOut_payload_0_15191 < _zz_dataOut_payload_0_15203);
  assign _zz_dataOut_payload_0_15215 = (_zz_dataOut_payload_0_15214 ? _zz_dataOut_payload_0_15191 : _zz_dataOut_payload_0_15203);
  assign _zz_dataOut_payload_0_15216 = (_zz_dataOut_payload_0_15214 ? _zz_dataOut_payload_0_15203 : _zz_dataOut_payload_0_15191);
  assign _zz_dataOut_payload_0_15217 = (_zz_dataOut_payload_0_15194 < _zz_dataOut_payload_0_15206);
  assign _zz_dataOut_payload_0_15218 = (_zz_dataOut_payload_0_15217 ? _zz_dataOut_payload_0_15194 : _zz_dataOut_payload_0_15206);
  assign _zz_dataOut_payload_0_15219 = (_zz_dataOut_payload_0_15217 ? _zz_dataOut_payload_0_15206 : _zz_dataOut_payload_0_15194);
  assign _zz_dataOut_payload_0_15220 = (_zz_dataOut_payload_0_15209 < _zz_dataOut_payload_0_15215);
  assign _zz_dataOut_payload_0_15221 = (_zz_dataOut_payload_0_15220 ? _zz_dataOut_payload_0_15209 : _zz_dataOut_payload_0_15215);
  assign _zz_dataOut_payload_0_15222 = (_zz_dataOut_payload_0_15220 ? _zz_dataOut_payload_0_15215 : _zz_dataOut_payload_0_15209);
  assign _zz_dataOut_payload_0_15223 = (_zz_dataOut_payload_0_15212 < _zz_dataOut_payload_0_15218);
  assign _zz_dataOut_payload_0_15224 = (_zz_dataOut_payload_0_15223 ? _zz_dataOut_payload_0_15212 : _zz_dataOut_payload_0_15218);
  assign _zz_dataOut_payload_0_15225 = (_zz_dataOut_payload_0_15223 ? _zz_dataOut_payload_0_15218 : _zz_dataOut_payload_0_15212);
  assign _zz_dataOut_payload_0_15226 = (_zz_dataOut_payload_0_15221 < _zz_dataOut_payload_0_15224);
  assign _zz_dataOut_payload_0_15227 = (_zz_dataOut_payload_0_15222 < _zz_dataOut_payload_0_15225);
  assign _zz_dataOut_payload_0_15232 = (_zz_dataOut_payload_0_15210 < _zz_dataOut_payload_0_15216);
  assign _zz_dataOut_payload_0_15233 = (_zz_dataOut_payload_0_15232 ? _zz_dataOut_payload_0_15210 : _zz_dataOut_payload_0_15216);
  assign _zz_dataOut_payload_0_15234 = (_zz_dataOut_payload_0_15232 ? _zz_dataOut_payload_0_15216 : _zz_dataOut_payload_0_15210);
  assign _zz_dataOut_payload_0_15235 = (_zz_dataOut_payload_0_15213 < _zz_dataOut_payload_0_15219);
  assign _zz_dataOut_payload_0_15236 = (_zz_dataOut_payload_0_15235 ? _zz_dataOut_payload_0_15213 : _zz_dataOut_payload_0_15219);
  assign _zz_dataOut_payload_0_15237 = (_zz_dataOut_payload_0_15235 ? _zz_dataOut_payload_0_15219 : _zz_dataOut_payload_0_15213);
  assign _zz_dataOut_payload_0_15238 = (_zz_dataOut_payload_0_15233 < _zz_dataOut_payload_0_15236);
  assign _zz_dataOut_payload_0_15239 = (_zz_dataOut_payload_0_15234 < _zz_dataOut_payload_0_15237);
  assign _zz_dataOut_payload_0_15252 = (_zz_dataOut_payload_0_15186 < _zz_dataOut_payload_0_15198);
  assign _zz_dataOut_payload_0_15253 = (_zz_dataOut_payload_0_15252 ? _zz_dataOut_payload_0_15186 : _zz_dataOut_payload_0_15198);
  assign _zz_dataOut_payload_0_15254 = (_zz_dataOut_payload_0_15252 ? _zz_dataOut_payload_0_15198 : _zz_dataOut_payload_0_15186);
  assign _zz_dataOut_payload_0_15255 = (_zz_dataOut_payload_0_15189 < _zz_dataOut_payload_0_15201);
  assign _zz_dataOut_payload_0_15256 = (_zz_dataOut_payload_0_15255 ? _zz_dataOut_payload_0_15189 : _zz_dataOut_payload_0_15201);
  assign _zz_dataOut_payload_0_15257 = (_zz_dataOut_payload_0_15255 ? _zz_dataOut_payload_0_15201 : _zz_dataOut_payload_0_15189);
  assign _zz_dataOut_payload_0_15258 = (_zz_dataOut_payload_0_15192 < _zz_dataOut_payload_0_15204);
  assign _zz_dataOut_payload_0_15259 = (_zz_dataOut_payload_0_15258 ? _zz_dataOut_payload_0_15192 : _zz_dataOut_payload_0_15204);
  assign _zz_dataOut_payload_0_15260 = (_zz_dataOut_payload_0_15258 ? _zz_dataOut_payload_0_15204 : _zz_dataOut_payload_0_15192);
  assign _zz_dataOut_payload_0_15261 = (_zz_dataOut_payload_0_15195 < _zz_dataOut_payload_0_15207);
  assign _zz_dataOut_payload_0_15262 = (_zz_dataOut_payload_0_15261 ? _zz_dataOut_payload_0_15195 : _zz_dataOut_payload_0_15207);
  assign _zz_dataOut_payload_0_15263 = (_zz_dataOut_payload_0_15261 ? _zz_dataOut_payload_0_15207 : _zz_dataOut_payload_0_15195);
  assign _zz_dataOut_payload_0_15264 = (_zz_dataOut_payload_0_15253 < _zz_dataOut_payload_0_15259);
  assign _zz_dataOut_payload_0_15265 = (_zz_dataOut_payload_0_15264 ? _zz_dataOut_payload_0_15253 : _zz_dataOut_payload_0_15259);
  assign _zz_dataOut_payload_0_15266 = (_zz_dataOut_payload_0_15264 ? _zz_dataOut_payload_0_15259 : _zz_dataOut_payload_0_15253);
  assign _zz_dataOut_payload_0_15267 = (_zz_dataOut_payload_0_15256 < _zz_dataOut_payload_0_15262);
  assign _zz_dataOut_payload_0_15268 = (_zz_dataOut_payload_0_15267 ? _zz_dataOut_payload_0_15256 : _zz_dataOut_payload_0_15262);
  assign _zz_dataOut_payload_0_15269 = (_zz_dataOut_payload_0_15267 ? _zz_dataOut_payload_0_15262 : _zz_dataOut_payload_0_15256);
  assign _zz_dataOut_payload_0_15270 = (_zz_dataOut_payload_0_15265 < _zz_dataOut_payload_0_15268);
  assign _zz_dataOut_payload_0_15271 = (_zz_dataOut_payload_0_15266 < _zz_dataOut_payload_0_15269);
  assign _zz_dataOut_payload_0_15276 = (_zz_dataOut_payload_0_15254 < _zz_dataOut_payload_0_15260);
  assign _zz_dataOut_payload_0_15277 = (_zz_dataOut_payload_0_15276 ? _zz_dataOut_payload_0_15254 : _zz_dataOut_payload_0_15260);
  assign _zz_dataOut_payload_0_15278 = (_zz_dataOut_payload_0_15276 ? _zz_dataOut_payload_0_15260 : _zz_dataOut_payload_0_15254);
  assign _zz_dataOut_payload_0_15279 = (_zz_dataOut_payload_0_15257 < _zz_dataOut_payload_0_15263);
  assign _zz_dataOut_payload_0_15280 = (_zz_dataOut_payload_0_15279 ? _zz_dataOut_payload_0_15257 : _zz_dataOut_payload_0_15263);
  assign _zz_dataOut_payload_0_15281 = (_zz_dataOut_payload_0_15279 ? _zz_dataOut_payload_0_15263 : _zz_dataOut_payload_0_15257);
  assign _zz_dataOut_payload_0_15282 = (_zz_dataOut_payload_0_15277 < _zz_dataOut_payload_0_15280);
  assign _zz_dataOut_payload_0_15283 = (_zz_dataOut_payload_0_15278 < _zz_dataOut_payload_0_15281);
  assign _zz_dataOut_payload_0_15344 = (_zz_dataOut_payload_0_14914 < _zz_dataOut_payload_0_14962);
  assign _zz_dataOut_payload_0_15345 = (_zz_dataOut_payload_0_15344 ? _zz_dataOut_payload_0_14914 : _zz_dataOut_payload_0_14962);
  assign _zz_dataOut_payload_0_15346 = (_zz_dataOut_payload_0_15344 ? _zz_dataOut_payload_0_14962 : _zz_dataOut_payload_0_14914);
  assign _zz_dataOut_payload_0_15347 = (_zz_dataOut_payload_0_14917 < _zz_dataOut_payload_0_14965);
  assign _zz_dataOut_payload_0_15348 = (_zz_dataOut_payload_0_15347 ? _zz_dataOut_payload_0_14917 : _zz_dataOut_payload_0_14965);
  assign _zz_dataOut_payload_0_15349 = (_zz_dataOut_payload_0_15347 ? _zz_dataOut_payload_0_14965 : _zz_dataOut_payload_0_14917);
  assign _zz_dataOut_payload_0_15350 = (_zz_dataOut_payload_0_14920 < _zz_dataOut_payload_0_14968);
  assign _zz_dataOut_payload_0_15351 = (_zz_dataOut_payload_0_15350 ? _zz_dataOut_payload_0_14920 : _zz_dataOut_payload_0_14968);
  assign _zz_dataOut_payload_0_15352 = (_zz_dataOut_payload_0_15350 ? _zz_dataOut_payload_0_14968 : _zz_dataOut_payload_0_14920);
  assign _zz_dataOut_payload_0_15353 = (_zz_dataOut_payload_0_14923 < _zz_dataOut_payload_0_14971);
  assign _zz_dataOut_payload_0_15354 = (_zz_dataOut_payload_0_15353 ? _zz_dataOut_payload_0_14923 : _zz_dataOut_payload_0_14971);
  assign _zz_dataOut_payload_0_15355 = (_zz_dataOut_payload_0_15353 ? _zz_dataOut_payload_0_14971 : _zz_dataOut_payload_0_14923);
  assign _zz_dataOut_payload_0_15356 = (_zz_dataOut_payload_0_14926 < _zz_dataOut_payload_0_14974);
  assign _zz_dataOut_payload_0_15357 = (_zz_dataOut_payload_0_15356 ? _zz_dataOut_payload_0_14926 : _zz_dataOut_payload_0_14974);
  assign _zz_dataOut_payload_0_15358 = (_zz_dataOut_payload_0_15356 ? _zz_dataOut_payload_0_14974 : _zz_dataOut_payload_0_14926);
  assign _zz_dataOut_payload_0_15359 = (_zz_dataOut_payload_0_14929 < _zz_dataOut_payload_0_14977);
  assign _zz_dataOut_payload_0_15360 = (_zz_dataOut_payload_0_15359 ? _zz_dataOut_payload_0_14929 : _zz_dataOut_payload_0_14977);
  assign _zz_dataOut_payload_0_15361 = (_zz_dataOut_payload_0_15359 ? _zz_dataOut_payload_0_14977 : _zz_dataOut_payload_0_14929);
  assign _zz_dataOut_payload_0_15362 = (_zz_dataOut_payload_0_14932 < _zz_dataOut_payload_0_14980);
  assign _zz_dataOut_payload_0_15363 = (_zz_dataOut_payload_0_15362 ? _zz_dataOut_payload_0_14932 : _zz_dataOut_payload_0_14980);
  assign _zz_dataOut_payload_0_15364 = (_zz_dataOut_payload_0_15362 ? _zz_dataOut_payload_0_14980 : _zz_dataOut_payload_0_14932);
  assign _zz_dataOut_payload_0_15365 = (_zz_dataOut_payload_0_14935 < _zz_dataOut_payload_0_14983);
  assign _zz_dataOut_payload_0_15366 = (_zz_dataOut_payload_0_15365 ? _zz_dataOut_payload_0_14935 : _zz_dataOut_payload_0_14983);
  assign _zz_dataOut_payload_0_15367 = (_zz_dataOut_payload_0_15365 ? _zz_dataOut_payload_0_14983 : _zz_dataOut_payload_0_14935);
  assign _zz_dataOut_payload_0_15368 = (_zz_dataOut_payload_0_14938 < _zz_dataOut_payload_0_14986);
  assign _zz_dataOut_payload_0_15369 = (_zz_dataOut_payload_0_15368 ? _zz_dataOut_payload_0_14938 : _zz_dataOut_payload_0_14986);
  assign _zz_dataOut_payload_0_15370 = (_zz_dataOut_payload_0_15368 ? _zz_dataOut_payload_0_14986 : _zz_dataOut_payload_0_14938);
  assign _zz_dataOut_payload_0_15371 = (_zz_dataOut_payload_0_14941 < _zz_dataOut_payload_0_14989);
  assign _zz_dataOut_payload_0_15372 = (_zz_dataOut_payload_0_15371 ? _zz_dataOut_payload_0_14941 : _zz_dataOut_payload_0_14989);
  assign _zz_dataOut_payload_0_15373 = (_zz_dataOut_payload_0_15371 ? _zz_dataOut_payload_0_14989 : _zz_dataOut_payload_0_14941);
  assign _zz_dataOut_payload_0_15374 = (_zz_dataOut_payload_0_14944 < _zz_dataOut_payload_0_14992);
  assign _zz_dataOut_payload_0_15375 = (_zz_dataOut_payload_0_15374 ? _zz_dataOut_payload_0_14944 : _zz_dataOut_payload_0_14992);
  assign _zz_dataOut_payload_0_15376 = (_zz_dataOut_payload_0_15374 ? _zz_dataOut_payload_0_14992 : _zz_dataOut_payload_0_14944);
  assign _zz_dataOut_payload_0_15377 = (_zz_dataOut_payload_0_14947 < _zz_dataOut_payload_0_14995);
  assign _zz_dataOut_payload_0_15378 = (_zz_dataOut_payload_0_15377 ? _zz_dataOut_payload_0_14947 : _zz_dataOut_payload_0_14995);
  assign _zz_dataOut_payload_0_15379 = (_zz_dataOut_payload_0_15377 ? _zz_dataOut_payload_0_14995 : _zz_dataOut_payload_0_14947);
  assign _zz_dataOut_payload_0_15380 = (_zz_dataOut_payload_0_14950 < _zz_dataOut_payload_0_14998);
  assign _zz_dataOut_payload_0_15381 = (_zz_dataOut_payload_0_15380 ? _zz_dataOut_payload_0_14950 : _zz_dataOut_payload_0_14998);
  assign _zz_dataOut_payload_0_15382 = (_zz_dataOut_payload_0_15380 ? _zz_dataOut_payload_0_14998 : _zz_dataOut_payload_0_14950);
  assign _zz_dataOut_payload_0_15383 = (_zz_dataOut_payload_0_14953 < _zz_dataOut_payload_0_15001);
  assign _zz_dataOut_payload_0_15384 = (_zz_dataOut_payload_0_15383 ? _zz_dataOut_payload_0_14953 : _zz_dataOut_payload_0_15001);
  assign _zz_dataOut_payload_0_15385 = (_zz_dataOut_payload_0_15383 ? _zz_dataOut_payload_0_15001 : _zz_dataOut_payload_0_14953);
  assign _zz_dataOut_payload_0_15386 = (_zz_dataOut_payload_0_14956 < _zz_dataOut_payload_0_15004);
  assign _zz_dataOut_payload_0_15387 = (_zz_dataOut_payload_0_15386 ? _zz_dataOut_payload_0_14956 : _zz_dataOut_payload_0_15004);
  assign _zz_dataOut_payload_0_15388 = (_zz_dataOut_payload_0_15386 ? _zz_dataOut_payload_0_15004 : _zz_dataOut_payload_0_14956);
  assign _zz_dataOut_payload_0_15389 = (_zz_dataOut_payload_0_14959 < _zz_dataOut_payload_0_15007);
  assign _zz_dataOut_payload_0_15390 = (_zz_dataOut_payload_0_15389 ? _zz_dataOut_payload_0_14959 : _zz_dataOut_payload_0_15007);
  assign _zz_dataOut_payload_0_15391 = (_zz_dataOut_payload_0_15389 ? _zz_dataOut_payload_0_15007 : _zz_dataOut_payload_0_14959);
  assign _zz_dataOut_payload_0_15392 = (_zz_dataOut_payload_0_15345 < _zz_dataOut_payload_0_15369);
  assign _zz_dataOut_payload_0_15393 = (_zz_dataOut_payload_0_15392 ? _zz_dataOut_payload_0_15345 : _zz_dataOut_payload_0_15369);
  assign _zz_dataOut_payload_0_15394 = (_zz_dataOut_payload_0_15392 ? _zz_dataOut_payload_0_15369 : _zz_dataOut_payload_0_15345);
  assign _zz_dataOut_payload_0_15395 = (_zz_dataOut_payload_0_15348 < _zz_dataOut_payload_0_15372);
  assign _zz_dataOut_payload_0_15396 = (_zz_dataOut_payload_0_15395 ? _zz_dataOut_payload_0_15348 : _zz_dataOut_payload_0_15372);
  assign _zz_dataOut_payload_0_15397 = (_zz_dataOut_payload_0_15395 ? _zz_dataOut_payload_0_15372 : _zz_dataOut_payload_0_15348);
  assign _zz_dataOut_payload_0_15398 = (_zz_dataOut_payload_0_15351 < _zz_dataOut_payload_0_15375);
  assign _zz_dataOut_payload_0_15399 = (_zz_dataOut_payload_0_15398 ? _zz_dataOut_payload_0_15351 : _zz_dataOut_payload_0_15375);
  assign _zz_dataOut_payload_0_15400 = (_zz_dataOut_payload_0_15398 ? _zz_dataOut_payload_0_15375 : _zz_dataOut_payload_0_15351);
  assign _zz_dataOut_payload_0_15401 = (_zz_dataOut_payload_0_15354 < _zz_dataOut_payload_0_15378);
  assign _zz_dataOut_payload_0_15402 = (_zz_dataOut_payload_0_15401 ? _zz_dataOut_payload_0_15354 : _zz_dataOut_payload_0_15378);
  assign _zz_dataOut_payload_0_15403 = (_zz_dataOut_payload_0_15401 ? _zz_dataOut_payload_0_15378 : _zz_dataOut_payload_0_15354);
  assign _zz_dataOut_payload_0_15404 = (_zz_dataOut_payload_0_15357 < _zz_dataOut_payload_0_15381);
  assign _zz_dataOut_payload_0_15405 = (_zz_dataOut_payload_0_15404 ? _zz_dataOut_payload_0_15357 : _zz_dataOut_payload_0_15381);
  assign _zz_dataOut_payload_0_15406 = (_zz_dataOut_payload_0_15404 ? _zz_dataOut_payload_0_15381 : _zz_dataOut_payload_0_15357);
  assign _zz_dataOut_payload_0_15407 = (_zz_dataOut_payload_0_15360 < _zz_dataOut_payload_0_15384);
  assign _zz_dataOut_payload_0_15408 = (_zz_dataOut_payload_0_15407 ? _zz_dataOut_payload_0_15360 : _zz_dataOut_payload_0_15384);
  assign _zz_dataOut_payload_0_15409 = (_zz_dataOut_payload_0_15407 ? _zz_dataOut_payload_0_15384 : _zz_dataOut_payload_0_15360);
  assign _zz_dataOut_payload_0_15410 = (_zz_dataOut_payload_0_15363 < _zz_dataOut_payload_0_15387);
  assign _zz_dataOut_payload_0_15411 = (_zz_dataOut_payload_0_15410 ? _zz_dataOut_payload_0_15363 : _zz_dataOut_payload_0_15387);
  assign _zz_dataOut_payload_0_15412 = (_zz_dataOut_payload_0_15410 ? _zz_dataOut_payload_0_15387 : _zz_dataOut_payload_0_15363);
  assign _zz_dataOut_payload_0_15413 = (_zz_dataOut_payload_0_15366 < _zz_dataOut_payload_0_15390);
  assign _zz_dataOut_payload_0_15414 = (_zz_dataOut_payload_0_15413 ? _zz_dataOut_payload_0_15366 : _zz_dataOut_payload_0_15390);
  assign _zz_dataOut_payload_0_15415 = (_zz_dataOut_payload_0_15413 ? _zz_dataOut_payload_0_15390 : _zz_dataOut_payload_0_15366);
  assign _zz_dataOut_payload_0_15416 = (_zz_dataOut_payload_0_15393 < _zz_dataOut_payload_0_15405);
  assign _zz_dataOut_payload_0_15417 = (_zz_dataOut_payload_0_15416 ? _zz_dataOut_payload_0_15393 : _zz_dataOut_payload_0_15405);
  assign _zz_dataOut_payload_0_15418 = (_zz_dataOut_payload_0_15416 ? _zz_dataOut_payload_0_15405 : _zz_dataOut_payload_0_15393);
  assign _zz_dataOut_payload_0_15419 = (_zz_dataOut_payload_0_15396 < _zz_dataOut_payload_0_15408);
  assign _zz_dataOut_payload_0_15420 = (_zz_dataOut_payload_0_15419 ? _zz_dataOut_payload_0_15396 : _zz_dataOut_payload_0_15408);
  assign _zz_dataOut_payload_0_15421 = (_zz_dataOut_payload_0_15419 ? _zz_dataOut_payload_0_15408 : _zz_dataOut_payload_0_15396);
  assign _zz_dataOut_payload_0_15422 = (_zz_dataOut_payload_0_15399 < _zz_dataOut_payload_0_15411);
  assign _zz_dataOut_payload_0_15423 = (_zz_dataOut_payload_0_15422 ? _zz_dataOut_payload_0_15399 : _zz_dataOut_payload_0_15411);
  assign _zz_dataOut_payload_0_15424 = (_zz_dataOut_payload_0_15422 ? _zz_dataOut_payload_0_15411 : _zz_dataOut_payload_0_15399);
  assign _zz_dataOut_payload_0_15425 = (_zz_dataOut_payload_0_15402 < _zz_dataOut_payload_0_15414);
  assign _zz_dataOut_payload_0_15426 = (_zz_dataOut_payload_0_15425 ? _zz_dataOut_payload_0_15402 : _zz_dataOut_payload_0_15414);
  assign _zz_dataOut_payload_0_15427 = (_zz_dataOut_payload_0_15425 ? _zz_dataOut_payload_0_15414 : _zz_dataOut_payload_0_15402);
  assign _zz_dataOut_payload_0_15428 = (_zz_dataOut_payload_0_15417 < _zz_dataOut_payload_0_15423);
  assign _zz_dataOut_payload_0_15429 = (_zz_dataOut_payload_0_15428 ? _zz_dataOut_payload_0_15417 : _zz_dataOut_payload_0_15423);
  assign _zz_dataOut_payload_0_15430 = (_zz_dataOut_payload_0_15428 ? _zz_dataOut_payload_0_15423 : _zz_dataOut_payload_0_15417);
  assign _zz_dataOut_payload_0_15431 = (_zz_dataOut_payload_0_15420 < _zz_dataOut_payload_0_15426);
  assign _zz_dataOut_payload_0_15432 = (_zz_dataOut_payload_0_15431 ? _zz_dataOut_payload_0_15420 : _zz_dataOut_payload_0_15426);
  assign _zz_dataOut_payload_0_15433 = (_zz_dataOut_payload_0_15431 ? _zz_dataOut_payload_0_15426 : _zz_dataOut_payload_0_15420);
  assign _zz_dataOut_payload_0_15434 = (_zz_dataOut_payload_0_15429 < _zz_dataOut_payload_0_15432);
  assign _zz_dataOut_payload_0_15435 = (_zz_dataOut_payload_0_15430 < _zz_dataOut_payload_0_15433);
  assign _zz_dataOut_payload_0_15440 = (_zz_dataOut_payload_0_15418 < _zz_dataOut_payload_0_15424);
  assign _zz_dataOut_payload_0_15441 = (_zz_dataOut_payload_0_15440 ? _zz_dataOut_payload_0_15418 : _zz_dataOut_payload_0_15424);
  assign _zz_dataOut_payload_0_15442 = (_zz_dataOut_payload_0_15440 ? _zz_dataOut_payload_0_15424 : _zz_dataOut_payload_0_15418);
  assign _zz_dataOut_payload_0_15443 = (_zz_dataOut_payload_0_15421 < _zz_dataOut_payload_0_15427);
  assign _zz_dataOut_payload_0_15444 = (_zz_dataOut_payload_0_15443 ? _zz_dataOut_payload_0_15421 : _zz_dataOut_payload_0_15427);
  assign _zz_dataOut_payload_0_15445 = (_zz_dataOut_payload_0_15443 ? _zz_dataOut_payload_0_15427 : _zz_dataOut_payload_0_15421);
  assign _zz_dataOut_payload_0_15446 = (_zz_dataOut_payload_0_15441 < _zz_dataOut_payload_0_15444);
  assign _zz_dataOut_payload_0_15447 = (_zz_dataOut_payload_0_15442 < _zz_dataOut_payload_0_15445);
  assign _zz_dataOut_payload_0_15460 = (_zz_dataOut_payload_0_15394 < _zz_dataOut_payload_0_15406);
  assign _zz_dataOut_payload_0_15461 = (_zz_dataOut_payload_0_15460 ? _zz_dataOut_payload_0_15394 : _zz_dataOut_payload_0_15406);
  assign _zz_dataOut_payload_0_15462 = (_zz_dataOut_payload_0_15460 ? _zz_dataOut_payload_0_15406 : _zz_dataOut_payload_0_15394);
  assign _zz_dataOut_payload_0_15463 = (_zz_dataOut_payload_0_15397 < _zz_dataOut_payload_0_15409);
  assign _zz_dataOut_payload_0_15464 = (_zz_dataOut_payload_0_15463 ? _zz_dataOut_payload_0_15397 : _zz_dataOut_payload_0_15409);
  assign _zz_dataOut_payload_0_15465 = (_zz_dataOut_payload_0_15463 ? _zz_dataOut_payload_0_15409 : _zz_dataOut_payload_0_15397);
  assign _zz_dataOut_payload_0_15466 = (_zz_dataOut_payload_0_15400 < _zz_dataOut_payload_0_15412);
  assign _zz_dataOut_payload_0_15467 = (_zz_dataOut_payload_0_15466 ? _zz_dataOut_payload_0_15400 : _zz_dataOut_payload_0_15412);
  assign _zz_dataOut_payload_0_15468 = (_zz_dataOut_payload_0_15466 ? _zz_dataOut_payload_0_15412 : _zz_dataOut_payload_0_15400);
  assign _zz_dataOut_payload_0_15469 = (_zz_dataOut_payload_0_15403 < _zz_dataOut_payload_0_15415);
  assign _zz_dataOut_payload_0_15470 = (_zz_dataOut_payload_0_15469 ? _zz_dataOut_payload_0_15403 : _zz_dataOut_payload_0_15415);
  assign _zz_dataOut_payload_0_15471 = (_zz_dataOut_payload_0_15469 ? _zz_dataOut_payload_0_15415 : _zz_dataOut_payload_0_15403);
  assign _zz_dataOut_payload_0_15472 = (_zz_dataOut_payload_0_15461 < _zz_dataOut_payload_0_15467);
  assign _zz_dataOut_payload_0_15473 = (_zz_dataOut_payload_0_15472 ? _zz_dataOut_payload_0_15461 : _zz_dataOut_payload_0_15467);
  assign _zz_dataOut_payload_0_15474 = (_zz_dataOut_payload_0_15472 ? _zz_dataOut_payload_0_15467 : _zz_dataOut_payload_0_15461);
  assign _zz_dataOut_payload_0_15475 = (_zz_dataOut_payload_0_15464 < _zz_dataOut_payload_0_15470);
  assign _zz_dataOut_payload_0_15476 = (_zz_dataOut_payload_0_15475 ? _zz_dataOut_payload_0_15464 : _zz_dataOut_payload_0_15470);
  assign _zz_dataOut_payload_0_15477 = (_zz_dataOut_payload_0_15475 ? _zz_dataOut_payload_0_15470 : _zz_dataOut_payload_0_15464);
  assign _zz_dataOut_payload_0_15478 = (_zz_dataOut_payload_0_15473 < _zz_dataOut_payload_0_15476);
  assign _zz_dataOut_payload_0_15479 = (_zz_dataOut_payload_0_15474 < _zz_dataOut_payload_0_15477);
  assign _zz_dataOut_payload_0_15484 = (_zz_dataOut_payload_0_15462 < _zz_dataOut_payload_0_15468);
  assign _zz_dataOut_payload_0_15485 = (_zz_dataOut_payload_0_15484 ? _zz_dataOut_payload_0_15462 : _zz_dataOut_payload_0_15468);
  assign _zz_dataOut_payload_0_15486 = (_zz_dataOut_payload_0_15484 ? _zz_dataOut_payload_0_15468 : _zz_dataOut_payload_0_15462);
  assign _zz_dataOut_payload_0_15487 = (_zz_dataOut_payload_0_15465 < _zz_dataOut_payload_0_15471);
  assign _zz_dataOut_payload_0_15488 = (_zz_dataOut_payload_0_15487 ? _zz_dataOut_payload_0_15465 : _zz_dataOut_payload_0_15471);
  assign _zz_dataOut_payload_0_15489 = (_zz_dataOut_payload_0_15487 ? _zz_dataOut_payload_0_15471 : _zz_dataOut_payload_0_15465);
  assign _zz_dataOut_payload_0_15490 = (_zz_dataOut_payload_0_15485 < _zz_dataOut_payload_0_15488);
  assign _zz_dataOut_payload_0_15491 = (_zz_dataOut_payload_0_15486 < _zz_dataOut_payload_0_15489);
  assign _zz_dataOut_payload_0_15520 = (_zz_dataOut_payload_0_15346 < _zz_dataOut_payload_0_15370);
  assign _zz_dataOut_payload_0_15521 = (_zz_dataOut_payload_0_15520 ? _zz_dataOut_payload_0_15346 : _zz_dataOut_payload_0_15370);
  assign _zz_dataOut_payload_0_15522 = (_zz_dataOut_payload_0_15520 ? _zz_dataOut_payload_0_15370 : _zz_dataOut_payload_0_15346);
  assign _zz_dataOut_payload_0_15523 = (_zz_dataOut_payload_0_15349 < _zz_dataOut_payload_0_15373);
  assign _zz_dataOut_payload_0_15524 = (_zz_dataOut_payload_0_15523 ? _zz_dataOut_payload_0_15349 : _zz_dataOut_payload_0_15373);
  assign _zz_dataOut_payload_0_15525 = (_zz_dataOut_payload_0_15523 ? _zz_dataOut_payload_0_15373 : _zz_dataOut_payload_0_15349);
  assign _zz_dataOut_payload_0_15526 = (_zz_dataOut_payload_0_15352 < _zz_dataOut_payload_0_15376);
  assign _zz_dataOut_payload_0_15527 = (_zz_dataOut_payload_0_15526 ? _zz_dataOut_payload_0_15352 : _zz_dataOut_payload_0_15376);
  assign _zz_dataOut_payload_0_15528 = (_zz_dataOut_payload_0_15526 ? _zz_dataOut_payload_0_15376 : _zz_dataOut_payload_0_15352);
  assign _zz_dataOut_payload_0_15529 = (_zz_dataOut_payload_0_15355 < _zz_dataOut_payload_0_15379);
  assign _zz_dataOut_payload_0_15530 = (_zz_dataOut_payload_0_15529 ? _zz_dataOut_payload_0_15355 : _zz_dataOut_payload_0_15379);
  assign _zz_dataOut_payload_0_15531 = (_zz_dataOut_payload_0_15529 ? _zz_dataOut_payload_0_15379 : _zz_dataOut_payload_0_15355);
  assign _zz_dataOut_payload_0_15532 = (_zz_dataOut_payload_0_15358 < _zz_dataOut_payload_0_15382);
  assign _zz_dataOut_payload_0_15533 = (_zz_dataOut_payload_0_15532 ? _zz_dataOut_payload_0_15358 : _zz_dataOut_payload_0_15382);
  assign _zz_dataOut_payload_0_15534 = (_zz_dataOut_payload_0_15532 ? _zz_dataOut_payload_0_15382 : _zz_dataOut_payload_0_15358);
  assign _zz_dataOut_payload_0_15535 = (_zz_dataOut_payload_0_15361 < _zz_dataOut_payload_0_15385);
  assign _zz_dataOut_payload_0_15536 = (_zz_dataOut_payload_0_15535 ? _zz_dataOut_payload_0_15361 : _zz_dataOut_payload_0_15385);
  assign _zz_dataOut_payload_0_15537 = (_zz_dataOut_payload_0_15535 ? _zz_dataOut_payload_0_15385 : _zz_dataOut_payload_0_15361);
  assign _zz_dataOut_payload_0_15538 = (_zz_dataOut_payload_0_15364 < _zz_dataOut_payload_0_15388);
  assign _zz_dataOut_payload_0_15539 = (_zz_dataOut_payload_0_15538 ? _zz_dataOut_payload_0_15364 : _zz_dataOut_payload_0_15388);
  assign _zz_dataOut_payload_0_15540 = (_zz_dataOut_payload_0_15538 ? _zz_dataOut_payload_0_15388 : _zz_dataOut_payload_0_15364);
  assign _zz_dataOut_payload_0_15541 = (_zz_dataOut_payload_0_15367 < _zz_dataOut_payload_0_15391);
  assign _zz_dataOut_payload_0_15542 = (_zz_dataOut_payload_0_15541 ? _zz_dataOut_payload_0_15367 : _zz_dataOut_payload_0_15391);
  assign _zz_dataOut_payload_0_15543 = (_zz_dataOut_payload_0_15541 ? _zz_dataOut_payload_0_15391 : _zz_dataOut_payload_0_15367);
  assign _zz_dataOut_payload_0_15544 = (_zz_dataOut_payload_0_15521 < _zz_dataOut_payload_0_15533);
  assign _zz_dataOut_payload_0_15545 = (_zz_dataOut_payload_0_15544 ? _zz_dataOut_payload_0_15521 : _zz_dataOut_payload_0_15533);
  assign _zz_dataOut_payload_0_15546 = (_zz_dataOut_payload_0_15544 ? _zz_dataOut_payload_0_15533 : _zz_dataOut_payload_0_15521);
  assign _zz_dataOut_payload_0_15547 = (_zz_dataOut_payload_0_15524 < _zz_dataOut_payload_0_15536);
  assign _zz_dataOut_payload_0_15548 = (_zz_dataOut_payload_0_15547 ? _zz_dataOut_payload_0_15524 : _zz_dataOut_payload_0_15536);
  assign _zz_dataOut_payload_0_15549 = (_zz_dataOut_payload_0_15547 ? _zz_dataOut_payload_0_15536 : _zz_dataOut_payload_0_15524);
  assign _zz_dataOut_payload_0_15550 = (_zz_dataOut_payload_0_15527 < _zz_dataOut_payload_0_15539);
  assign _zz_dataOut_payload_0_15551 = (_zz_dataOut_payload_0_15550 ? _zz_dataOut_payload_0_15527 : _zz_dataOut_payload_0_15539);
  assign _zz_dataOut_payload_0_15552 = (_zz_dataOut_payload_0_15550 ? _zz_dataOut_payload_0_15539 : _zz_dataOut_payload_0_15527);
  assign _zz_dataOut_payload_0_15553 = (_zz_dataOut_payload_0_15530 < _zz_dataOut_payload_0_15542);
  assign _zz_dataOut_payload_0_15554 = (_zz_dataOut_payload_0_15553 ? _zz_dataOut_payload_0_15530 : _zz_dataOut_payload_0_15542);
  assign _zz_dataOut_payload_0_15555 = (_zz_dataOut_payload_0_15553 ? _zz_dataOut_payload_0_15542 : _zz_dataOut_payload_0_15530);
  assign _zz_dataOut_payload_0_15556 = (_zz_dataOut_payload_0_15545 < _zz_dataOut_payload_0_15551);
  assign _zz_dataOut_payload_0_15557 = (_zz_dataOut_payload_0_15556 ? _zz_dataOut_payload_0_15545 : _zz_dataOut_payload_0_15551);
  assign _zz_dataOut_payload_0_15558 = (_zz_dataOut_payload_0_15556 ? _zz_dataOut_payload_0_15551 : _zz_dataOut_payload_0_15545);
  assign _zz_dataOut_payload_0_15559 = (_zz_dataOut_payload_0_15548 < _zz_dataOut_payload_0_15554);
  assign _zz_dataOut_payload_0_15560 = (_zz_dataOut_payload_0_15559 ? _zz_dataOut_payload_0_15548 : _zz_dataOut_payload_0_15554);
  assign _zz_dataOut_payload_0_15561 = (_zz_dataOut_payload_0_15559 ? _zz_dataOut_payload_0_15554 : _zz_dataOut_payload_0_15548);
  assign _zz_dataOut_payload_0_15562 = (_zz_dataOut_payload_0_15557 < _zz_dataOut_payload_0_15560);
  assign _zz_dataOut_payload_0_15563 = (_zz_dataOut_payload_0_15558 < _zz_dataOut_payload_0_15561);
  assign _zz_dataOut_payload_0_15568 = (_zz_dataOut_payload_0_15546 < _zz_dataOut_payload_0_15552);
  assign _zz_dataOut_payload_0_15569 = (_zz_dataOut_payload_0_15568 ? _zz_dataOut_payload_0_15546 : _zz_dataOut_payload_0_15552);
  assign _zz_dataOut_payload_0_15570 = (_zz_dataOut_payload_0_15568 ? _zz_dataOut_payload_0_15552 : _zz_dataOut_payload_0_15546);
  assign _zz_dataOut_payload_0_15571 = (_zz_dataOut_payload_0_15549 < _zz_dataOut_payload_0_15555);
  assign _zz_dataOut_payload_0_15572 = (_zz_dataOut_payload_0_15571 ? _zz_dataOut_payload_0_15549 : _zz_dataOut_payload_0_15555);
  assign _zz_dataOut_payload_0_15573 = (_zz_dataOut_payload_0_15571 ? _zz_dataOut_payload_0_15555 : _zz_dataOut_payload_0_15549);
  assign _zz_dataOut_payload_0_15574 = (_zz_dataOut_payload_0_15569 < _zz_dataOut_payload_0_15572);
  assign _zz_dataOut_payload_0_15575 = (_zz_dataOut_payload_0_15570 < _zz_dataOut_payload_0_15573);
  assign _zz_dataOut_payload_0_15588 = (_zz_dataOut_payload_0_15522 < _zz_dataOut_payload_0_15534);
  assign _zz_dataOut_payload_0_15589 = (_zz_dataOut_payload_0_15588 ? _zz_dataOut_payload_0_15522 : _zz_dataOut_payload_0_15534);
  assign _zz_dataOut_payload_0_15590 = (_zz_dataOut_payload_0_15588 ? _zz_dataOut_payload_0_15534 : _zz_dataOut_payload_0_15522);
  assign _zz_dataOut_payload_0_15591 = (_zz_dataOut_payload_0_15525 < _zz_dataOut_payload_0_15537);
  assign _zz_dataOut_payload_0_15592 = (_zz_dataOut_payload_0_15591 ? _zz_dataOut_payload_0_15525 : _zz_dataOut_payload_0_15537);
  assign _zz_dataOut_payload_0_15593 = (_zz_dataOut_payload_0_15591 ? _zz_dataOut_payload_0_15537 : _zz_dataOut_payload_0_15525);
  assign _zz_dataOut_payload_0_15594 = (_zz_dataOut_payload_0_15528 < _zz_dataOut_payload_0_15540);
  assign _zz_dataOut_payload_0_15595 = (_zz_dataOut_payload_0_15594 ? _zz_dataOut_payload_0_15528 : _zz_dataOut_payload_0_15540);
  assign _zz_dataOut_payload_0_15596 = (_zz_dataOut_payload_0_15594 ? _zz_dataOut_payload_0_15540 : _zz_dataOut_payload_0_15528);
  assign _zz_dataOut_payload_0_15597 = (_zz_dataOut_payload_0_15531 < _zz_dataOut_payload_0_15543);
  assign _zz_dataOut_payload_0_15598 = (_zz_dataOut_payload_0_15597 ? _zz_dataOut_payload_0_15531 : _zz_dataOut_payload_0_15543);
  assign _zz_dataOut_payload_0_15599 = (_zz_dataOut_payload_0_15597 ? _zz_dataOut_payload_0_15543 : _zz_dataOut_payload_0_15531);
  assign _zz_dataOut_payload_0_15600 = (_zz_dataOut_payload_0_15589 < _zz_dataOut_payload_0_15595);
  assign _zz_dataOut_payload_0_15601 = (_zz_dataOut_payload_0_15600 ? _zz_dataOut_payload_0_15589 : _zz_dataOut_payload_0_15595);
  assign _zz_dataOut_payload_0_15602 = (_zz_dataOut_payload_0_15600 ? _zz_dataOut_payload_0_15595 : _zz_dataOut_payload_0_15589);
  assign _zz_dataOut_payload_0_15603 = (_zz_dataOut_payload_0_15592 < _zz_dataOut_payload_0_15598);
  assign _zz_dataOut_payload_0_15604 = (_zz_dataOut_payload_0_15603 ? _zz_dataOut_payload_0_15592 : _zz_dataOut_payload_0_15598);
  assign _zz_dataOut_payload_0_15605 = (_zz_dataOut_payload_0_15603 ? _zz_dataOut_payload_0_15598 : _zz_dataOut_payload_0_15592);
  assign _zz_dataOut_payload_0_15606 = (_zz_dataOut_payload_0_15601 < _zz_dataOut_payload_0_15604);
  assign _zz_dataOut_payload_0_15607 = (_zz_dataOut_payload_0_15602 < _zz_dataOut_payload_0_15605);
  assign _zz_dataOut_payload_0_15612 = (_zz_dataOut_payload_0_15590 < _zz_dataOut_payload_0_15596);
  assign _zz_dataOut_payload_0_15613 = (_zz_dataOut_payload_0_15612 ? _zz_dataOut_payload_0_15590 : _zz_dataOut_payload_0_15596);
  assign _zz_dataOut_payload_0_15614 = (_zz_dataOut_payload_0_15612 ? _zz_dataOut_payload_0_15596 : _zz_dataOut_payload_0_15590);
  assign _zz_dataOut_payload_0_15615 = (_zz_dataOut_payload_0_15593 < _zz_dataOut_payload_0_15599);
  assign _zz_dataOut_payload_0_15616 = (_zz_dataOut_payload_0_15615 ? _zz_dataOut_payload_0_15593 : _zz_dataOut_payload_0_15599);
  assign _zz_dataOut_payload_0_15617 = (_zz_dataOut_payload_0_15615 ? _zz_dataOut_payload_0_15599 : _zz_dataOut_payload_0_15593);
  assign _zz_dataOut_payload_0_15618 = (_zz_dataOut_payload_0_15613 < _zz_dataOut_payload_0_15616);
  assign _zz_dataOut_payload_0_15619 = (_zz_dataOut_payload_0_15614 < _zz_dataOut_payload_0_15617);
  assign _zz_dataOut_payload_0_16128 = (_zz_dataOut_payload_0_15872 < _zz_dataOut_payload_0_16127);
  assign _zz_dataOut_payload_0_16129 = (_zz_dataOut_payload_0_16128 ? _zz_dataOut_payload_0_15872 : _zz_dataOut_payload_0_16127);
  assign _zz_dataOut_payload_128 = (_zz_dataOut_payload_0_16128 ? _zz_dataOut_payload_0_16127 : _zz_dataOut_payload_0_15872);
  assign _zz_dataOut_payload_0_16130 = (_zz_dataOut_payload_0_15873 < _zz_dataOut_payload_0_16126);
  assign _zz_dataOut_payload_0_16131 = (_zz_dataOut_payload_0_16130 ? _zz_dataOut_payload_0_15873 : _zz_dataOut_payload_0_16126);
  assign _zz_dataOut_payload_128_1 = (_zz_dataOut_payload_0_16130 ? _zz_dataOut_payload_0_16126 : _zz_dataOut_payload_0_15873);
  assign _zz_dataOut_payload_0_16132 = (_zz_dataOut_payload_0_15874 < _zz_dataOut_payload_0_16125);
  assign _zz_dataOut_payload_0_16133 = (_zz_dataOut_payload_0_16132 ? _zz_dataOut_payload_0_15874 : _zz_dataOut_payload_0_16125);
  assign _zz_dataOut_payload_128_2 = (_zz_dataOut_payload_0_16132 ? _zz_dataOut_payload_0_16125 : _zz_dataOut_payload_0_15874);
  assign _zz_dataOut_payload_0_16134 = (_zz_dataOut_payload_0_15875 < _zz_dataOut_payload_0_16124);
  assign _zz_dataOut_payload_0_16135 = (_zz_dataOut_payload_0_16134 ? _zz_dataOut_payload_0_15875 : _zz_dataOut_payload_0_16124);
  assign _zz_dataOut_payload_128_3 = (_zz_dataOut_payload_0_16134 ? _zz_dataOut_payload_0_16124 : _zz_dataOut_payload_0_15875);
  assign _zz_dataOut_payload_0_16136 = (_zz_dataOut_payload_0_15876 < _zz_dataOut_payload_0_16123);
  assign _zz_dataOut_payload_0_16137 = (_zz_dataOut_payload_0_16136 ? _zz_dataOut_payload_0_15876 : _zz_dataOut_payload_0_16123);
  assign _zz_dataOut_payload_128_4 = (_zz_dataOut_payload_0_16136 ? _zz_dataOut_payload_0_16123 : _zz_dataOut_payload_0_15876);
  assign _zz_dataOut_payload_0_16138 = (_zz_dataOut_payload_0_15877 < _zz_dataOut_payload_0_16122);
  assign _zz_dataOut_payload_0_16139 = (_zz_dataOut_payload_0_16138 ? _zz_dataOut_payload_0_15877 : _zz_dataOut_payload_0_16122);
  assign _zz_dataOut_payload_128_5 = (_zz_dataOut_payload_0_16138 ? _zz_dataOut_payload_0_16122 : _zz_dataOut_payload_0_15877);
  assign _zz_dataOut_payload_0_16140 = (_zz_dataOut_payload_0_15878 < _zz_dataOut_payload_0_16121);
  assign _zz_dataOut_payload_0_16141 = (_zz_dataOut_payload_0_16140 ? _zz_dataOut_payload_0_15878 : _zz_dataOut_payload_0_16121);
  assign _zz_dataOut_payload_128_6 = (_zz_dataOut_payload_0_16140 ? _zz_dataOut_payload_0_16121 : _zz_dataOut_payload_0_15878);
  assign _zz_dataOut_payload_0_16142 = (_zz_dataOut_payload_0_15879 < _zz_dataOut_payload_0_16120);
  assign _zz_dataOut_payload_0_16143 = (_zz_dataOut_payload_0_16142 ? _zz_dataOut_payload_0_15879 : _zz_dataOut_payload_0_16120);
  assign _zz_dataOut_payload_128_7 = (_zz_dataOut_payload_0_16142 ? _zz_dataOut_payload_0_16120 : _zz_dataOut_payload_0_15879);
  assign _zz_dataOut_payload_0_16144 = (_zz_dataOut_payload_0_15880 < _zz_dataOut_payload_0_16119);
  assign _zz_dataOut_payload_0_16145 = (_zz_dataOut_payload_0_16144 ? _zz_dataOut_payload_0_15880 : _zz_dataOut_payload_0_16119);
  assign _zz_dataOut_payload_128_8 = (_zz_dataOut_payload_0_16144 ? _zz_dataOut_payload_0_16119 : _zz_dataOut_payload_0_15880);
  assign _zz_dataOut_payload_0_16146 = (_zz_dataOut_payload_0_15881 < _zz_dataOut_payload_0_16118);
  assign _zz_dataOut_payload_0_16147 = (_zz_dataOut_payload_0_16146 ? _zz_dataOut_payload_0_15881 : _zz_dataOut_payload_0_16118);
  assign _zz_dataOut_payload_128_9 = (_zz_dataOut_payload_0_16146 ? _zz_dataOut_payload_0_16118 : _zz_dataOut_payload_0_15881);
  assign _zz_dataOut_payload_0_16148 = (_zz_dataOut_payload_0_15882 < _zz_dataOut_payload_0_16117);
  assign _zz_dataOut_payload_0_16149 = (_zz_dataOut_payload_0_16148 ? _zz_dataOut_payload_0_15882 : _zz_dataOut_payload_0_16117);
  assign _zz_dataOut_payload_128_10 = (_zz_dataOut_payload_0_16148 ? _zz_dataOut_payload_0_16117 : _zz_dataOut_payload_0_15882);
  assign _zz_dataOut_payload_0_16150 = (_zz_dataOut_payload_0_15883 < _zz_dataOut_payload_0_16116);
  assign _zz_dataOut_payload_0_16151 = (_zz_dataOut_payload_0_16150 ? _zz_dataOut_payload_0_15883 : _zz_dataOut_payload_0_16116);
  assign _zz_dataOut_payload_128_11 = (_zz_dataOut_payload_0_16150 ? _zz_dataOut_payload_0_16116 : _zz_dataOut_payload_0_15883);
  assign _zz_dataOut_payload_0_16152 = (_zz_dataOut_payload_0_15884 < _zz_dataOut_payload_0_16115);
  assign _zz_dataOut_payload_0_16153 = (_zz_dataOut_payload_0_16152 ? _zz_dataOut_payload_0_15884 : _zz_dataOut_payload_0_16115);
  assign _zz_dataOut_payload_128_12 = (_zz_dataOut_payload_0_16152 ? _zz_dataOut_payload_0_16115 : _zz_dataOut_payload_0_15884);
  assign _zz_dataOut_payload_0_16154 = (_zz_dataOut_payload_0_15885 < _zz_dataOut_payload_0_16114);
  assign _zz_dataOut_payload_0_16155 = (_zz_dataOut_payload_0_16154 ? _zz_dataOut_payload_0_15885 : _zz_dataOut_payload_0_16114);
  assign _zz_dataOut_payload_128_13 = (_zz_dataOut_payload_0_16154 ? _zz_dataOut_payload_0_16114 : _zz_dataOut_payload_0_15885);
  assign _zz_dataOut_payload_0_16156 = (_zz_dataOut_payload_0_15886 < _zz_dataOut_payload_0_16113);
  assign _zz_dataOut_payload_0_16157 = (_zz_dataOut_payload_0_16156 ? _zz_dataOut_payload_0_15886 : _zz_dataOut_payload_0_16113);
  assign _zz_dataOut_payload_128_14 = (_zz_dataOut_payload_0_16156 ? _zz_dataOut_payload_0_16113 : _zz_dataOut_payload_0_15886);
  assign _zz_dataOut_payload_0_16158 = (_zz_dataOut_payload_0_15887 < _zz_dataOut_payload_0_16112);
  assign _zz_dataOut_payload_0_16159 = (_zz_dataOut_payload_0_16158 ? _zz_dataOut_payload_0_15887 : _zz_dataOut_payload_0_16112);
  assign _zz_dataOut_payload_128_15 = (_zz_dataOut_payload_0_16158 ? _zz_dataOut_payload_0_16112 : _zz_dataOut_payload_0_15887);
  assign _zz_dataOut_payload_0_16160 = (_zz_dataOut_payload_0_15888 < _zz_dataOut_payload_0_16111);
  assign _zz_dataOut_payload_0_16161 = (_zz_dataOut_payload_0_16160 ? _zz_dataOut_payload_0_15888 : _zz_dataOut_payload_0_16111);
  assign _zz_dataOut_payload_128_16 = (_zz_dataOut_payload_0_16160 ? _zz_dataOut_payload_0_16111 : _zz_dataOut_payload_0_15888);
  assign _zz_dataOut_payload_0_16162 = (_zz_dataOut_payload_0_15889 < _zz_dataOut_payload_0_16110);
  assign _zz_dataOut_payload_0_16163 = (_zz_dataOut_payload_0_16162 ? _zz_dataOut_payload_0_15889 : _zz_dataOut_payload_0_16110);
  assign _zz_dataOut_payload_128_17 = (_zz_dataOut_payload_0_16162 ? _zz_dataOut_payload_0_16110 : _zz_dataOut_payload_0_15889);
  assign _zz_dataOut_payload_0_16164 = (_zz_dataOut_payload_0_15890 < _zz_dataOut_payload_0_16109);
  assign _zz_dataOut_payload_0_16165 = (_zz_dataOut_payload_0_16164 ? _zz_dataOut_payload_0_15890 : _zz_dataOut_payload_0_16109);
  assign _zz_dataOut_payload_128_18 = (_zz_dataOut_payload_0_16164 ? _zz_dataOut_payload_0_16109 : _zz_dataOut_payload_0_15890);
  assign _zz_dataOut_payload_0_16166 = (_zz_dataOut_payload_0_15891 < _zz_dataOut_payload_0_16108);
  assign _zz_dataOut_payload_0_16167 = (_zz_dataOut_payload_0_16166 ? _zz_dataOut_payload_0_15891 : _zz_dataOut_payload_0_16108);
  assign _zz_dataOut_payload_128_19 = (_zz_dataOut_payload_0_16166 ? _zz_dataOut_payload_0_16108 : _zz_dataOut_payload_0_15891);
  assign _zz_dataOut_payload_0_16168 = (_zz_dataOut_payload_0_15892 < _zz_dataOut_payload_0_16107);
  assign _zz_dataOut_payload_0_16169 = (_zz_dataOut_payload_0_16168 ? _zz_dataOut_payload_0_15892 : _zz_dataOut_payload_0_16107);
  assign _zz_dataOut_payload_128_20 = (_zz_dataOut_payload_0_16168 ? _zz_dataOut_payload_0_16107 : _zz_dataOut_payload_0_15892);
  assign _zz_dataOut_payload_0_16170 = (_zz_dataOut_payload_0_15893 < _zz_dataOut_payload_0_16106);
  assign _zz_dataOut_payload_0_16171 = (_zz_dataOut_payload_0_16170 ? _zz_dataOut_payload_0_15893 : _zz_dataOut_payload_0_16106);
  assign _zz_dataOut_payload_128_21 = (_zz_dataOut_payload_0_16170 ? _zz_dataOut_payload_0_16106 : _zz_dataOut_payload_0_15893);
  assign _zz_dataOut_payload_0_16172 = (_zz_dataOut_payload_0_15894 < _zz_dataOut_payload_0_16105);
  assign _zz_dataOut_payload_0_16173 = (_zz_dataOut_payload_0_16172 ? _zz_dataOut_payload_0_15894 : _zz_dataOut_payload_0_16105);
  assign _zz_dataOut_payload_128_22 = (_zz_dataOut_payload_0_16172 ? _zz_dataOut_payload_0_16105 : _zz_dataOut_payload_0_15894);
  assign _zz_dataOut_payload_0_16174 = (_zz_dataOut_payload_0_15895 < _zz_dataOut_payload_0_16104);
  assign _zz_dataOut_payload_0_16175 = (_zz_dataOut_payload_0_16174 ? _zz_dataOut_payload_0_15895 : _zz_dataOut_payload_0_16104);
  assign _zz_dataOut_payload_128_23 = (_zz_dataOut_payload_0_16174 ? _zz_dataOut_payload_0_16104 : _zz_dataOut_payload_0_15895);
  assign _zz_dataOut_payload_0_16176 = (_zz_dataOut_payload_0_15896 < _zz_dataOut_payload_0_16103);
  assign _zz_dataOut_payload_0_16177 = (_zz_dataOut_payload_0_16176 ? _zz_dataOut_payload_0_15896 : _zz_dataOut_payload_0_16103);
  assign _zz_dataOut_payload_128_24 = (_zz_dataOut_payload_0_16176 ? _zz_dataOut_payload_0_16103 : _zz_dataOut_payload_0_15896);
  assign _zz_dataOut_payload_0_16178 = (_zz_dataOut_payload_0_15897 < _zz_dataOut_payload_0_16102);
  assign _zz_dataOut_payload_0_16179 = (_zz_dataOut_payload_0_16178 ? _zz_dataOut_payload_0_15897 : _zz_dataOut_payload_0_16102);
  assign _zz_dataOut_payload_128_25 = (_zz_dataOut_payload_0_16178 ? _zz_dataOut_payload_0_16102 : _zz_dataOut_payload_0_15897);
  assign _zz_dataOut_payload_0_16180 = (_zz_dataOut_payload_0_15898 < _zz_dataOut_payload_0_16101);
  assign _zz_dataOut_payload_0_16181 = (_zz_dataOut_payload_0_16180 ? _zz_dataOut_payload_0_15898 : _zz_dataOut_payload_0_16101);
  assign _zz_dataOut_payload_128_26 = (_zz_dataOut_payload_0_16180 ? _zz_dataOut_payload_0_16101 : _zz_dataOut_payload_0_15898);
  assign _zz_dataOut_payload_0_16182 = (_zz_dataOut_payload_0_15899 < _zz_dataOut_payload_0_16100);
  assign _zz_dataOut_payload_0_16183 = (_zz_dataOut_payload_0_16182 ? _zz_dataOut_payload_0_15899 : _zz_dataOut_payload_0_16100);
  assign _zz_dataOut_payload_128_27 = (_zz_dataOut_payload_0_16182 ? _zz_dataOut_payload_0_16100 : _zz_dataOut_payload_0_15899);
  assign _zz_dataOut_payload_0_16184 = (_zz_dataOut_payload_0_15900 < _zz_dataOut_payload_0_16099);
  assign _zz_dataOut_payload_0_16185 = (_zz_dataOut_payload_0_16184 ? _zz_dataOut_payload_0_15900 : _zz_dataOut_payload_0_16099);
  assign _zz_dataOut_payload_128_28 = (_zz_dataOut_payload_0_16184 ? _zz_dataOut_payload_0_16099 : _zz_dataOut_payload_0_15900);
  assign _zz_dataOut_payload_0_16186 = (_zz_dataOut_payload_0_15901 < _zz_dataOut_payload_0_16098);
  assign _zz_dataOut_payload_0_16187 = (_zz_dataOut_payload_0_16186 ? _zz_dataOut_payload_0_15901 : _zz_dataOut_payload_0_16098);
  assign _zz_dataOut_payload_128_29 = (_zz_dataOut_payload_0_16186 ? _zz_dataOut_payload_0_16098 : _zz_dataOut_payload_0_15901);
  assign _zz_dataOut_payload_0_16188 = (_zz_dataOut_payload_0_15902 < _zz_dataOut_payload_0_16097);
  assign _zz_dataOut_payload_0_16189 = (_zz_dataOut_payload_0_16188 ? _zz_dataOut_payload_0_15902 : _zz_dataOut_payload_0_16097);
  assign _zz_dataOut_payload_128_30 = (_zz_dataOut_payload_0_16188 ? _zz_dataOut_payload_0_16097 : _zz_dataOut_payload_0_15902);
  assign _zz_dataOut_payload_0_16190 = (_zz_dataOut_payload_0_15903 < _zz_dataOut_payload_0_16096);
  assign _zz_dataOut_payload_0_16191 = (_zz_dataOut_payload_0_16190 ? _zz_dataOut_payload_0_15903 : _zz_dataOut_payload_0_16096);
  assign _zz_dataOut_payload_128_31 = (_zz_dataOut_payload_0_16190 ? _zz_dataOut_payload_0_16096 : _zz_dataOut_payload_0_15903);
  assign _zz_dataOut_payload_0_16192 = (_zz_dataOut_payload_0_15904 < _zz_dataOut_payload_0_16095);
  assign _zz_dataOut_payload_0_16193 = (_zz_dataOut_payload_0_16192 ? _zz_dataOut_payload_0_15904 : _zz_dataOut_payload_0_16095);
  assign _zz_dataOut_payload_128_32 = (_zz_dataOut_payload_0_16192 ? _zz_dataOut_payload_0_16095 : _zz_dataOut_payload_0_15904);
  assign _zz_dataOut_payload_0_16194 = (_zz_dataOut_payload_0_15905 < _zz_dataOut_payload_0_16094);
  assign _zz_dataOut_payload_0_16195 = (_zz_dataOut_payload_0_16194 ? _zz_dataOut_payload_0_15905 : _zz_dataOut_payload_0_16094);
  assign _zz_dataOut_payload_128_33 = (_zz_dataOut_payload_0_16194 ? _zz_dataOut_payload_0_16094 : _zz_dataOut_payload_0_15905);
  assign _zz_dataOut_payload_0_16196 = (_zz_dataOut_payload_0_15906 < _zz_dataOut_payload_0_16093);
  assign _zz_dataOut_payload_0_16197 = (_zz_dataOut_payload_0_16196 ? _zz_dataOut_payload_0_15906 : _zz_dataOut_payload_0_16093);
  assign _zz_dataOut_payload_128_34 = (_zz_dataOut_payload_0_16196 ? _zz_dataOut_payload_0_16093 : _zz_dataOut_payload_0_15906);
  assign _zz_dataOut_payload_0_16198 = (_zz_dataOut_payload_0_15907 < _zz_dataOut_payload_0_16092);
  assign _zz_dataOut_payload_0_16199 = (_zz_dataOut_payload_0_16198 ? _zz_dataOut_payload_0_15907 : _zz_dataOut_payload_0_16092);
  assign _zz_dataOut_payload_128_35 = (_zz_dataOut_payload_0_16198 ? _zz_dataOut_payload_0_16092 : _zz_dataOut_payload_0_15907);
  assign _zz_dataOut_payload_0_16200 = (_zz_dataOut_payload_0_15908 < _zz_dataOut_payload_0_16091);
  assign _zz_dataOut_payload_0_16201 = (_zz_dataOut_payload_0_16200 ? _zz_dataOut_payload_0_15908 : _zz_dataOut_payload_0_16091);
  assign _zz_dataOut_payload_128_36 = (_zz_dataOut_payload_0_16200 ? _zz_dataOut_payload_0_16091 : _zz_dataOut_payload_0_15908);
  assign _zz_dataOut_payload_0_16202 = (_zz_dataOut_payload_0_15909 < _zz_dataOut_payload_0_16090);
  assign _zz_dataOut_payload_0_16203 = (_zz_dataOut_payload_0_16202 ? _zz_dataOut_payload_0_15909 : _zz_dataOut_payload_0_16090);
  assign _zz_dataOut_payload_128_37 = (_zz_dataOut_payload_0_16202 ? _zz_dataOut_payload_0_16090 : _zz_dataOut_payload_0_15909);
  assign _zz_dataOut_payload_0_16204 = (_zz_dataOut_payload_0_15910 < _zz_dataOut_payload_0_16089);
  assign _zz_dataOut_payload_0_16205 = (_zz_dataOut_payload_0_16204 ? _zz_dataOut_payload_0_15910 : _zz_dataOut_payload_0_16089);
  assign _zz_dataOut_payload_128_38 = (_zz_dataOut_payload_0_16204 ? _zz_dataOut_payload_0_16089 : _zz_dataOut_payload_0_15910);
  assign _zz_dataOut_payload_0_16206 = (_zz_dataOut_payload_0_15911 < _zz_dataOut_payload_0_16088);
  assign _zz_dataOut_payload_0_16207 = (_zz_dataOut_payload_0_16206 ? _zz_dataOut_payload_0_15911 : _zz_dataOut_payload_0_16088);
  assign _zz_dataOut_payload_128_39 = (_zz_dataOut_payload_0_16206 ? _zz_dataOut_payload_0_16088 : _zz_dataOut_payload_0_15911);
  assign _zz_dataOut_payload_0_16208 = (_zz_dataOut_payload_0_15912 < _zz_dataOut_payload_0_16087);
  assign _zz_dataOut_payload_0_16209 = (_zz_dataOut_payload_0_16208 ? _zz_dataOut_payload_0_15912 : _zz_dataOut_payload_0_16087);
  assign _zz_dataOut_payload_128_40 = (_zz_dataOut_payload_0_16208 ? _zz_dataOut_payload_0_16087 : _zz_dataOut_payload_0_15912);
  assign _zz_dataOut_payload_0_16210 = (_zz_dataOut_payload_0_15913 < _zz_dataOut_payload_0_16086);
  assign _zz_dataOut_payload_0_16211 = (_zz_dataOut_payload_0_16210 ? _zz_dataOut_payload_0_15913 : _zz_dataOut_payload_0_16086);
  assign _zz_dataOut_payload_128_41 = (_zz_dataOut_payload_0_16210 ? _zz_dataOut_payload_0_16086 : _zz_dataOut_payload_0_15913);
  assign _zz_dataOut_payload_0_16212 = (_zz_dataOut_payload_0_15914 < _zz_dataOut_payload_0_16085);
  assign _zz_dataOut_payload_0_16213 = (_zz_dataOut_payload_0_16212 ? _zz_dataOut_payload_0_15914 : _zz_dataOut_payload_0_16085);
  assign _zz_dataOut_payload_128_42 = (_zz_dataOut_payload_0_16212 ? _zz_dataOut_payload_0_16085 : _zz_dataOut_payload_0_15914);
  assign _zz_dataOut_payload_0_16214 = (_zz_dataOut_payload_0_15915 < _zz_dataOut_payload_0_16084);
  assign _zz_dataOut_payload_0_16215 = (_zz_dataOut_payload_0_16214 ? _zz_dataOut_payload_0_15915 : _zz_dataOut_payload_0_16084);
  assign _zz_dataOut_payload_128_43 = (_zz_dataOut_payload_0_16214 ? _zz_dataOut_payload_0_16084 : _zz_dataOut_payload_0_15915);
  assign _zz_dataOut_payload_0_16216 = (_zz_dataOut_payload_0_15916 < _zz_dataOut_payload_0_16083);
  assign _zz_dataOut_payload_0_16217 = (_zz_dataOut_payload_0_16216 ? _zz_dataOut_payload_0_15916 : _zz_dataOut_payload_0_16083);
  assign _zz_dataOut_payload_128_44 = (_zz_dataOut_payload_0_16216 ? _zz_dataOut_payload_0_16083 : _zz_dataOut_payload_0_15916);
  assign _zz_dataOut_payload_0_16218 = (_zz_dataOut_payload_0_15917 < _zz_dataOut_payload_0_16082);
  assign _zz_dataOut_payload_0_16219 = (_zz_dataOut_payload_0_16218 ? _zz_dataOut_payload_0_15917 : _zz_dataOut_payload_0_16082);
  assign _zz_dataOut_payload_128_45 = (_zz_dataOut_payload_0_16218 ? _zz_dataOut_payload_0_16082 : _zz_dataOut_payload_0_15917);
  assign _zz_dataOut_payload_0_16220 = (_zz_dataOut_payload_0_15918 < _zz_dataOut_payload_0_16081);
  assign _zz_dataOut_payload_0_16221 = (_zz_dataOut_payload_0_16220 ? _zz_dataOut_payload_0_15918 : _zz_dataOut_payload_0_16081);
  assign _zz_dataOut_payload_128_46 = (_zz_dataOut_payload_0_16220 ? _zz_dataOut_payload_0_16081 : _zz_dataOut_payload_0_15918);
  assign _zz_dataOut_payload_0_16222 = (_zz_dataOut_payload_0_15919 < _zz_dataOut_payload_0_16080);
  assign _zz_dataOut_payload_0_16223 = (_zz_dataOut_payload_0_16222 ? _zz_dataOut_payload_0_15919 : _zz_dataOut_payload_0_16080);
  assign _zz_dataOut_payload_128_47 = (_zz_dataOut_payload_0_16222 ? _zz_dataOut_payload_0_16080 : _zz_dataOut_payload_0_15919);
  assign _zz_dataOut_payload_0_16224 = (_zz_dataOut_payload_0_15920 < _zz_dataOut_payload_0_16079);
  assign _zz_dataOut_payload_0_16225 = (_zz_dataOut_payload_0_16224 ? _zz_dataOut_payload_0_15920 : _zz_dataOut_payload_0_16079);
  assign _zz_dataOut_payload_128_48 = (_zz_dataOut_payload_0_16224 ? _zz_dataOut_payload_0_16079 : _zz_dataOut_payload_0_15920);
  assign _zz_dataOut_payload_0_16226 = (_zz_dataOut_payload_0_15921 < _zz_dataOut_payload_0_16078);
  assign _zz_dataOut_payload_0_16227 = (_zz_dataOut_payload_0_16226 ? _zz_dataOut_payload_0_15921 : _zz_dataOut_payload_0_16078);
  assign _zz_dataOut_payload_128_49 = (_zz_dataOut_payload_0_16226 ? _zz_dataOut_payload_0_16078 : _zz_dataOut_payload_0_15921);
  assign _zz_dataOut_payload_0_16228 = (_zz_dataOut_payload_0_15922 < _zz_dataOut_payload_0_16077);
  assign _zz_dataOut_payload_0_16229 = (_zz_dataOut_payload_0_16228 ? _zz_dataOut_payload_0_15922 : _zz_dataOut_payload_0_16077);
  assign _zz_dataOut_payload_128_50 = (_zz_dataOut_payload_0_16228 ? _zz_dataOut_payload_0_16077 : _zz_dataOut_payload_0_15922);
  assign _zz_dataOut_payload_0_16230 = (_zz_dataOut_payload_0_15923 < _zz_dataOut_payload_0_16076);
  assign _zz_dataOut_payload_0_16231 = (_zz_dataOut_payload_0_16230 ? _zz_dataOut_payload_0_15923 : _zz_dataOut_payload_0_16076);
  assign _zz_dataOut_payload_128_51 = (_zz_dataOut_payload_0_16230 ? _zz_dataOut_payload_0_16076 : _zz_dataOut_payload_0_15923);
  assign _zz_dataOut_payload_0_16232 = (_zz_dataOut_payload_0_15924 < _zz_dataOut_payload_0_16075);
  assign _zz_dataOut_payload_0_16233 = (_zz_dataOut_payload_0_16232 ? _zz_dataOut_payload_0_15924 : _zz_dataOut_payload_0_16075);
  assign _zz_dataOut_payload_128_52 = (_zz_dataOut_payload_0_16232 ? _zz_dataOut_payload_0_16075 : _zz_dataOut_payload_0_15924);
  assign _zz_dataOut_payload_0_16234 = (_zz_dataOut_payload_0_15925 < _zz_dataOut_payload_0_16074);
  assign _zz_dataOut_payload_0_16235 = (_zz_dataOut_payload_0_16234 ? _zz_dataOut_payload_0_15925 : _zz_dataOut_payload_0_16074);
  assign _zz_dataOut_payload_128_53 = (_zz_dataOut_payload_0_16234 ? _zz_dataOut_payload_0_16074 : _zz_dataOut_payload_0_15925);
  assign _zz_dataOut_payload_0_16236 = (_zz_dataOut_payload_0_15926 < _zz_dataOut_payload_0_16073);
  assign _zz_dataOut_payload_0_16237 = (_zz_dataOut_payload_0_16236 ? _zz_dataOut_payload_0_15926 : _zz_dataOut_payload_0_16073);
  assign _zz_dataOut_payload_128_54 = (_zz_dataOut_payload_0_16236 ? _zz_dataOut_payload_0_16073 : _zz_dataOut_payload_0_15926);
  assign _zz_dataOut_payload_0_16238 = (_zz_dataOut_payload_0_15927 < _zz_dataOut_payload_0_16072);
  assign _zz_dataOut_payload_0_16239 = (_zz_dataOut_payload_0_16238 ? _zz_dataOut_payload_0_15927 : _zz_dataOut_payload_0_16072);
  assign _zz_dataOut_payload_128_55 = (_zz_dataOut_payload_0_16238 ? _zz_dataOut_payload_0_16072 : _zz_dataOut_payload_0_15927);
  assign _zz_dataOut_payload_0_16240 = (_zz_dataOut_payload_0_15928 < _zz_dataOut_payload_0_16071);
  assign _zz_dataOut_payload_0_16241 = (_zz_dataOut_payload_0_16240 ? _zz_dataOut_payload_0_15928 : _zz_dataOut_payload_0_16071);
  assign _zz_dataOut_payload_128_56 = (_zz_dataOut_payload_0_16240 ? _zz_dataOut_payload_0_16071 : _zz_dataOut_payload_0_15928);
  assign _zz_dataOut_payload_0_16242 = (_zz_dataOut_payload_0_15929 < _zz_dataOut_payload_0_16070);
  assign _zz_dataOut_payload_0_16243 = (_zz_dataOut_payload_0_16242 ? _zz_dataOut_payload_0_15929 : _zz_dataOut_payload_0_16070);
  assign _zz_dataOut_payload_128_57 = (_zz_dataOut_payload_0_16242 ? _zz_dataOut_payload_0_16070 : _zz_dataOut_payload_0_15929);
  assign _zz_dataOut_payload_0_16244 = (_zz_dataOut_payload_0_15930 < _zz_dataOut_payload_0_16069);
  assign _zz_dataOut_payload_0_16245 = (_zz_dataOut_payload_0_16244 ? _zz_dataOut_payload_0_15930 : _zz_dataOut_payload_0_16069);
  assign _zz_dataOut_payload_128_58 = (_zz_dataOut_payload_0_16244 ? _zz_dataOut_payload_0_16069 : _zz_dataOut_payload_0_15930);
  assign _zz_dataOut_payload_0_16246 = (_zz_dataOut_payload_0_15931 < _zz_dataOut_payload_0_16068);
  assign _zz_dataOut_payload_0_16247 = (_zz_dataOut_payload_0_16246 ? _zz_dataOut_payload_0_15931 : _zz_dataOut_payload_0_16068);
  assign _zz_dataOut_payload_128_59 = (_zz_dataOut_payload_0_16246 ? _zz_dataOut_payload_0_16068 : _zz_dataOut_payload_0_15931);
  assign _zz_dataOut_payload_0_16248 = (_zz_dataOut_payload_0_15932 < _zz_dataOut_payload_0_16067);
  assign _zz_dataOut_payload_0_16249 = (_zz_dataOut_payload_0_16248 ? _zz_dataOut_payload_0_15932 : _zz_dataOut_payload_0_16067);
  assign _zz_dataOut_payload_128_60 = (_zz_dataOut_payload_0_16248 ? _zz_dataOut_payload_0_16067 : _zz_dataOut_payload_0_15932);
  assign _zz_dataOut_payload_0_16250 = (_zz_dataOut_payload_0_15933 < _zz_dataOut_payload_0_16066);
  assign _zz_dataOut_payload_0_16251 = (_zz_dataOut_payload_0_16250 ? _zz_dataOut_payload_0_15933 : _zz_dataOut_payload_0_16066);
  assign _zz_dataOut_payload_128_61 = (_zz_dataOut_payload_0_16250 ? _zz_dataOut_payload_0_16066 : _zz_dataOut_payload_0_15933);
  assign _zz_dataOut_payload_0_16252 = (_zz_dataOut_payload_0_15934 < _zz_dataOut_payload_0_16065);
  assign _zz_dataOut_payload_0_16253 = (_zz_dataOut_payload_0_16252 ? _zz_dataOut_payload_0_15934 : _zz_dataOut_payload_0_16065);
  assign _zz_dataOut_payload_128_62 = (_zz_dataOut_payload_0_16252 ? _zz_dataOut_payload_0_16065 : _zz_dataOut_payload_0_15934);
  assign _zz_dataOut_payload_0_16254 = (_zz_dataOut_payload_0_15935 < _zz_dataOut_payload_0_16064);
  assign _zz_dataOut_payload_0_16255 = (_zz_dataOut_payload_0_16254 ? _zz_dataOut_payload_0_15935 : _zz_dataOut_payload_0_16064);
  assign _zz_dataOut_payload_128_63 = (_zz_dataOut_payload_0_16254 ? _zz_dataOut_payload_0_16064 : _zz_dataOut_payload_0_15935);
  assign _zz_dataOut_payload_0_16256 = (_zz_dataOut_payload_0_15936 < _zz_dataOut_payload_0_16063);
  assign _zz_dataOut_payload_0_16257 = (_zz_dataOut_payload_0_16256 ? _zz_dataOut_payload_0_15936 : _zz_dataOut_payload_0_16063);
  assign _zz_dataOut_payload_128_64 = (_zz_dataOut_payload_0_16256 ? _zz_dataOut_payload_0_16063 : _zz_dataOut_payload_0_15936);
  assign _zz_dataOut_payload_0_16258 = (_zz_dataOut_payload_0_15937 < _zz_dataOut_payload_0_16062);
  assign _zz_dataOut_payload_0_16259 = (_zz_dataOut_payload_0_16258 ? _zz_dataOut_payload_0_15937 : _zz_dataOut_payload_0_16062);
  assign _zz_dataOut_payload_128_65 = (_zz_dataOut_payload_0_16258 ? _zz_dataOut_payload_0_16062 : _zz_dataOut_payload_0_15937);
  assign _zz_dataOut_payload_0_16260 = (_zz_dataOut_payload_0_15938 < _zz_dataOut_payload_0_16061);
  assign _zz_dataOut_payload_0_16261 = (_zz_dataOut_payload_0_16260 ? _zz_dataOut_payload_0_15938 : _zz_dataOut_payload_0_16061);
  assign _zz_dataOut_payload_128_66 = (_zz_dataOut_payload_0_16260 ? _zz_dataOut_payload_0_16061 : _zz_dataOut_payload_0_15938);
  assign _zz_dataOut_payload_0_16262 = (_zz_dataOut_payload_0_15939 < _zz_dataOut_payload_0_16060);
  assign _zz_dataOut_payload_0_16263 = (_zz_dataOut_payload_0_16262 ? _zz_dataOut_payload_0_15939 : _zz_dataOut_payload_0_16060);
  assign _zz_dataOut_payload_128_67 = (_zz_dataOut_payload_0_16262 ? _zz_dataOut_payload_0_16060 : _zz_dataOut_payload_0_15939);
  assign _zz_dataOut_payload_0_16264 = (_zz_dataOut_payload_0_15940 < _zz_dataOut_payload_0_16059);
  assign _zz_dataOut_payload_0_16265 = (_zz_dataOut_payload_0_16264 ? _zz_dataOut_payload_0_15940 : _zz_dataOut_payload_0_16059);
  assign _zz_dataOut_payload_128_68 = (_zz_dataOut_payload_0_16264 ? _zz_dataOut_payload_0_16059 : _zz_dataOut_payload_0_15940);
  assign _zz_dataOut_payload_0_16266 = (_zz_dataOut_payload_0_15941 < _zz_dataOut_payload_0_16058);
  assign _zz_dataOut_payload_0_16267 = (_zz_dataOut_payload_0_16266 ? _zz_dataOut_payload_0_15941 : _zz_dataOut_payload_0_16058);
  assign _zz_dataOut_payload_128_69 = (_zz_dataOut_payload_0_16266 ? _zz_dataOut_payload_0_16058 : _zz_dataOut_payload_0_15941);
  assign _zz_dataOut_payload_0_16268 = (_zz_dataOut_payload_0_15942 < _zz_dataOut_payload_0_16057);
  assign _zz_dataOut_payload_0_16269 = (_zz_dataOut_payload_0_16268 ? _zz_dataOut_payload_0_15942 : _zz_dataOut_payload_0_16057);
  assign _zz_dataOut_payload_128_70 = (_zz_dataOut_payload_0_16268 ? _zz_dataOut_payload_0_16057 : _zz_dataOut_payload_0_15942);
  assign _zz_dataOut_payload_0_16270 = (_zz_dataOut_payload_0_15943 < _zz_dataOut_payload_0_16056);
  assign _zz_dataOut_payload_0_16271 = (_zz_dataOut_payload_0_16270 ? _zz_dataOut_payload_0_15943 : _zz_dataOut_payload_0_16056);
  assign _zz_dataOut_payload_128_71 = (_zz_dataOut_payload_0_16270 ? _zz_dataOut_payload_0_16056 : _zz_dataOut_payload_0_15943);
  assign _zz_dataOut_payload_0_16272 = (_zz_dataOut_payload_0_15944 < _zz_dataOut_payload_0_16055);
  assign _zz_dataOut_payload_0_16273 = (_zz_dataOut_payload_0_16272 ? _zz_dataOut_payload_0_15944 : _zz_dataOut_payload_0_16055);
  assign _zz_dataOut_payload_128_72 = (_zz_dataOut_payload_0_16272 ? _zz_dataOut_payload_0_16055 : _zz_dataOut_payload_0_15944);
  assign _zz_dataOut_payload_0_16274 = (_zz_dataOut_payload_0_15945 < _zz_dataOut_payload_0_16054);
  assign _zz_dataOut_payload_0_16275 = (_zz_dataOut_payload_0_16274 ? _zz_dataOut_payload_0_15945 : _zz_dataOut_payload_0_16054);
  assign _zz_dataOut_payload_128_73 = (_zz_dataOut_payload_0_16274 ? _zz_dataOut_payload_0_16054 : _zz_dataOut_payload_0_15945);
  assign _zz_dataOut_payload_0_16276 = (_zz_dataOut_payload_0_15946 < _zz_dataOut_payload_0_16053);
  assign _zz_dataOut_payload_0_16277 = (_zz_dataOut_payload_0_16276 ? _zz_dataOut_payload_0_15946 : _zz_dataOut_payload_0_16053);
  assign _zz_dataOut_payload_128_74 = (_zz_dataOut_payload_0_16276 ? _zz_dataOut_payload_0_16053 : _zz_dataOut_payload_0_15946);
  assign _zz_dataOut_payload_0_16278 = (_zz_dataOut_payload_0_15947 < _zz_dataOut_payload_0_16052);
  assign _zz_dataOut_payload_0_16279 = (_zz_dataOut_payload_0_16278 ? _zz_dataOut_payload_0_15947 : _zz_dataOut_payload_0_16052);
  assign _zz_dataOut_payload_128_75 = (_zz_dataOut_payload_0_16278 ? _zz_dataOut_payload_0_16052 : _zz_dataOut_payload_0_15947);
  assign _zz_dataOut_payload_0_16280 = (_zz_dataOut_payload_0_15948 < _zz_dataOut_payload_0_16051);
  assign _zz_dataOut_payload_0_16281 = (_zz_dataOut_payload_0_16280 ? _zz_dataOut_payload_0_15948 : _zz_dataOut_payload_0_16051);
  assign _zz_dataOut_payload_128_76 = (_zz_dataOut_payload_0_16280 ? _zz_dataOut_payload_0_16051 : _zz_dataOut_payload_0_15948);
  assign _zz_dataOut_payload_0_16282 = (_zz_dataOut_payload_0_15949 < _zz_dataOut_payload_0_16050);
  assign _zz_dataOut_payload_0_16283 = (_zz_dataOut_payload_0_16282 ? _zz_dataOut_payload_0_15949 : _zz_dataOut_payload_0_16050);
  assign _zz_dataOut_payload_128_77 = (_zz_dataOut_payload_0_16282 ? _zz_dataOut_payload_0_16050 : _zz_dataOut_payload_0_15949);
  assign _zz_dataOut_payload_0_16284 = (_zz_dataOut_payload_0_15950 < _zz_dataOut_payload_0_16049);
  assign _zz_dataOut_payload_0_16285 = (_zz_dataOut_payload_0_16284 ? _zz_dataOut_payload_0_15950 : _zz_dataOut_payload_0_16049);
  assign _zz_dataOut_payload_128_78 = (_zz_dataOut_payload_0_16284 ? _zz_dataOut_payload_0_16049 : _zz_dataOut_payload_0_15950);
  assign _zz_dataOut_payload_0_16286 = (_zz_dataOut_payload_0_15951 < _zz_dataOut_payload_0_16048);
  assign _zz_dataOut_payload_0_16287 = (_zz_dataOut_payload_0_16286 ? _zz_dataOut_payload_0_15951 : _zz_dataOut_payload_0_16048);
  assign _zz_dataOut_payload_128_79 = (_zz_dataOut_payload_0_16286 ? _zz_dataOut_payload_0_16048 : _zz_dataOut_payload_0_15951);
  assign _zz_dataOut_payload_0_16288 = (_zz_dataOut_payload_0_15952 < _zz_dataOut_payload_0_16047);
  assign _zz_dataOut_payload_0_16289 = (_zz_dataOut_payload_0_16288 ? _zz_dataOut_payload_0_15952 : _zz_dataOut_payload_0_16047);
  assign _zz_dataOut_payload_128_80 = (_zz_dataOut_payload_0_16288 ? _zz_dataOut_payload_0_16047 : _zz_dataOut_payload_0_15952);
  assign _zz_dataOut_payload_0_16290 = (_zz_dataOut_payload_0_15953 < _zz_dataOut_payload_0_16046);
  assign _zz_dataOut_payload_0_16291 = (_zz_dataOut_payload_0_16290 ? _zz_dataOut_payload_0_15953 : _zz_dataOut_payload_0_16046);
  assign _zz_dataOut_payload_128_81 = (_zz_dataOut_payload_0_16290 ? _zz_dataOut_payload_0_16046 : _zz_dataOut_payload_0_15953);
  assign _zz_dataOut_payload_0_16292 = (_zz_dataOut_payload_0_15954 < _zz_dataOut_payload_0_16045);
  assign _zz_dataOut_payload_0_16293 = (_zz_dataOut_payload_0_16292 ? _zz_dataOut_payload_0_15954 : _zz_dataOut_payload_0_16045);
  assign _zz_dataOut_payload_128_82 = (_zz_dataOut_payload_0_16292 ? _zz_dataOut_payload_0_16045 : _zz_dataOut_payload_0_15954);
  assign _zz_dataOut_payload_0_16294 = (_zz_dataOut_payload_0_15955 < _zz_dataOut_payload_0_16044);
  assign _zz_dataOut_payload_0_16295 = (_zz_dataOut_payload_0_16294 ? _zz_dataOut_payload_0_15955 : _zz_dataOut_payload_0_16044);
  assign _zz_dataOut_payload_128_83 = (_zz_dataOut_payload_0_16294 ? _zz_dataOut_payload_0_16044 : _zz_dataOut_payload_0_15955);
  assign _zz_dataOut_payload_0_16296 = (_zz_dataOut_payload_0_15956 < _zz_dataOut_payload_0_16043);
  assign _zz_dataOut_payload_0_16297 = (_zz_dataOut_payload_0_16296 ? _zz_dataOut_payload_0_15956 : _zz_dataOut_payload_0_16043);
  assign _zz_dataOut_payload_128_84 = (_zz_dataOut_payload_0_16296 ? _zz_dataOut_payload_0_16043 : _zz_dataOut_payload_0_15956);
  assign _zz_dataOut_payload_0_16298 = (_zz_dataOut_payload_0_15957 < _zz_dataOut_payload_0_16042);
  assign _zz_dataOut_payload_0_16299 = (_zz_dataOut_payload_0_16298 ? _zz_dataOut_payload_0_15957 : _zz_dataOut_payload_0_16042);
  assign _zz_dataOut_payload_128_85 = (_zz_dataOut_payload_0_16298 ? _zz_dataOut_payload_0_16042 : _zz_dataOut_payload_0_15957);
  assign _zz_dataOut_payload_0_16300 = (_zz_dataOut_payload_0_15958 < _zz_dataOut_payload_0_16041);
  assign _zz_dataOut_payload_0_16301 = (_zz_dataOut_payload_0_16300 ? _zz_dataOut_payload_0_15958 : _zz_dataOut_payload_0_16041);
  assign _zz_dataOut_payload_128_86 = (_zz_dataOut_payload_0_16300 ? _zz_dataOut_payload_0_16041 : _zz_dataOut_payload_0_15958);
  assign _zz_dataOut_payload_0_16302 = (_zz_dataOut_payload_0_15959 < _zz_dataOut_payload_0_16040);
  assign _zz_dataOut_payload_0_16303 = (_zz_dataOut_payload_0_16302 ? _zz_dataOut_payload_0_15959 : _zz_dataOut_payload_0_16040);
  assign _zz_dataOut_payload_128_87 = (_zz_dataOut_payload_0_16302 ? _zz_dataOut_payload_0_16040 : _zz_dataOut_payload_0_15959);
  assign _zz_dataOut_payload_0_16304 = (_zz_dataOut_payload_0_15960 < _zz_dataOut_payload_0_16039);
  assign _zz_dataOut_payload_0_16305 = (_zz_dataOut_payload_0_16304 ? _zz_dataOut_payload_0_15960 : _zz_dataOut_payload_0_16039);
  assign _zz_dataOut_payload_128_88 = (_zz_dataOut_payload_0_16304 ? _zz_dataOut_payload_0_16039 : _zz_dataOut_payload_0_15960);
  assign _zz_dataOut_payload_0_16306 = (_zz_dataOut_payload_0_15961 < _zz_dataOut_payload_0_16038);
  assign _zz_dataOut_payload_0_16307 = (_zz_dataOut_payload_0_16306 ? _zz_dataOut_payload_0_15961 : _zz_dataOut_payload_0_16038);
  assign _zz_dataOut_payload_128_89 = (_zz_dataOut_payload_0_16306 ? _zz_dataOut_payload_0_16038 : _zz_dataOut_payload_0_15961);
  assign _zz_dataOut_payload_0_16308 = (_zz_dataOut_payload_0_15962 < _zz_dataOut_payload_0_16037);
  assign _zz_dataOut_payload_0_16309 = (_zz_dataOut_payload_0_16308 ? _zz_dataOut_payload_0_15962 : _zz_dataOut_payload_0_16037);
  assign _zz_dataOut_payload_128_90 = (_zz_dataOut_payload_0_16308 ? _zz_dataOut_payload_0_16037 : _zz_dataOut_payload_0_15962);
  assign _zz_dataOut_payload_0_16310 = (_zz_dataOut_payload_0_15963 < _zz_dataOut_payload_0_16036);
  assign _zz_dataOut_payload_0_16311 = (_zz_dataOut_payload_0_16310 ? _zz_dataOut_payload_0_15963 : _zz_dataOut_payload_0_16036);
  assign _zz_dataOut_payload_128_91 = (_zz_dataOut_payload_0_16310 ? _zz_dataOut_payload_0_16036 : _zz_dataOut_payload_0_15963);
  assign _zz_dataOut_payload_0_16312 = (_zz_dataOut_payload_0_15964 < _zz_dataOut_payload_0_16035);
  assign _zz_dataOut_payload_0_16313 = (_zz_dataOut_payload_0_16312 ? _zz_dataOut_payload_0_15964 : _zz_dataOut_payload_0_16035);
  assign _zz_dataOut_payload_128_92 = (_zz_dataOut_payload_0_16312 ? _zz_dataOut_payload_0_16035 : _zz_dataOut_payload_0_15964);
  assign _zz_dataOut_payload_0_16314 = (_zz_dataOut_payload_0_15965 < _zz_dataOut_payload_0_16034);
  assign _zz_dataOut_payload_0_16315 = (_zz_dataOut_payload_0_16314 ? _zz_dataOut_payload_0_15965 : _zz_dataOut_payload_0_16034);
  assign _zz_dataOut_payload_128_93 = (_zz_dataOut_payload_0_16314 ? _zz_dataOut_payload_0_16034 : _zz_dataOut_payload_0_15965);
  assign _zz_dataOut_payload_0_16316 = (_zz_dataOut_payload_0_15966 < _zz_dataOut_payload_0_16033);
  assign _zz_dataOut_payload_0_16317 = (_zz_dataOut_payload_0_16316 ? _zz_dataOut_payload_0_15966 : _zz_dataOut_payload_0_16033);
  assign _zz_dataOut_payload_128_94 = (_zz_dataOut_payload_0_16316 ? _zz_dataOut_payload_0_16033 : _zz_dataOut_payload_0_15966);
  assign _zz_dataOut_payload_0_16318 = (_zz_dataOut_payload_0_15967 < _zz_dataOut_payload_0_16032);
  assign _zz_dataOut_payload_0_16319 = (_zz_dataOut_payload_0_16318 ? _zz_dataOut_payload_0_15967 : _zz_dataOut_payload_0_16032);
  assign _zz_dataOut_payload_128_95 = (_zz_dataOut_payload_0_16318 ? _zz_dataOut_payload_0_16032 : _zz_dataOut_payload_0_15967);
  assign _zz_dataOut_payload_0_16320 = (_zz_dataOut_payload_0_15968 < _zz_dataOut_payload_0_16031);
  assign _zz_dataOut_payload_0_16321 = (_zz_dataOut_payload_0_16320 ? _zz_dataOut_payload_0_15968 : _zz_dataOut_payload_0_16031);
  assign _zz_dataOut_payload_128_96 = (_zz_dataOut_payload_0_16320 ? _zz_dataOut_payload_0_16031 : _zz_dataOut_payload_0_15968);
  assign _zz_dataOut_payload_0_16322 = (_zz_dataOut_payload_0_15969 < _zz_dataOut_payload_0_16030);
  assign _zz_dataOut_payload_0_16323 = (_zz_dataOut_payload_0_16322 ? _zz_dataOut_payload_0_15969 : _zz_dataOut_payload_0_16030);
  assign _zz_dataOut_payload_128_97 = (_zz_dataOut_payload_0_16322 ? _zz_dataOut_payload_0_16030 : _zz_dataOut_payload_0_15969);
  assign _zz_dataOut_payload_0_16324 = (_zz_dataOut_payload_0_15970 < _zz_dataOut_payload_0_16029);
  assign _zz_dataOut_payload_0_16325 = (_zz_dataOut_payload_0_16324 ? _zz_dataOut_payload_0_15970 : _zz_dataOut_payload_0_16029);
  assign _zz_dataOut_payload_128_98 = (_zz_dataOut_payload_0_16324 ? _zz_dataOut_payload_0_16029 : _zz_dataOut_payload_0_15970);
  assign _zz_dataOut_payload_0_16326 = (_zz_dataOut_payload_0_15971 < _zz_dataOut_payload_0_16028);
  assign _zz_dataOut_payload_0_16327 = (_zz_dataOut_payload_0_16326 ? _zz_dataOut_payload_0_15971 : _zz_dataOut_payload_0_16028);
  assign _zz_dataOut_payload_128_99 = (_zz_dataOut_payload_0_16326 ? _zz_dataOut_payload_0_16028 : _zz_dataOut_payload_0_15971);
  assign _zz_dataOut_payload_0_16328 = (_zz_dataOut_payload_0_15972 < _zz_dataOut_payload_0_16027);
  assign _zz_dataOut_payload_0_16329 = (_zz_dataOut_payload_0_16328 ? _zz_dataOut_payload_0_15972 : _zz_dataOut_payload_0_16027);
  assign _zz_dataOut_payload_128_100 = (_zz_dataOut_payload_0_16328 ? _zz_dataOut_payload_0_16027 : _zz_dataOut_payload_0_15972);
  assign _zz_dataOut_payload_0_16330 = (_zz_dataOut_payload_0_15973 < _zz_dataOut_payload_0_16026);
  assign _zz_dataOut_payload_0_16331 = (_zz_dataOut_payload_0_16330 ? _zz_dataOut_payload_0_15973 : _zz_dataOut_payload_0_16026);
  assign _zz_dataOut_payload_128_101 = (_zz_dataOut_payload_0_16330 ? _zz_dataOut_payload_0_16026 : _zz_dataOut_payload_0_15973);
  assign _zz_dataOut_payload_0_16332 = (_zz_dataOut_payload_0_15974 < _zz_dataOut_payload_0_16025);
  assign _zz_dataOut_payload_0_16333 = (_zz_dataOut_payload_0_16332 ? _zz_dataOut_payload_0_15974 : _zz_dataOut_payload_0_16025);
  assign _zz_dataOut_payload_128_102 = (_zz_dataOut_payload_0_16332 ? _zz_dataOut_payload_0_16025 : _zz_dataOut_payload_0_15974);
  assign _zz_dataOut_payload_0_16334 = (_zz_dataOut_payload_0_15975 < _zz_dataOut_payload_0_16024);
  assign _zz_dataOut_payload_0_16335 = (_zz_dataOut_payload_0_16334 ? _zz_dataOut_payload_0_15975 : _zz_dataOut_payload_0_16024);
  assign _zz_dataOut_payload_128_103 = (_zz_dataOut_payload_0_16334 ? _zz_dataOut_payload_0_16024 : _zz_dataOut_payload_0_15975);
  assign _zz_dataOut_payload_0_16336 = (_zz_dataOut_payload_0_15976 < _zz_dataOut_payload_0_16023);
  assign _zz_dataOut_payload_0_16337 = (_zz_dataOut_payload_0_16336 ? _zz_dataOut_payload_0_15976 : _zz_dataOut_payload_0_16023);
  assign _zz_dataOut_payload_128_104 = (_zz_dataOut_payload_0_16336 ? _zz_dataOut_payload_0_16023 : _zz_dataOut_payload_0_15976);
  assign _zz_dataOut_payload_0_16338 = (_zz_dataOut_payload_0_15977 < _zz_dataOut_payload_0_16022);
  assign _zz_dataOut_payload_0_16339 = (_zz_dataOut_payload_0_16338 ? _zz_dataOut_payload_0_15977 : _zz_dataOut_payload_0_16022);
  assign _zz_dataOut_payload_128_105 = (_zz_dataOut_payload_0_16338 ? _zz_dataOut_payload_0_16022 : _zz_dataOut_payload_0_15977);
  assign _zz_dataOut_payload_0_16340 = (_zz_dataOut_payload_0_15978 < _zz_dataOut_payload_0_16021);
  assign _zz_dataOut_payload_0_16341 = (_zz_dataOut_payload_0_16340 ? _zz_dataOut_payload_0_15978 : _zz_dataOut_payload_0_16021);
  assign _zz_dataOut_payload_128_106 = (_zz_dataOut_payload_0_16340 ? _zz_dataOut_payload_0_16021 : _zz_dataOut_payload_0_15978);
  assign _zz_dataOut_payload_0_16342 = (_zz_dataOut_payload_0_15979 < _zz_dataOut_payload_0_16020);
  assign _zz_dataOut_payload_0_16343 = (_zz_dataOut_payload_0_16342 ? _zz_dataOut_payload_0_15979 : _zz_dataOut_payload_0_16020);
  assign _zz_dataOut_payload_128_107 = (_zz_dataOut_payload_0_16342 ? _zz_dataOut_payload_0_16020 : _zz_dataOut_payload_0_15979);
  assign _zz_dataOut_payload_0_16344 = (_zz_dataOut_payload_0_15980 < _zz_dataOut_payload_0_16019);
  assign _zz_dataOut_payload_0_16345 = (_zz_dataOut_payload_0_16344 ? _zz_dataOut_payload_0_15980 : _zz_dataOut_payload_0_16019);
  assign _zz_dataOut_payload_128_108 = (_zz_dataOut_payload_0_16344 ? _zz_dataOut_payload_0_16019 : _zz_dataOut_payload_0_15980);
  assign _zz_dataOut_payload_0_16346 = (_zz_dataOut_payload_0_15981 < _zz_dataOut_payload_0_16018);
  assign _zz_dataOut_payload_0_16347 = (_zz_dataOut_payload_0_16346 ? _zz_dataOut_payload_0_15981 : _zz_dataOut_payload_0_16018);
  assign _zz_dataOut_payload_128_109 = (_zz_dataOut_payload_0_16346 ? _zz_dataOut_payload_0_16018 : _zz_dataOut_payload_0_15981);
  assign _zz_dataOut_payload_0_16348 = (_zz_dataOut_payload_0_15982 < _zz_dataOut_payload_0_16017);
  assign _zz_dataOut_payload_0_16349 = (_zz_dataOut_payload_0_16348 ? _zz_dataOut_payload_0_15982 : _zz_dataOut_payload_0_16017);
  assign _zz_dataOut_payload_128_110 = (_zz_dataOut_payload_0_16348 ? _zz_dataOut_payload_0_16017 : _zz_dataOut_payload_0_15982);
  assign _zz_dataOut_payload_0_16350 = (_zz_dataOut_payload_0_15983 < _zz_dataOut_payload_0_16016);
  assign _zz_dataOut_payload_0_16351 = (_zz_dataOut_payload_0_16350 ? _zz_dataOut_payload_0_15983 : _zz_dataOut_payload_0_16016);
  assign _zz_dataOut_payload_128_111 = (_zz_dataOut_payload_0_16350 ? _zz_dataOut_payload_0_16016 : _zz_dataOut_payload_0_15983);
  assign _zz_dataOut_payload_0_16352 = (_zz_dataOut_payload_0_15984 < _zz_dataOut_payload_0_16015);
  assign _zz_dataOut_payload_0_16353 = (_zz_dataOut_payload_0_16352 ? _zz_dataOut_payload_0_15984 : _zz_dataOut_payload_0_16015);
  assign _zz_dataOut_payload_128_112 = (_zz_dataOut_payload_0_16352 ? _zz_dataOut_payload_0_16015 : _zz_dataOut_payload_0_15984);
  assign _zz_dataOut_payload_0_16354 = (_zz_dataOut_payload_0_15985 < _zz_dataOut_payload_0_16014);
  assign _zz_dataOut_payload_0_16355 = (_zz_dataOut_payload_0_16354 ? _zz_dataOut_payload_0_15985 : _zz_dataOut_payload_0_16014);
  assign _zz_dataOut_payload_128_113 = (_zz_dataOut_payload_0_16354 ? _zz_dataOut_payload_0_16014 : _zz_dataOut_payload_0_15985);
  assign _zz_dataOut_payload_0_16356 = (_zz_dataOut_payload_0_15986 < _zz_dataOut_payload_0_16013);
  assign _zz_dataOut_payload_0_16357 = (_zz_dataOut_payload_0_16356 ? _zz_dataOut_payload_0_15986 : _zz_dataOut_payload_0_16013);
  assign _zz_dataOut_payload_128_114 = (_zz_dataOut_payload_0_16356 ? _zz_dataOut_payload_0_16013 : _zz_dataOut_payload_0_15986);
  assign _zz_dataOut_payload_0_16358 = (_zz_dataOut_payload_0_15987 < _zz_dataOut_payload_0_16012);
  assign _zz_dataOut_payload_0_16359 = (_zz_dataOut_payload_0_16358 ? _zz_dataOut_payload_0_15987 : _zz_dataOut_payload_0_16012);
  assign _zz_dataOut_payload_128_115 = (_zz_dataOut_payload_0_16358 ? _zz_dataOut_payload_0_16012 : _zz_dataOut_payload_0_15987);
  assign _zz_dataOut_payload_0_16360 = (_zz_dataOut_payload_0_15988 < _zz_dataOut_payload_0_16011);
  assign _zz_dataOut_payload_0_16361 = (_zz_dataOut_payload_0_16360 ? _zz_dataOut_payload_0_15988 : _zz_dataOut_payload_0_16011);
  assign _zz_dataOut_payload_128_116 = (_zz_dataOut_payload_0_16360 ? _zz_dataOut_payload_0_16011 : _zz_dataOut_payload_0_15988);
  assign _zz_dataOut_payload_0_16362 = (_zz_dataOut_payload_0_15989 < _zz_dataOut_payload_0_16010);
  assign _zz_dataOut_payload_0_16363 = (_zz_dataOut_payload_0_16362 ? _zz_dataOut_payload_0_15989 : _zz_dataOut_payload_0_16010);
  assign _zz_dataOut_payload_128_117 = (_zz_dataOut_payload_0_16362 ? _zz_dataOut_payload_0_16010 : _zz_dataOut_payload_0_15989);
  assign _zz_dataOut_payload_0_16364 = (_zz_dataOut_payload_0_15990 < _zz_dataOut_payload_0_16009);
  assign _zz_dataOut_payload_0_16365 = (_zz_dataOut_payload_0_16364 ? _zz_dataOut_payload_0_15990 : _zz_dataOut_payload_0_16009);
  assign _zz_dataOut_payload_128_118 = (_zz_dataOut_payload_0_16364 ? _zz_dataOut_payload_0_16009 : _zz_dataOut_payload_0_15990);
  assign _zz_dataOut_payload_0_16366 = (_zz_dataOut_payload_0_15991 < _zz_dataOut_payload_0_16008);
  assign _zz_dataOut_payload_0_16367 = (_zz_dataOut_payload_0_16366 ? _zz_dataOut_payload_0_15991 : _zz_dataOut_payload_0_16008);
  assign _zz_dataOut_payload_128_119 = (_zz_dataOut_payload_0_16366 ? _zz_dataOut_payload_0_16008 : _zz_dataOut_payload_0_15991);
  assign _zz_dataOut_payload_0_16368 = (_zz_dataOut_payload_0_15992 < _zz_dataOut_payload_0_16007);
  assign _zz_dataOut_payload_0_16369 = (_zz_dataOut_payload_0_16368 ? _zz_dataOut_payload_0_15992 : _zz_dataOut_payload_0_16007);
  assign _zz_dataOut_payload_128_120 = (_zz_dataOut_payload_0_16368 ? _zz_dataOut_payload_0_16007 : _zz_dataOut_payload_0_15992);
  assign _zz_dataOut_payload_0_16370 = (_zz_dataOut_payload_0_15993 < _zz_dataOut_payload_0_16006);
  assign _zz_dataOut_payload_0_16371 = (_zz_dataOut_payload_0_16370 ? _zz_dataOut_payload_0_15993 : _zz_dataOut_payload_0_16006);
  assign _zz_dataOut_payload_128_121 = (_zz_dataOut_payload_0_16370 ? _zz_dataOut_payload_0_16006 : _zz_dataOut_payload_0_15993);
  assign _zz_dataOut_payload_0_16372 = (_zz_dataOut_payload_0_15994 < _zz_dataOut_payload_0_16005);
  assign _zz_dataOut_payload_0_16373 = (_zz_dataOut_payload_0_16372 ? _zz_dataOut_payload_0_15994 : _zz_dataOut_payload_0_16005);
  assign _zz_dataOut_payload_128_122 = (_zz_dataOut_payload_0_16372 ? _zz_dataOut_payload_0_16005 : _zz_dataOut_payload_0_15994);
  assign _zz_dataOut_payload_0_16374 = (_zz_dataOut_payload_0_15995 < _zz_dataOut_payload_0_16004);
  assign _zz_dataOut_payload_0_16375 = (_zz_dataOut_payload_0_16374 ? _zz_dataOut_payload_0_15995 : _zz_dataOut_payload_0_16004);
  assign _zz_dataOut_payload_128_123 = (_zz_dataOut_payload_0_16374 ? _zz_dataOut_payload_0_16004 : _zz_dataOut_payload_0_15995);
  assign _zz_dataOut_payload_0_16376 = (_zz_dataOut_payload_0_15996 < _zz_dataOut_payload_0_16003);
  assign _zz_dataOut_payload_0_16377 = (_zz_dataOut_payload_0_16376 ? _zz_dataOut_payload_0_15996 : _zz_dataOut_payload_0_16003);
  assign _zz_dataOut_payload_128_124 = (_zz_dataOut_payload_0_16376 ? _zz_dataOut_payload_0_16003 : _zz_dataOut_payload_0_15996);
  assign _zz_dataOut_payload_0_16378 = (_zz_dataOut_payload_0_15997 < _zz_dataOut_payload_0_16002);
  assign _zz_dataOut_payload_0_16379 = (_zz_dataOut_payload_0_16378 ? _zz_dataOut_payload_0_15997 : _zz_dataOut_payload_0_16002);
  assign _zz_dataOut_payload_128_125 = (_zz_dataOut_payload_0_16378 ? _zz_dataOut_payload_0_16002 : _zz_dataOut_payload_0_15997);
  assign _zz_dataOut_payload_0_16380 = (_zz_dataOut_payload_0_15998 < _zz_dataOut_payload_0_16001);
  assign _zz_dataOut_payload_0_16381 = (_zz_dataOut_payload_0_16380 ? _zz_dataOut_payload_0_15998 : _zz_dataOut_payload_0_16001);
  assign _zz_dataOut_payload_128_126 = (_zz_dataOut_payload_0_16380 ? _zz_dataOut_payload_0_16001 : _zz_dataOut_payload_0_15998);
  assign _zz_dataOut_payload_0_16382 = (_zz_dataOut_payload_0_15999 < _zz_dataOut_payload_0_16000);
  assign _zz_dataOut_payload_0_16383 = (_zz_dataOut_payload_0_16382 ? _zz_dataOut_payload_0_15999 : _zz_dataOut_payload_0_16000);
  assign _zz_dataOut_payload_128_127 = (_zz_dataOut_payload_0_16382 ? _zz_dataOut_payload_0_16000 : _zz_dataOut_payload_0_15999);
  assign _zz_dataOut_payload_0_16384 = (_zz_dataOut_payload_0_16129 < _zz_dataOut_payload_0_16257);
  assign _zz_dataOut_payload_0_16385 = (_zz_dataOut_payload_0_16384 ? _zz_dataOut_payload_0_16129 : _zz_dataOut_payload_0_16257);
  assign _zz_dataOut_payload_64 = (_zz_dataOut_payload_0_16384 ? _zz_dataOut_payload_0_16257 : _zz_dataOut_payload_0_16129);
  assign _zz_dataOut_payload_0_16386 = (_zz_dataOut_payload_0_16131 < _zz_dataOut_payload_0_16259);
  assign _zz_dataOut_payload_0_16387 = (_zz_dataOut_payload_0_16386 ? _zz_dataOut_payload_0_16131 : _zz_dataOut_payload_0_16259);
  assign _zz_dataOut_payload_64_1 = (_zz_dataOut_payload_0_16386 ? _zz_dataOut_payload_0_16259 : _zz_dataOut_payload_0_16131);
  assign _zz_dataOut_payload_0_16388 = (_zz_dataOut_payload_0_16133 < _zz_dataOut_payload_0_16261);
  assign _zz_dataOut_payload_0_16389 = (_zz_dataOut_payload_0_16388 ? _zz_dataOut_payload_0_16133 : _zz_dataOut_payload_0_16261);
  assign _zz_dataOut_payload_64_2 = (_zz_dataOut_payload_0_16388 ? _zz_dataOut_payload_0_16261 : _zz_dataOut_payload_0_16133);
  assign _zz_dataOut_payload_0_16390 = (_zz_dataOut_payload_0_16135 < _zz_dataOut_payload_0_16263);
  assign _zz_dataOut_payload_0_16391 = (_zz_dataOut_payload_0_16390 ? _zz_dataOut_payload_0_16135 : _zz_dataOut_payload_0_16263);
  assign _zz_dataOut_payload_64_3 = (_zz_dataOut_payload_0_16390 ? _zz_dataOut_payload_0_16263 : _zz_dataOut_payload_0_16135);
  assign _zz_dataOut_payload_0_16392 = (_zz_dataOut_payload_0_16137 < _zz_dataOut_payload_0_16265);
  assign _zz_dataOut_payload_0_16393 = (_zz_dataOut_payload_0_16392 ? _zz_dataOut_payload_0_16137 : _zz_dataOut_payload_0_16265);
  assign _zz_dataOut_payload_64_4 = (_zz_dataOut_payload_0_16392 ? _zz_dataOut_payload_0_16265 : _zz_dataOut_payload_0_16137);
  assign _zz_dataOut_payload_0_16394 = (_zz_dataOut_payload_0_16139 < _zz_dataOut_payload_0_16267);
  assign _zz_dataOut_payload_0_16395 = (_zz_dataOut_payload_0_16394 ? _zz_dataOut_payload_0_16139 : _zz_dataOut_payload_0_16267);
  assign _zz_dataOut_payload_64_5 = (_zz_dataOut_payload_0_16394 ? _zz_dataOut_payload_0_16267 : _zz_dataOut_payload_0_16139);
  assign _zz_dataOut_payload_0_16396 = (_zz_dataOut_payload_0_16141 < _zz_dataOut_payload_0_16269);
  assign _zz_dataOut_payload_0_16397 = (_zz_dataOut_payload_0_16396 ? _zz_dataOut_payload_0_16141 : _zz_dataOut_payload_0_16269);
  assign _zz_dataOut_payload_64_6 = (_zz_dataOut_payload_0_16396 ? _zz_dataOut_payload_0_16269 : _zz_dataOut_payload_0_16141);
  assign _zz_dataOut_payload_0_16398 = (_zz_dataOut_payload_0_16143 < _zz_dataOut_payload_0_16271);
  assign _zz_dataOut_payload_0_16399 = (_zz_dataOut_payload_0_16398 ? _zz_dataOut_payload_0_16143 : _zz_dataOut_payload_0_16271);
  assign _zz_dataOut_payload_64_7 = (_zz_dataOut_payload_0_16398 ? _zz_dataOut_payload_0_16271 : _zz_dataOut_payload_0_16143);
  assign _zz_dataOut_payload_0_16400 = (_zz_dataOut_payload_0_16145 < _zz_dataOut_payload_0_16273);
  assign _zz_dataOut_payload_0_16401 = (_zz_dataOut_payload_0_16400 ? _zz_dataOut_payload_0_16145 : _zz_dataOut_payload_0_16273);
  assign _zz_dataOut_payload_64_8 = (_zz_dataOut_payload_0_16400 ? _zz_dataOut_payload_0_16273 : _zz_dataOut_payload_0_16145);
  assign _zz_dataOut_payload_0_16402 = (_zz_dataOut_payload_0_16147 < _zz_dataOut_payload_0_16275);
  assign _zz_dataOut_payload_0_16403 = (_zz_dataOut_payload_0_16402 ? _zz_dataOut_payload_0_16147 : _zz_dataOut_payload_0_16275);
  assign _zz_dataOut_payload_64_9 = (_zz_dataOut_payload_0_16402 ? _zz_dataOut_payload_0_16275 : _zz_dataOut_payload_0_16147);
  assign _zz_dataOut_payload_0_16404 = (_zz_dataOut_payload_0_16149 < _zz_dataOut_payload_0_16277);
  assign _zz_dataOut_payload_0_16405 = (_zz_dataOut_payload_0_16404 ? _zz_dataOut_payload_0_16149 : _zz_dataOut_payload_0_16277);
  assign _zz_dataOut_payload_64_10 = (_zz_dataOut_payload_0_16404 ? _zz_dataOut_payload_0_16277 : _zz_dataOut_payload_0_16149);
  assign _zz_dataOut_payload_0_16406 = (_zz_dataOut_payload_0_16151 < _zz_dataOut_payload_0_16279);
  assign _zz_dataOut_payload_0_16407 = (_zz_dataOut_payload_0_16406 ? _zz_dataOut_payload_0_16151 : _zz_dataOut_payload_0_16279);
  assign _zz_dataOut_payload_64_11 = (_zz_dataOut_payload_0_16406 ? _zz_dataOut_payload_0_16279 : _zz_dataOut_payload_0_16151);
  assign _zz_dataOut_payload_0_16408 = (_zz_dataOut_payload_0_16153 < _zz_dataOut_payload_0_16281);
  assign _zz_dataOut_payload_0_16409 = (_zz_dataOut_payload_0_16408 ? _zz_dataOut_payload_0_16153 : _zz_dataOut_payload_0_16281);
  assign _zz_dataOut_payload_64_12 = (_zz_dataOut_payload_0_16408 ? _zz_dataOut_payload_0_16281 : _zz_dataOut_payload_0_16153);
  assign _zz_dataOut_payload_0_16410 = (_zz_dataOut_payload_0_16155 < _zz_dataOut_payload_0_16283);
  assign _zz_dataOut_payload_0_16411 = (_zz_dataOut_payload_0_16410 ? _zz_dataOut_payload_0_16155 : _zz_dataOut_payload_0_16283);
  assign _zz_dataOut_payload_64_13 = (_zz_dataOut_payload_0_16410 ? _zz_dataOut_payload_0_16283 : _zz_dataOut_payload_0_16155);
  assign _zz_dataOut_payload_0_16412 = (_zz_dataOut_payload_0_16157 < _zz_dataOut_payload_0_16285);
  assign _zz_dataOut_payload_0_16413 = (_zz_dataOut_payload_0_16412 ? _zz_dataOut_payload_0_16157 : _zz_dataOut_payload_0_16285);
  assign _zz_dataOut_payload_64_14 = (_zz_dataOut_payload_0_16412 ? _zz_dataOut_payload_0_16285 : _zz_dataOut_payload_0_16157);
  assign _zz_dataOut_payload_0_16414 = (_zz_dataOut_payload_0_16159 < _zz_dataOut_payload_0_16287);
  assign _zz_dataOut_payload_0_16415 = (_zz_dataOut_payload_0_16414 ? _zz_dataOut_payload_0_16159 : _zz_dataOut_payload_0_16287);
  assign _zz_dataOut_payload_64_15 = (_zz_dataOut_payload_0_16414 ? _zz_dataOut_payload_0_16287 : _zz_dataOut_payload_0_16159);
  assign _zz_dataOut_payload_0_16416 = (_zz_dataOut_payload_0_16161 < _zz_dataOut_payload_0_16289);
  assign _zz_dataOut_payload_0_16417 = (_zz_dataOut_payload_0_16416 ? _zz_dataOut_payload_0_16161 : _zz_dataOut_payload_0_16289);
  assign _zz_dataOut_payload_64_16 = (_zz_dataOut_payload_0_16416 ? _zz_dataOut_payload_0_16289 : _zz_dataOut_payload_0_16161);
  assign _zz_dataOut_payload_0_16418 = (_zz_dataOut_payload_0_16163 < _zz_dataOut_payload_0_16291);
  assign _zz_dataOut_payload_0_16419 = (_zz_dataOut_payload_0_16418 ? _zz_dataOut_payload_0_16163 : _zz_dataOut_payload_0_16291);
  assign _zz_dataOut_payload_64_17 = (_zz_dataOut_payload_0_16418 ? _zz_dataOut_payload_0_16291 : _zz_dataOut_payload_0_16163);
  assign _zz_dataOut_payload_0_16420 = (_zz_dataOut_payload_0_16165 < _zz_dataOut_payload_0_16293);
  assign _zz_dataOut_payload_0_16421 = (_zz_dataOut_payload_0_16420 ? _zz_dataOut_payload_0_16165 : _zz_dataOut_payload_0_16293);
  assign _zz_dataOut_payload_64_18 = (_zz_dataOut_payload_0_16420 ? _zz_dataOut_payload_0_16293 : _zz_dataOut_payload_0_16165);
  assign _zz_dataOut_payload_0_16422 = (_zz_dataOut_payload_0_16167 < _zz_dataOut_payload_0_16295);
  assign _zz_dataOut_payload_0_16423 = (_zz_dataOut_payload_0_16422 ? _zz_dataOut_payload_0_16167 : _zz_dataOut_payload_0_16295);
  assign _zz_dataOut_payload_64_19 = (_zz_dataOut_payload_0_16422 ? _zz_dataOut_payload_0_16295 : _zz_dataOut_payload_0_16167);
  assign _zz_dataOut_payload_0_16424 = (_zz_dataOut_payload_0_16169 < _zz_dataOut_payload_0_16297);
  assign _zz_dataOut_payload_0_16425 = (_zz_dataOut_payload_0_16424 ? _zz_dataOut_payload_0_16169 : _zz_dataOut_payload_0_16297);
  assign _zz_dataOut_payload_64_20 = (_zz_dataOut_payload_0_16424 ? _zz_dataOut_payload_0_16297 : _zz_dataOut_payload_0_16169);
  assign _zz_dataOut_payload_0_16426 = (_zz_dataOut_payload_0_16171 < _zz_dataOut_payload_0_16299);
  assign _zz_dataOut_payload_0_16427 = (_zz_dataOut_payload_0_16426 ? _zz_dataOut_payload_0_16171 : _zz_dataOut_payload_0_16299);
  assign _zz_dataOut_payload_64_21 = (_zz_dataOut_payload_0_16426 ? _zz_dataOut_payload_0_16299 : _zz_dataOut_payload_0_16171);
  assign _zz_dataOut_payload_0_16428 = (_zz_dataOut_payload_0_16173 < _zz_dataOut_payload_0_16301);
  assign _zz_dataOut_payload_0_16429 = (_zz_dataOut_payload_0_16428 ? _zz_dataOut_payload_0_16173 : _zz_dataOut_payload_0_16301);
  assign _zz_dataOut_payload_64_22 = (_zz_dataOut_payload_0_16428 ? _zz_dataOut_payload_0_16301 : _zz_dataOut_payload_0_16173);
  assign _zz_dataOut_payload_0_16430 = (_zz_dataOut_payload_0_16175 < _zz_dataOut_payload_0_16303);
  assign _zz_dataOut_payload_0_16431 = (_zz_dataOut_payload_0_16430 ? _zz_dataOut_payload_0_16175 : _zz_dataOut_payload_0_16303);
  assign _zz_dataOut_payload_64_23 = (_zz_dataOut_payload_0_16430 ? _zz_dataOut_payload_0_16303 : _zz_dataOut_payload_0_16175);
  assign _zz_dataOut_payload_0_16432 = (_zz_dataOut_payload_0_16177 < _zz_dataOut_payload_0_16305);
  assign _zz_dataOut_payload_0_16433 = (_zz_dataOut_payload_0_16432 ? _zz_dataOut_payload_0_16177 : _zz_dataOut_payload_0_16305);
  assign _zz_dataOut_payload_64_24 = (_zz_dataOut_payload_0_16432 ? _zz_dataOut_payload_0_16305 : _zz_dataOut_payload_0_16177);
  assign _zz_dataOut_payload_0_16434 = (_zz_dataOut_payload_0_16179 < _zz_dataOut_payload_0_16307);
  assign _zz_dataOut_payload_0_16435 = (_zz_dataOut_payload_0_16434 ? _zz_dataOut_payload_0_16179 : _zz_dataOut_payload_0_16307);
  assign _zz_dataOut_payload_64_25 = (_zz_dataOut_payload_0_16434 ? _zz_dataOut_payload_0_16307 : _zz_dataOut_payload_0_16179);
  assign _zz_dataOut_payload_0_16436 = (_zz_dataOut_payload_0_16181 < _zz_dataOut_payload_0_16309);
  assign _zz_dataOut_payload_0_16437 = (_zz_dataOut_payload_0_16436 ? _zz_dataOut_payload_0_16181 : _zz_dataOut_payload_0_16309);
  assign _zz_dataOut_payload_64_26 = (_zz_dataOut_payload_0_16436 ? _zz_dataOut_payload_0_16309 : _zz_dataOut_payload_0_16181);
  assign _zz_dataOut_payload_0_16438 = (_zz_dataOut_payload_0_16183 < _zz_dataOut_payload_0_16311);
  assign _zz_dataOut_payload_0_16439 = (_zz_dataOut_payload_0_16438 ? _zz_dataOut_payload_0_16183 : _zz_dataOut_payload_0_16311);
  assign _zz_dataOut_payload_64_27 = (_zz_dataOut_payload_0_16438 ? _zz_dataOut_payload_0_16311 : _zz_dataOut_payload_0_16183);
  assign _zz_dataOut_payload_0_16440 = (_zz_dataOut_payload_0_16185 < _zz_dataOut_payload_0_16313);
  assign _zz_dataOut_payload_0_16441 = (_zz_dataOut_payload_0_16440 ? _zz_dataOut_payload_0_16185 : _zz_dataOut_payload_0_16313);
  assign _zz_dataOut_payload_64_28 = (_zz_dataOut_payload_0_16440 ? _zz_dataOut_payload_0_16313 : _zz_dataOut_payload_0_16185);
  assign _zz_dataOut_payload_0_16442 = (_zz_dataOut_payload_0_16187 < _zz_dataOut_payload_0_16315);
  assign _zz_dataOut_payload_0_16443 = (_zz_dataOut_payload_0_16442 ? _zz_dataOut_payload_0_16187 : _zz_dataOut_payload_0_16315);
  assign _zz_dataOut_payload_64_29 = (_zz_dataOut_payload_0_16442 ? _zz_dataOut_payload_0_16315 : _zz_dataOut_payload_0_16187);
  assign _zz_dataOut_payload_0_16444 = (_zz_dataOut_payload_0_16189 < _zz_dataOut_payload_0_16317);
  assign _zz_dataOut_payload_0_16445 = (_zz_dataOut_payload_0_16444 ? _zz_dataOut_payload_0_16189 : _zz_dataOut_payload_0_16317);
  assign _zz_dataOut_payload_64_30 = (_zz_dataOut_payload_0_16444 ? _zz_dataOut_payload_0_16317 : _zz_dataOut_payload_0_16189);
  assign _zz_dataOut_payload_0_16446 = (_zz_dataOut_payload_0_16191 < _zz_dataOut_payload_0_16319);
  assign _zz_dataOut_payload_0_16447 = (_zz_dataOut_payload_0_16446 ? _zz_dataOut_payload_0_16191 : _zz_dataOut_payload_0_16319);
  assign _zz_dataOut_payload_64_31 = (_zz_dataOut_payload_0_16446 ? _zz_dataOut_payload_0_16319 : _zz_dataOut_payload_0_16191);
  assign _zz_dataOut_payload_0_16448 = (_zz_dataOut_payload_0_16193 < _zz_dataOut_payload_0_16321);
  assign _zz_dataOut_payload_0_16449 = (_zz_dataOut_payload_0_16448 ? _zz_dataOut_payload_0_16193 : _zz_dataOut_payload_0_16321);
  assign _zz_dataOut_payload_64_32 = (_zz_dataOut_payload_0_16448 ? _zz_dataOut_payload_0_16321 : _zz_dataOut_payload_0_16193);
  assign _zz_dataOut_payload_0_16450 = (_zz_dataOut_payload_0_16195 < _zz_dataOut_payload_0_16323);
  assign _zz_dataOut_payload_0_16451 = (_zz_dataOut_payload_0_16450 ? _zz_dataOut_payload_0_16195 : _zz_dataOut_payload_0_16323);
  assign _zz_dataOut_payload_64_33 = (_zz_dataOut_payload_0_16450 ? _zz_dataOut_payload_0_16323 : _zz_dataOut_payload_0_16195);
  assign _zz_dataOut_payload_0_16452 = (_zz_dataOut_payload_0_16197 < _zz_dataOut_payload_0_16325);
  assign _zz_dataOut_payload_0_16453 = (_zz_dataOut_payload_0_16452 ? _zz_dataOut_payload_0_16197 : _zz_dataOut_payload_0_16325);
  assign _zz_dataOut_payload_64_34 = (_zz_dataOut_payload_0_16452 ? _zz_dataOut_payload_0_16325 : _zz_dataOut_payload_0_16197);
  assign _zz_dataOut_payload_0_16454 = (_zz_dataOut_payload_0_16199 < _zz_dataOut_payload_0_16327);
  assign _zz_dataOut_payload_0_16455 = (_zz_dataOut_payload_0_16454 ? _zz_dataOut_payload_0_16199 : _zz_dataOut_payload_0_16327);
  assign _zz_dataOut_payload_64_35 = (_zz_dataOut_payload_0_16454 ? _zz_dataOut_payload_0_16327 : _zz_dataOut_payload_0_16199);
  assign _zz_dataOut_payload_0_16456 = (_zz_dataOut_payload_0_16201 < _zz_dataOut_payload_0_16329);
  assign _zz_dataOut_payload_0_16457 = (_zz_dataOut_payload_0_16456 ? _zz_dataOut_payload_0_16201 : _zz_dataOut_payload_0_16329);
  assign _zz_dataOut_payload_64_36 = (_zz_dataOut_payload_0_16456 ? _zz_dataOut_payload_0_16329 : _zz_dataOut_payload_0_16201);
  assign _zz_dataOut_payload_0_16458 = (_zz_dataOut_payload_0_16203 < _zz_dataOut_payload_0_16331);
  assign _zz_dataOut_payload_0_16459 = (_zz_dataOut_payload_0_16458 ? _zz_dataOut_payload_0_16203 : _zz_dataOut_payload_0_16331);
  assign _zz_dataOut_payload_64_37 = (_zz_dataOut_payload_0_16458 ? _zz_dataOut_payload_0_16331 : _zz_dataOut_payload_0_16203);
  assign _zz_dataOut_payload_0_16460 = (_zz_dataOut_payload_0_16205 < _zz_dataOut_payload_0_16333);
  assign _zz_dataOut_payload_0_16461 = (_zz_dataOut_payload_0_16460 ? _zz_dataOut_payload_0_16205 : _zz_dataOut_payload_0_16333);
  assign _zz_dataOut_payload_64_38 = (_zz_dataOut_payload_0_16460 ? _zz_dataOut_payload_0_16333 : _zz_dataOut_payload_0_16205);
  assign _zz_dataOut_payload_0_16462 = (_zz_dataOut_payload_0_16207 < _zz_dataOut_payload_0_16335);
  assign _zz_dataOut_payload_0_16463 = (_zz_dataOut_payload_0_16462 ? _zz_dataOut_payload_0_16207 : _zz_dataOut_payload_0_16335);
  assign _zz_dataOut_payload_64_39 = (_zz_dataOut_payload_0_16462 ? _zz_dataOut_payload_0_16335 : _zz_dataOut_payload_0_16207);
  assign _zz_dataOut_payload_0_16464 = (_zz_dataOut_payload_0_16209 < _zz_dataOut_payload_0_16337);
  assign _zz_dataOut_payload_0_16465 = (_zz_dataOut_payload_0_16464 ? _zz_dataOut_payload_0_16209 : _zz_dataOut_payload_0_16337);
  assign _zz_dataOut_payload_64_40 = (_zz_dataOut_payload_0_16464 ? _zz_dataOut_payload_0_16337 : _zz_dataOut_payload_0_16209);
  assign _zz_dataOut_payload_0_16466 = (_zz_dataOut_payload_0_16211 < _zz_dataOut_payload_0_16339);
  assign _zz_dataOut_payload_0_16467 = (_zz_dataOut_payload_0_16466 ? _zz_dataOut_payload_0_16211 : _zz_dataOut_payload_0_16339);
  assign _zz_dataOut_payload_64_41 = (_zz_dataOut_payload_0_16466 ? _zz_dataOut_payload_0_16339 : _zz_dataOut_payload_0_16211);
  assign _zz_dataOut_payload_0_16468 = (_zz_dataOut_payload_0_16213 < _zz_dataOut_payload_0_16341);
  assign _zz_dataOut_payload_0_16469 = (_zz_dataOut_payload_0_16468 ? _zz_dataOut_payload_0_16213 : _zz_dataOut_payload_0_16341);
  assign _zz_dataOut_payload_64_42 = (_zz_dataOut_payload_0_16468 ? _zz_dataOut_payload_0_16341 : _zz_dataOut_payload_0_16213);
  assign _zz_dataOut_payload_0_16470 = (_zz_dataOut_payload_0_16215 < _zz_dataOut_payload_0_16343);
  assign _zz_dataOut_payload_0_16471 = (_zz_dataOut_payload_0_16470 ? _zz_dataOut_payload_0_16215 : _zz_dataOut_payload_0_16343);
  assign _zz_dataOut_payload_64_43 = (_zz_dataOut_payload_0_16470 ? _zz_dataOut_payload_0_16343 : _zz_dataOut_payload_0_16215);
  assign _zz_dataOut_payload_0_16472 = (_zz_dataOut_payload_0_16217 < _zz_dataOut_payload_0_16345);
  assign _zz_dataOut_payload_0_16473 = (_zz_dataOut_payload_0_16472 ? _zz_dataOut_payload_0_16217 : _zz_dataOut_payload_0_16345);
  assign _zz_dataOut_payload_64_44 = (_zz_dataOut_payload_0_16472 ? _zz_dataOut_payload_0_16345 : _zz_dataOut_payload_0_16217);
  assign _zz_dataOut_payload_0_16474 = (_zz_dataOut_payload_0_16219 < _zz_dataOut_payload_0_16347);
  assign _zz_dataOut_payload_0_16475 = (_zz_dataOut_payload_0_16474 ? _zz_dataOut_payload_0_16219 : _zz_dataOut_payload_0_16347);
  assign _zz_dataOut_payload_64_45 = (_zz_dataOut_payload_0_16474 ? _zz_dataOut_payload_0_16347 : _zz_dataOut_payload_0_16219);
  assign _zz_dataOut_payload_0_16476 = (_zz_dataOut_payload_0_16221 < _zz_dataOut_payload_0_16349);
  assign _zz_dataOut_payload_0_16477 = (_zz_dataOut_payload_0_16476 ? _zz_dataOut_payload_0_16221 : _zz_dataOut_payload_0_16349);
  assign _zz_dataOut_payload_64_46 = (_zz_dataOut_payload_0_16476 ? _zz_dataOut_payload_0_16349 : _zz_dataOut_payload_0_16221);
  assign _zz_dataOut_payload_0_16478 = (_zz_dataOut_payload_0_16223 < _zz_dataOut_payload_0_16351);
  assign _zz_dataOut_payload_0_16479 = (_zz_dataOut_payload_0_16478 ? _zz_dataOut_payload_0_16223 : _zz_dataOut_payload_0_16351);
  assign _zz_dataOut_payload_64_47 = (_zz_dataOut_payload_0_16478 ? _zz_dataOut_payload_0_16351 : _zz_dataOut_payload_0_16223);
  assign _zz_dataOut_payload_0_16480 = (_zz_dataOut_payload_0_16225 < _zz_dataOut_payload_0_16353);
  assign _zz_dataOut_payload_0_16481 = (_zz_dataOut_payload_0_16480 ? _zz_dataOut_payload_0_16225 : _zz_dataOut_payload_0_16353);
  assign _zz_dataOut_payload_64_48 = (_zz_dataOut_payload_0_16480 ? _zz_dataOut_payload_0_16353 : _zz_dataOut_payload_0_16225);
  assign _zz_dataOut_payload_0_16482 = (_zz_dataOut_payload_0_16227 < _zz_dataOut_payload_0_16355);
  assign _zz_dataOut_payload_0_16483 = (_zz_dataOut_payload_0_16482 ? _zz_dataOut_payload_0_16227 : _zz_dataOut_payload_0_16355);
  assign _zz_dataOut_payload_64_49 = (_zz_dataOut_payload_0_16482 ? _zz_dataOut_payload_0_16355 : _zz_dataOut_payload_0_16227);
  assign _zz_dataOut_payload_0_16484 = (_zz_dataOut_payload_0_16229 < _zz_dataOut_payload_0_16357);
  assign _zz_dataOut_payload_0_16485 = (_zz_dataOut_payload_0_16484 ? _zz_dataOut_payload_0_16229 : _zz_dataOut_payload_0_16357);
  assign _zz_dataOut_payload_64_50 = (_zz_dataOut_payload_0_16484 ? _zz_dataOut_payload_0_16357 : _zz_dataOut_payload_0_16229);
  assign _zz_dataOut_payload_0_16486 = (_zz_dataOut_payload_0_16231 < _zz_dataOut_payload_0_16359);
  assign _zz_dataOut_payload_0_16487 = (_zz_dataOut_payload_0_16486 ? _zz_dataOut_payload_0_16231 : _zz_dataOut_payload_0_16359);
  assign _zz_dataOut_payload_64_51 = (_zz_dataOut_payload_0_16486 ? _zz_dataOut_payload_0_16359 : _zz_dataOut_payload_0_16231);
  assign _zz_dataOut_payload_0_16488 = (_zz_dataOut_payload_0_16233 < _zz_dataOut_payload_0_16361);
  assign _zz_dataOut_payload_0_16489 = (_zz_dataOut_payload_0_16488 ? _zz_dataOut_payload_0_16233 : _zz_dataOut_payload_0_16361);
  assign _zz_dataOut_payload_64_52 = (_zz_dataOut_payload_0_16488 ? _zz_dataOut_payload_0_16361 : _zz_dataOut_payload_0_16233);
  assign _zz_dataOut_payload_0_16490 = (_zz_dataOut_payload_0_16235 < _zz_dataOut_payload_0_16363);
  assign _zz_dataOut_payload_0_16491 = (_zz_dataOut_payload_0_16490 ? _zz_dataOut_payload_0_16235 : _zz_dataOut_payload_0_16363);
  assign _zz_dataOut_payload_64_53 = (_zz_dataOut_payload_0_16490 ? _zz_dataOut_payload_0_16363 : _zz_dataOut_payload_0_16235);
  assign _zz_dataOut_payload_0_16492 = (_zz_dataOut_payload_0_16237 < _zz_dataOut_payload_0_16365);
  assign _zz_dataOut_payload_0_16493 = (_zz_dataOut_payload_0_16492 ? _zz_dataOut_payload_0_16237 : _zz_dataOut_payload_0_16365);
  assign _zz_dataOut_payload_64_54 = (_zz_dataOut_payload_0_16492 ? _zz_dataOut_payload_0_16365 : _zz_dataOut_payload_0_16237);
  assign _zz_dataOut_payload_0_16494 = (_zz_dataOut_payload_0_16239 < _zz_dataOut_payload_0_16367);
  assign _zz_dataOut_payload_0_16495 = (_zz_dataOut_payload_0_16494 ? _zz_dataOut_payload_0_16239 : _zz_dataOut_payload_0_16367);
  assign _zz_dataOut_payload_64_55 = (_zz_dataOut_payload_0_16494 ? _zz_dataOut_payload_0_16367 : _zz_dataOut_payload_0_16239);
  assign _zz_dataOut_payload_0_16496 = (_zz_dataOut_payload_0_16241 < _zz_dataOut_payload_0_16369);
  assign _zz_dataOut_payload_0_16497 = (_zz_dataOut_payload_0_16496 ? _zz_dataOut_payload_0_16241 : _zz_dataOut_payload_0_16369);
  assign _zz_dataOut_payload_64_56 = (_zz_dataOut_payload_0_16496 ? _zz_dataOut_payload_0_16369 : _zz_dataOut_payload_0_16241);
  assign _zz_dataOut_payload_0_16498 = (_zz_dataOut_payload_0_16243 < _zz_dataOut_payload_0_16371);
  assign _zz_dataOut_payload_0_16499 = (_zz_dataOut_payload_0_16498 ? _zz_dataOut_payload_0_16243 : _zz_dataOut_payload_0_16371);
  assign _zz_dataOut_payload_64_57 = (_zz_dataOut_payload_0_16498 ? _zz_dataOut_payload_0_16371 : _zz_dataOut_payload_0_16243);
  assign _zz_dataOut_payload_0_16500 = (_zz_dataOut_payload_0_16245 < _zz_dataOut_payload_0_16373);
  assign _zz_dataOut_payload_0_16501 = (_zz_dataOut_payload_0_16500 ? _zz_dataOut_payload_0_16245 : _zz_dataOut_payload_0_16373);
  assign _zz_dataOut_payload_64_58 = (_zz_dataOut_payload_0_16500 ? _zz_dataOut_payload_0_16373 : _zz_dataOut_payload_0_16245);
  assign _zz_dataOut_payload_0_16502 = (_zz_dataOut_payload_0_16247 < _zz_dataOut_payload_0_16375);
  assign _zz_dataOut_payload_0_16503 = (_zz_dataOut_payload_0_16502 ? _zz_dataOut_payload_0_16247 : _zz_dataOut_payload_0_16375);
  assign _zz_dataOut_payload_64_59 = (_zz_dataOut_payload_0_16502 ? _zz_dataOut_payload_0_16375 : _zz_dataOut_payload_0_16247);
  assign _zz_dataOut_payload_0_16504 = (_zz_dataOut_payload_0_16249 < _zz_dataOut_payload_0_16377);
  assign _zz_dataOut_payload_0_16505 = (_zz_dataOut_payload_0_16504 ? _zz_dataOut_payload_0_16249 : _zz_dataOut_payload_0_16377);
  assign _zz_dataOut_payload_64_60 = (_zz_dataOut_payload_0_16504 ? _zz_dataOut_payload_0_16377 : _zz_dataOut_payload_0_16249);
  assign _zz_dataOut_payload_0_16506 = (_zz_dataOut_payload_0_16251 < _zz_dataOut_payload_0_16379);
  assign _zz_dataOut_payload_0_16507 = (_zz_dataOut_payload_0_16506 ? _zz_dataOut_payload_0_16251 : _zz_dataOut_payload_0_16379);
  assign _zz_dataOut_payload_64_61 = (_zz_dataOut_payload_0_16506 ? _zz_dataOut_payload_0_16379 : _zz_dataOut_payload_0_16251);
  assign _zz_dataOut_payload_0_16508 = (_zz_dataOut_payload_0_16253 < _zz_dataOut_payload_0_16381);
  assign _zz_dataOut_payload_0_16509 = (_zz_dataOut_payload_0_16508 ? _zz_dataOut_payload_0_16253 : _zz_dataOut_payload_0_16381);
  assign _zz_dataOut_payload_64_62 = (_zz_dataOut_payload_0_16508 ? _zz_dataOut_payload_0_16381 : _zz_dataOut_payload_0_16253);
  assign _zz_dataOut_payload_0_16510 = (_zz_dataOut_payload_0_16255 < _zz_dataOut_payload_0_16383);
  assign _zz_dataOut_payload_0_16511 = (_zz_dataOut_payload_0_16510 ? _zz_dataOut_payload_0_16255 : _zz_dataOut_payload_0_16383);
  assign _zz_dataOut_payload_64_63 = (_zz_dataOut_payload_0_16510 ? _zz_dataOut_payload_0_16383 : _zz_dataOut_payload_0_16255);
  assign _zz_dataOut_payload_0_16512 = (_zz_dataOut_payload_0_16385 < _zz_dataOut_payload_0_16449);
  assign _zz_dataOut_payload_0_16513 = (_zz_dataOut_payload_0_16512 ? _zz_dataOut_payload_0_16385 : _zz_dataOut_payload_0_16449);
  assign _zz_dataOut_payload_32 = (_zz_dataOut_payload_0_16512 ? _zz_dataOut_payload_0_16449 : _zz_dataOut_payload_0_16385);
  assign _zz_dataOut_payload_0_16514 = (_zz_dataOut_payload_0_16387 < _zz_dataOut_payload_0_16451);
  assign _zz_dataOut_payload_0_16515 = (_zz_dataOut_payload_0_16514 ? _zz_dataOut_payload_0_16387 : _zz_dataOut_payload_0_16451);
  assign _zz_dataOut_payload_32_1 = (_zz_dataOut_payload_0_16514 ? _zz_dataOut_payload_0_16451 : _zz_dataOut_payload_0_16387);
  assign _zz_dataOut_payload_0_16516 = (_zz_dataOut_payload_0_16389 < _zz_dataOut_payload_0_16453);
  assign _zz_dataOut_payload_0_16517 = (_zz_dataOut_payload_0_16516 ? _zz_dataOut_payload_0_16389 : _zz_dataOut_payload_0_16453);
  assign _zz_dataOut_payload_32_2 = (_zz_dataOut_payload_0_16516 ? _zz_dataOut_payload_0_16453 : _zz_dataOut_payload_0_16389);
  assign _zz_dataOut_payload_0_16518 = (_zz_dataOut_payload_0_16391 < _zz_dataOut_payload_0_16455);
  assign _zz_dataOut_payload_0_16519 = (_zz_dataOut_payload_0_16518 ? _zz_dataOut_payload_0_16391 : _zz_dataOut_payload_0_16455);
  assign _zz_dataOut_payload_32_3 = (_zz_dataOut_payload_0_16518 ? _zz_dataOut_payload_0_16455 : _zz_dataOut_payload_0_16391);
  assign _zz_dataOut_payload_0_16520 = (_zz_dataOut_payload_0_16393 < _zz_dataOut_payload_0_16457);
  assign _zz_dataOut_payload_0_16521 = (_zz_dataOut_payload_0_16520 ? _zz_dataOut_payload_0_16393 : _zz_dataOut_payload_0_16457);
  assign _zz_dataOut_payload_32_4 = (_zz_dataOut_payload_0_16520 ? _zz_dataOut_payload_0_16457 : _zz_dataOut_payload_0_16393);
  assign _zz_dataOut_payload_0_16522 = (_zz_dataOut_payload_0_16395 < _zz_dataOut_payload_0_16459);
  assign _zz_dataOut_payload_0_16523 = (_zz_dataOut_payload_0_16522 ? _zz_dataOut_payload_0_16395 : _zz_dataOut_payload_0_16459);
  assign _zz_dataOut_payload_32_5 = (_zz_dataOut_payload_0_16522 ? _zz_dataOut_payload_0_16459 : _zz_dataOut_payload_0_16395);
  assign _zz_dataOut_payload_0_16524 = (_zz_dataOut_payload_0_16397 < _zz_dataOut_payload_0_16461);
  assign _zz_dataOut_payload_0_16525 = (_zz_dataOut_payload_0_16524 ? _zz_dataOut_payload_0_16397 : _zz_dataOut_payload_0_16461);
  assign _zz_dataOut_payload_32_6 = (_zz_dataOut_payload_0_16524 ? _zz_dataOut_payload_0_16461 : _zz_dataOut_payload_0_16397);
  assign _zz_dataOut_payload_0_16526 = (_zz_dataOut_payload_0_16399 < _zz_dataOut_payload_0_16463);
  assign _zz_dataOut_payload_0_16527 = (_zz_dataOut_payload_0_16526 ? _zz_dataOut_payload_0_16399 : _zz_dataOut_payload_0_16463);
  assign _zz_dataOut_payload_32_7 = (_zz_dataOut_payload_0_16526 ? _zz_dataOut_payload_0_16463 : _zz_dataOut_payload_0_16399);
  assign _zz_dataOut_payload_0_16528 = (_zz_dataOut_payload_0_16401 < _zz_dataOut_payload_0_16465);
  assign _zz_dataOut_payload_0_16529 = (_zz_dataOut_payload_0_16528 ? _zz_dataOut_payload_0_16401 : _zz_dataOut_payload_0_16465);
  assign _zz_dataOut_payload_32_8 = (_zz_dataOut_payload_0_16528 ? _zz_dataOut_payload_0_16465 : _zz_dataOut_payload_0_16401);
  assign _zz_dataOut_payload_0_16530 = (_zz_dataOut_payload_0_16403 < _zz_dataOut_payload_0_16467);
  assign _zz_dataOut_payload_0_16531 = (_zz_dataOut_payload_0_16530 ? _zz_dataOut_payload_0_16403 : _zz_dataOut_payload_0_16467);
  assign _zz_dataOut_payload_32_9 = (_zz_dataOut_payload_0_16530 ? _zz_dataOut_payload_0_16467 : _zz_dataOut_payload_0_16403);
  assign _zz_dataOut_payload_0_16532 = (_zz_dataOut_payload_0_16405 < _zz_dataOut_payload_0_16469);
  assign _zz_dataOut_payload_0_16533 = (_zz_dataOut_payload_0_16532 ? _zz_dataOut_payload_0_16405 : _zz_dataOut_payload_0_16469);
  assign _zz_dataOut_payload_32_10 = (_zz_dataOut_payload_0_16532 ? _zz_dataOut_payload_0_16469 : _zz_dataOut_payload_0_16405);
  assign _zz_dataOut_payload_0_16534 = (_zz_dataOut_payload_0_16407 < _zz_dataOut_payload_0_16471);
  assign _zz_dataOut_payload_0_16535 = (_zz_dataOut_payload_0_16534 ? _zz_dataOut_payload_0_16407 : _zz_dataOut_payload_0_16471);
  assign _zz_dataOut_payload_32_11 = (_zz_dataOut_payload_0_16534 ? _zz_dataOut_payload_0_16471 : _zz_dataOut_payload_0_16407);
  assign _zz_dataOut_payload_0_16536 = (_zz_dataOut_payload_0_16409 < _zz_dataOut_payload_0_16473);
  assign _zz_dataOut_payload_0_16537 = (_zz_dataOut_payload_0_16536 ? _zz_dataOut_payload_0_16409 : _zz_dataOut_payload_0_16473);
  assign _zz_dataOut_payload_32_12 = (_zz_dataOut_payload_0_16536 ? _zz_dataOut_payload_0_16473 : _zz_dataOut_payload_0_16409);
  assign _zz_dataOut_payload_0_16538 = (_zz_dataOut_payload_0_16411 < _zz_dataOut_payload_0_16475);
  assign _zz_dataOut_payload_0_16539 = (_zz_dataOut_payload_0_16538 ? _zz_dataOut_payload_0_16411 : _zz_dataOut_payload_0_16475);
  assign _zz_dataOut_payload_32_13 = (_zz_dataOut_payload_0_16538 ? _zz_dataOut_payload_0_16475 : _zz_dataOut_payload_0_16411);
  assign _zz_dataOut_payload_0_16540 = (_zz_dataOut_payload_0_16413 < _zz_dataOut_payload_0_16477);
  assign _zz_dataOut_payload_0_16541 = (_zz_dataOut_payload_0_16540 ? _zz_dataOut_payload_0_16413 : _zz_dataOut_payload_0_16477);
  assign _zz_dataOut_payload_32_14 = (_zz_dataOut_payload_0_16540 ? _zz_dataOut_payload_0_16477 : _zz_dataOut_payload_0_16413);
  assign _zz_dataOut_payload_0_16542 = (_zz_dataOut_payload_0_16415 < _zz_dataOut_payload_0_16479);
  assign _zz_dataOut_payload_0_16543 = (_zz_dataOut_payload_0_16542 ? _zz_dataOut_payload_0_16415 : _zz_dataOut_payload_0_16479);
  assign _zz_dataOut_payload_32_15 = (_zz_dataOut_payload_0_16542 ? _zz_dataOut_payload_0_16479 : _zz_dataOut_payload_0_16415);
  assign _zz_dataOut_payload_0_16544 = (_zz_dataOut_payload_0_16417 < _zz_dataOut_payload_0_16481);
  assign _zz_dataOut_payload_0_16545 = (_zz_dataOut_payload_0_16544 ? _zz_dataOut_payload_0_16417 : _zz_dataOut_payload_0_16481);
  assign _zz_dataOut_payload_32_16 = (_zz_dataOut_payload_0_16544 ? _zz_dataOut_payload_0_16481 : _zz_dataOut_payload_0_16417);
  assign _zz_dataOut_payload_0_16546 = (_zz_dataOut_payload_0_16419 < _zz_dataOut_payload_0_16483);
  assign _zz_dataOut_payload_0_16547 = (_zz_dataOut_payload_0_16546 ? _zz_dataOut_payload_0_16419 : _zz_dataOut_payload_0_16483);
  assign _zz_dataOut_payload_32_17 = (_zz_dataOut_payload_0_16546 ? _zz_dataOut_payload_0_16483 : _zz_dataOut_payload_0_16419);
  assign _zz_dataOut_payload_0_16548 = (_zz_dataOut_payload_0_16421 < _zz_dataOut_payload_0_16485);
  assign _zz_dataOut_payload_0_16549 = (_zz_dataOut_payload_0_16548 ? _zz_dataOut_payload_0_16421 : _zz_dataOut_payload_0_16485);
  assign _zz_dataOut_payload_32_18 = (_zz_dataOut_payload_0_16548 ? _zz_dataOut_payload_0_16485 : _zz_dataOut_payload_0_16421);
  assign _zz_dataOut_payload_0_16550 = (_zz_dataOut_payload_0_16423 < _zz_dataOut_payload_0_16487);
  assign _zz_dataOut_payload_0_16551 = (_zz_dataOut_payload_0_16550 ? _zz_dataOut_payload_0_16423 : _zz_dataOut_payload_0_16487);
  assign _zz_dataOut_payload_32_19 = (_zz_dataOut_payload_0_16550 ? _zz_dataOut_payload_0_16487 : _zz_dataOut_payload_0_16423);
  assign _zz_dataOut_payload_0_16552 = (_zz_dataOut_payload_0_16425 < _zz_dataOut_payload_0_16489);
  assign _zz_dataOut_payload_0_16553 = (_zz_dataOut_payload_0_16552 ? _zz_dataOut_payload_0_16425 : _zz_dataOut_payload_0_16489);
  assign _zz_dataOut_payload_32_20 = (_zz_dataOut_payload_0_16552 ? _zz_dataOut_payload_0_16489 : _zz_dataOut_payload_0_16425);
  assign _zz_dataOut_payload_0_16554 = (_zz_dataOut_payload_0_16427 < _zz_dataOut_payload_0_16491);
  assign _zz_dataOut_payload_0_16555 = (_zz_dataOut_payload_0_16554 ? _zz_dataOut_payload_0_16427 : _zz_dataOut_payload_0_16491);
  assign _zz_dataOut_payload_32_21 = (_zz_dataOut_payload_0_16554 ? _zz_dataOut_payload_0_16491 : _zz_dataOut_payload_0_16427);
  assign _zz_dataOut_payload_0_16556 = (_zz_dataOut_payload_0_16429 < _zz_dataOut_payload_0_16493);
  assign _zz_dataOut_payload_0_16557 = (_zz_dataOut_payload_0_16556 ? _zz_dataOut_payload_0_16429 : _zz_dataOut_payload_0_16493);
  assign _zz_dataOut_payload_32_22 = (_zz_dataOut_payload_0_16556 ? _zz_dataOut_payload_0_16493 : _zz_dataOut_payload_0_16429);
  assign _zz_dataOut_payload_0_16558 = (_zz_dataOut_payload_0_16431 < _zz_dataOut_payload_0_16495);
  assign _zz_dataOut_payload_0_16559 = (_zz_dataOut_payload_0_16558 ? _zz_dataOut_payload_0_16431 : _zz_dataOut_payload_0_16495);
  assign _zz_dataOut_payload_32_23 = (_zz_dataOut_payload_0_16558 ? _zz_dataOut_payload_0_16495 : _zz_dataOut_payload_0_16431);
  assign _zz_dataOut_payload_0_16560 = (_zz_dataOut_payload_0_16433 < _zz_dataOut_payload_0_16497);
  assign _zz_dataOut_payload_0_16561 = (_zz_dataOut_payload_0_16560 ? _zz_dataOut_payload_0_16433 : _zz_dataOut_payload_0_16497);
  assign _zz_dataOut_payload_32_24 = (_zz_dataOut_payload_0_16560 ? _zz_dataOut_payload_0_16497 : _zz_dataOut_payload_0_16433);
  assign _zz_dataOut_payload_0_16562 = (_zz_dataOut_payload_0_16435 < _zz_dataOut_payload_0_16499);
  assign _zz_dataOut_payload_0_16563 = (_zz_dataOut_payload_0_16562 ? _zz_dataOut_payload_0_16435 : _zz_dataOut_payload_0_16499);
  assign _zz_dataOut_payload_32_25 = (_zz_dataOut_payload_0_16562 ? _zz_dataOut_payload_0_16499 : _zz_dataOut_payload_0_16435);
  assign _zz_dataOut_payload_0_16564 = (_zz_dataOut_payload_0_16437 < _zz_dataOut_payload_0_16501);
  assign _zz_dataOut_payload_0_16565 = (_zz_dataOut_payload_0_16564 ? _zz_dataOut_payload_0_16437 : _zz_dataOut_payload_0_16501);
  assign _zz_dataOut_payload_32_26 = (_zz_dataOut_payload_0_16564 ? _zz_dataOut_payload_0_16501 : _zz_dataOut_payload_0_16437);
  assign _zz_dataOut_payload_0_16566 = (_zz_dataOut_payload_0_16439 < _zz_dataOut_payload_0_16503);
  assign _zz_dataOut_payload_0_16567 = (_zz_dataOut_payload_0_16566 ? _zz_dataOut_payload_0_16439 : _zz_dataOut_payload_0_16503);
  assign _zz_dataOut_payload_32_27 = (_zz_dataOut_payload_0_16566 ? _zz_dataOut_payload_0_16503 : _zz_dataOut_payload_0_16439);
  assign _zz_dataOut_payload_0_16568 = (_zz_dataOut_payload_0_16441 < _zz_dataOut_payload_0_16505);
  assign _zz_dataOut_payload_0_16569 = (_zz_dataOut_payload_0_16568 ? _zz_dataOut_payload_0_16441 : _zz_dataOut_payload_0_16505);
  assign _zz_dataOut_payload_32_28 = (_zz_dataOut_payload_0_16568 ? _zz_dataOut_payload_0_16505 : _zz_dataOut_payload_0_16441);
  assign _zz_dataOut_payload_0_16570 = (_zz_dataOut_payload_0_16443 < _zz_dataOut_payload_0_16507);
  assign _zz_dataOut_payload_0_16571 = (_zz_dataOut_payload_0_16570 ? _zz_dataOut_payload_0_16443 : _zz_dataOut_payload_0_16507);
  assign _zz_dataOut_payload_32_29 = (_zz_dataOut_payload_0_16570 ? _zz_dataOut_payload_0_16507 : _zz_dataOut_payload_0_16443);
  assign _zz_dataOut_payload_0_16572 = (_zz_dataOut_payload_0_16445 < _zz_dataOut_payload_0_16509);
  assign _zz_dataOut_payload_0_16573 = (_zz_dataOut_payload_0_16572 ? _zz_dataOut_payload_0_16445 : _zz_dataOut_payload_0_16509);
  assign _zz_dataOut_payload_32_30 = (_zz_dataOut_payload_0_16572 ? _zz_dataOut_payload_0_16509 : _zz_dataOut_payload_0_16445);
  assign _zz_dataOut_payload_0_16574 = (_zz_dataOut_payload_0_16447 < _zz_dataOut_payload_0_16511);
  assign _zz_dataOut_payload_0_16575 = (_zz_dataOut_payload_0_16574 ? _zz_dataOut_payload_0_16447 : _zz_dataOut_payload_0_16511);
  assign _zz_dataOut_payload_32_31 = (_zz_dataOut_payload_0_16574 ? _zz_dataOut_payload_0_16511 : _zz_dataOut_payload_0_16447);
  assign _zz_dataOut_payload_0_16576 = (_zz_dataOut_payload_0_16513 < _zz_dataOut_payload_0_16545);
  assign _zz_dataOut_payload_0_16577 = (_zz_dataOut_payload_0_16576 ? _zz_dataOut_payload_0_16513 : _zz_dataOut_payload_0_16545);
  assign _zz_dataOut_payload_16 = (_zz_dataOut_payload_0_16576 ? _zz_dataOut_payload_0_16545 : _zz_dataOut_payload_0_16513);
  assign _zz_dataOut_payload_0_16578 = (_zz_dataOut_payload_0_16515 < _zz_dataOut_payload_0_16547);
  assign _zz_dataOut_payload_0_16579 = (_zz_dataOut_payload_0_16578 ? _zz_dataOut_payload_0_16515 : _zz_dataOut_payload_0_16547);
  assign _zz_dataOut_payload_16_1 = (_zz_dataOut_payload_0_16578 ? _zz_dataOut_payload_0_16547 : _zz_dataOut_payload_0_16515);
  assign _zz_dataOut_payload_0_16580 = (_zz_dataOut_payload_0_16517 < _zz_dataOut_payload_0_16549);
  assign _zz_dataOut_payload_0_16581 = (_zz_dataOut_payload_0_16580 ? _zz_dataOut_payload_0_16517 : _zz_dataOut_payload_0_16549);
  assign _zz_dataOut_payload_16_2 = (_zz_dataOut_payload_0_16580 ? _zz_dataOut_payload_0_16549 : _zz_dataOut_payload_0_16517);
  assign _zz_dataOut_payload_0_16582 = (_zz_dataOut_payload_0_16519 < _zz_dataOut_payload_0_16551);
  assign _zz_dataOut_payload_0_16583 = (_zz_dataOut_payload_0_16582 ? _zz_dataOut_payload_0_16519 : _zz_dataOut_payload_0_16551);
  assign _zz_dataOut_payload_16_3 = (_zz_dataOut_payload_0_16582 ? _zz_dataOut_payload_0_16551 : _zz_dataOut_payload_0_16519);
  assign _zz_dataOut_payload_0_16584 = (_zz_dataOut_payload_0_16521 < _zz_dataOut_payload_0_16553);
  assign _zz_dataOut_payload_0_16585 = (_zz_dataOut_payload_0_16584 ? _zz_dataOut_payload_0_16521 : _zz_dataOut_payload_0_16553);
  assign _zz_dataOut_payload_16_4 = (_zz_dataOut_payload_0_16584 ? _zz_dataOut_payload_0_16553 : _zz_dataOut_payload_0_16521);
  assign _zz_dataOut_payload_0_16586 = (_zz_dataOut_payload_0_16523 < _zz_dataOut_payload_0_16555);
  assign _zz_dataOut_payload_0_16587 = (_zz_dataOut_payload_0_16586 ? _zz_dataOut_payload_0_16523 : _zz_dataOut_payload_0_16555);
  assign _zz_dataOut_payload_16_5 = (_zz_dataOut_payload_0_16586 ? _zz_dataOut_payload_0_16555 : _zz_dataOut_payload_0_16523);
  assign _zz_dataOut_payload_0_16588 = (_zz_dataOut_payload_0_16525 < _zz_dataOut_payload_0_16557);
  assign _zz_dataOut_payload_0_16589 = (_zz_dataOut_payload_0_16588 ? _zz_dataOut_payload_0_16525 : _zz_dataOut_payload_0_16557);
  assign _zz_dataOut_payload_16_6 = (_zz_dataOut_payload_0_16588 ? _zz_dataOut_payload_0_16557 : _zz_dataOut_payload_0_16525);
  assign _zz_dataOut_payload_0_16590 = (_zz_dataOut_payload_0_16527 < _zz_dataOut_payload_0_16559);
  assign _zz_dataOut_payload_0_16591 = (_zz_dataOut_payload_0_16590 ? _zz_dataOut_payload_0_16527 : _zz_dataOut_payload_0_16559);
  assign _zz_dataOut_payload_16_7 = (_zz_dataOut_payload_0_16590 ? _zz_dataOut_payload_0_16559 : _zz_dataOut_payload_0_16527);
  assign _zz_dataOut_payload_0_16592 = (_zz_dataOut_payload_0_16529 < _zz_dataOut_payload_0_16561);
  assign _zz_dataOut_payload_0_16593 = (_zz_dataOut_payload_0_16592 ? _zz_dataOut_payload_0_16529 : _zz_dataOut_payload_0_16561);
  assign _zz_dataOut_payload_16_8 = (_zz_dataOut_payload_0_16592 ? _zz_dataOut_payload_0_16561 : _zz_dataOut_payload_0_16529);
  assign _zz_dataOut_payload_0_16594 = (_zz_dataOut_payload_0_16531 < _zz_dataOut_payload_0_16563);
  assign _zz_dataOut_payload_0_16595 = (_zz_dataOut_payload_0_16594 ? _zz_dataOut_payload_0_16531 : _zz_dataOut_payload_0_16563);
  assign _zz_dataOut_payload_16_9 = (_zz_dataOut_payload_0_16594 ? _zz_dataOut_payload_0_16563 : _zz_dataOut_payload_0_16531);
  assign _zz_dataOut_payload_0_16596 = (_zz_dataOut_payload_0_16533 < _zz_dataOut_payload_0_16565);
  assign _zz_dataOut_payload_0_16597 = (_zz_dataOut_payload_0_16596 ? _zz_dataOut_payload_0_16533 : _zz_dataOut_payload_0_16565);
  assign _zz_dataOut_payload_16_10 = (_zz_dataOut_payload_0_16596 ? _zz_dataOut_payload_0_16565 : _zz_dataOut_payload_0_16533);
  assign _zz_dataOut_payload_0_16598 = (_zz_dataOut_payload_0_16535 < _zz_dataOut_payload_0_16567);
  assign _zz_dataOut_payload_0_16599 = (_zz_dataOut_payload_0_16598 ? _zz_dataOut_payload_0_16535 : _zz_dataOut_payload_0_16567);
  assign _zz_dataOut_payload_16_11 = (_zz_dataOut_payload_0_16598 ? _zz_dataOut_payload_0_16567 : _zz_dataOut_payload_0_16535);
  assign _zz_dataOut_payload_0_16600 = (_zz_dataOut_payload_0_16537 < _zz_dataOut_payload_0_16569);
  assign _zz_dataOut_payload_0_16601 = (_zz_dataOut_payload_0_16600 ? _zz_dataOut_payload_0_16537 : _zz_dataOut_payload_0_16569);
  assign _zz_dataOut_payload_16_12 = (_zz_dataOut_payload_0_16600 ? _zz_dataOut_payload_0_16569 : _zz_dataOut_payload_0_16537);
  assign _zz_dataOut_payload_0_16602 = (_zz_dataOut_payload_0_16539 < _zz_dataOut_payload_0_16571);
  assign _zz_dataOut_payload_0_16603 = (_zz_dataOut_payload_0_16602 ? _zz_dataOut_payload_0_16539 : _zz_dataOut_payload_0_16571);
  assign _zz_dataOut_payload_16_13 = (_zz_dataOut_payload_0_16602 ? _zz_dataOut_payload_0_16571 : _zz_dataOut_payload_0_16539);
  assign _zz_dataOut_payload_0_16604 = (_zz_dataOut_payload_0_16541 < _zz_dataOut_payload_0_16573);
  assign _zz_dataOut_payload_0_16605 = (_zz_dataOut_payload_0_16604 ? _zz_dataOut_payload_0_16541 : _zz_dataOut_payload_0_16573);
  assign _zz_dataOut_payload_16_14 = (_zz_dataOut_payload_0_16604 ? _zz_dataOut_payload_0_16573 : _zz_dataOut_payload_0_16541);
  assign _zz_dataOut_payload_0_16606 = (_zz_dataOut_payload_0_16543 < _zz_dataOut_payload_0_16575);
  assign _zz_dataOut_payload_0_16607 = (_zz_dataOut_payload_0_16606 ? _zz_dataOut_payload_0_16543 : _zz_dataOut_payload_0_16575);
  assign _zz_dataOut_payload_16_15 = (_zz_dataOut_payload_0_16606 ? _zz_dataOut_payload_0_16575 : _zz_dataOut_payload_0_16543);
  assign _zz_dataOut_payload_0_16608 = (_zz_dataOut_payload_0_16577 < _zz_dataOut_payload_0_16593);
  assign _zz_dataOut_payload_0_16609 = (_zz_dataOut_payload_0_16608 ? _zz_dataOut_payload_0_16577 : _zz_dataOut_payload_0_16593);
  assign _zz_dataOut_payload_8 = (_zz_dataOut_payload_0_16608 ? _zz_dataOut_payload_0_16593 : _zz_dataOut_payload_0_16577);
  assign _zz_dataOut_payload_0_16610 = (_zz_dataOut_payload_0_16579 < _zz_dataOut_payload_0_16595);
  assign _zz_dataOut_payload_0_16611 = (_zz_dataOut_payload_0_16610 ? _zz_dataOut_payload_0_16579 : _zz_dataOut_payload_0_16595);
  assign _zz_dataOut_payload_8_1 = (_zz_dataOut_payload_0_16610 ? _zz_dataOut_payload_0_16595 : _zz_dataOut_payload_0_16579);
  assign _zz_dataOut_payload_0_16612 = (_zz_dataOut_payload_0_16581 < _zz_dataOut_payload_0_16597);
  assign _zz_dataOut_payload_0_16613 = (_zz_dataOut_payload_0_16612 ? _zz_dataOut_payload_0_16581 : _zz_dataOut_payload_0_16597);
  assign _zz_dataOut_payload_8_2 = (_zz_dataOut_payload_0_16612 ? _zz_dataOut_payload_0_16597 : _zz_dataOut_payload_0_16581);
  assign _zz_dataOut_payload_0_16614 = (_zz_dataOut_payload_0_16583 < _zz_dataOut_payload_0_16599);
  assign _zz_dataOut_payload_0_16615 = (_zz_dataOut_payload_0_16614 ? _zz_dataOut_payload_0_16583 : _zz_dataOut_payload_0_16599);
  assign _zz_dataOut_payload_8_3 = (_zz_dataOut_payload_0_16614 ? _zz_dataOut_payload_0_16599 : _zz_dataOut_payload_0_16583);
  assign _zz_dataOut_payload_0_16616 = (_zz_dataOut_payload_0_16585 < _zz_dataOut_payload_0_16601);
  assign _zz_dataOut_payload_0_16617 = (_zz_dataOut_payload_0_16616 ? _zz_dataOut_payload_0_16585 : _zz_dataOut_payload_0_16601);
  assign _zz_dataOut_payload_8_4 = (_zz_dataOut_payload_0_16616 ? _zz_dataOut_payload_0_16601 : _zz_dataOut_payload_0_16585);
  assign _zz_dataOut_payload_0_16618 = (_zz_dataOut_payload_0_16587 < _zz_dataOut_payload_0_16603);
  assign _zz_dataOut_payload_0_16619 = (_zz_dataOut_payload_0_16618 ? _zz_dataOut_payload_0_16587 : _zz_dataOut_payload_0_16603);
  assign _zz_dataOut_payload_8_5 = (_zz_dataOut_payload_0_16618 ? _zz_dataOut_payload_0_16603 : _zz_dataOut_payload_0_16587);
  assign _zz_dataOut_payload_0_16620 = (_zz_dataOut_payload_0_16589 < _zz_dataOut_payload_0_16605);
  assign _zz_dataOut_payload_0_16621 = (_zz_dataOut_payload_0_16620 ? _zz_dataOut_payload_0_16589 : _zz_dataOut_payload_0_16605);
  assign _zz_dataOut_payload_8_6 = (_zz_dataOut_payload_0_16620 ? _zz_dataOut_payload_0_16605 : _zz_dataOut_payload_0_16589);
  assign _zz_dataOut_payload_0_16622 = (_zz_dataOut_payload_0_16591 < _zz_dataOut_payload_0_16607);
  assign _zz_dataOut_payload_0_16623 = (_zz_dataOut_payload_0_16622 ? _zz_dataOut_payload_0_16591 : _zz_dataOut_payload_0_16607);
  assign _zz_dataOut_payload_8_7 = (_zz_dataOut_payload_0_16622 ? _zz_dataOut_payload_0_16607 : _zz_dataOut_payload_0_16591);
  assign _zz_dataOut_payload_0_16624 = (_zz_dataOut_payload_0_16609 < _zz_dataOut_payload_0_16617);
  assign _zz_dataOut_payload_0_16625 = (_zz_dataOut_payload_0_16624 ? _zz_dataOut_payload_0_16609 : _zz_dataOut_payload_0_16617);
  assign _zz_dataOut_payload_4 = (_zz_dataOut_payload_0_16624 ? _zz_dataOut_payload_0_16617 : _zz_dataOut_payload_0_16609);
  assign _zz_dataOut_payload_0_16626 = (_zz_dataOut_payload_0_16611 < _zz_dataOut_payload_0_16619);
  assign _zz_dataOut_payload_0_16627 = (_zz_dataOut_payload_0_16626 ? _zz_dataOut_payload_0_16611 : _zz_dataOut_payload_0_16619);
  assign _zz_dataOut_payload_4_1 = (_zz_dataOut_payload_0_16626 ? _zz_dataOut_payload_0_16619 : _zz_dataOut_payload_0_16611);
  assign _zz_dataOut_payload_0_16628 = (_zz_dataOut_payload_0_16613 < _zz_dataOut_payload_0_16621);
  assign _zz_dataOut_payload_0_16629 = (_zz_dataOut_payload_0_16628 ? _zz_dataOut_payload_0_16613 : _zz_dataOut_payload_0_16621);
  assign _zz_dataOut_payload_4_2 = (_zz_dataOut_payload_0_16628 ? _zz_dataOut_payload_0_16621 : _zz_dataOut_payload_0_16613);
  assign _zz_dataOut_payload_0_16630 = (_zz_dataOut_payload_0_16615 < _zz_dataOut_payload_0_16623);
  assign _zz_dataOut_payload_0_16631 = (_zz_dataOut_payload_0_16630 ? _zz_dataOut_payload_0_16615 : _zz_dataOut_payload_0_16623);
  assign _zz_dataOut_payload_4_3 = (_zz_dataOut_payload_0_16630 ? _zz_dataOut_payload_0_16623 : _zz_dataOut_payload_0_16615);
  assign _zz_dataOut_payload_0_16632 = (_zz_dataOut_payload_0_16625 < _zz_dataOut_payload_0_16629);
  assign _zz_dataOut_payload_0_16633 = (_zz_dataOut_payload_0_16632 ? _zz_dataOut_payload_0_16625 : _zz_dataOut_payload_0_16629);
  assign _zz_dataOut_payload_2 = (_zz_dataOut_payload_0_16632 ? _zz_dataOut_payload_0_16629 : _zz_dataOut_payload_0_16625);
  assign _zz_dataOut_payload_0_16634 = (_zz_dataOut_payload_0_16627 < _zz_dataOut_payload_0_16631);
  assign _zz_dataOut_payload_0_16635 = (_zz_dataOut_payload_0_16634 ? _zz_dataOut_payload_0_16627 : _zz_dataOut_payload_0_16631);
  assign _zz_dataOut_payload_2_1 = (_zz_dataOut_payload_0_16634 ? _zz_dataOut_payload_0_16631 : _zz_dataOut_payload_0_16627);
  assign _zz_dataOut_payload_0_16636 = (_zz_dataOut_payload_0_16633 < _zz_dataOut_payload_0_16635);
  assign _zz_dataOut_payload_2_2 = (_zz_dataOut_payload_2 < _zz_dataOut_payload_2_1);
  assign _zz_dataOut_payload_4_4 = (_zz_dataOut_payload_4 < _zz_dataOut_payload_4_2);
  assign _zz_dataOut_payload_4_5 = (_zz_dataOut_payload_4_4 ? _zz_dataOut_payload_4 : _zz_dataOut_payload_4_2);
  assign _zz_dataOut_payload_6 = (_zz_dataOut_payload_4_4 ? _zz_dataOut_payload_4_2 : _zz_dataOut_payload_4);
  assign _zz_dataOut_payload_4_6 = (_zz_dataOut_payload_4_1 < _zz_dataOut_payload_4_3);
  assign _zz_dataOut_payload_4_7 = (_zz_dataOut_payload_4_6 ? _zz_dataOut_payload_4_1 : _zz_dataOut_payload_4_3);
  assign _zz_dataOut_payload_6_1 = (_zz_dataOut_payload_4_6 ? _zz_dataOut_payload_4_3 : _zz_dataOut_payload_4_1);
  assign _zz_dataOut_payload_4_8 = (_zz_dataOut_payload_4_5 < _zz_dataOut_payload_4_7);
  assign _zz_dataOut_payload_6_2 = (_zz_dataOut_payload_6 < _zz_dataOut_payload_6_1);
  assign _zz_dataOut_payload_8_8 = (_zz_dataOut_payload_8 < _zz_dataOut_payload_8_4);
  assign _zz_dataOut_payload_8_9 = (_zz_dataOut_payload_8_8 ? _zz_dataOut_payload_8 : _zz_dataOut_payload_8_4);
  assign _zz_dataOut_payload_12 = (_zz_dataOut_payload_8_8 ? _zz_dataOut_payload_8_4 : _zz_dataOut_payload_8);
  assign _zz_dataOut_payload_8_10 = (_zz_dataOut_payload_8_1 < _zz_dataOut_payload_8_5);
  assign _zz_dataOut_payload_8_11 = (_zz_dataOut_payload_8_10 ? _zz_dataOut_payload_8_1 : _zz_dataOut_payload_8_5);
  assign _zz_dataOut_payload_12_1 = (_zz_dataOut_payload_8_10 ? _zz_dataOut_payload_8_5 : _zz_dataOut_payload_8_1);
  assign _zz_dataOut_payload_8_12 = (_zz_dataOut_payload_8_2 < _zz_dataOut_payload_8_6);
  assign _zz_dataOut_payload_8_13 = (_zz_dataOut_payload_8_12 ? _zz_dataOut_payload_8_2 : _zz_dataOut_payload_8_6);
  assign _zz_dataOut_payload_12_2 = (_zz_dataOut_payload_8_12 ? _zz_dataOut_payload_8_6 : _zz_dataOut_payload_8_2);
  assign _zz_dataOut_payload_8_14 = (_zz_dataOut_payload_8_3 < _zz_dataOut_payload_8_7);
  assign _zz_dataOut_payload_8_15 = (_zz_dataOut_payload_8_14 ? _zz_dataOut_payload_8_3 : _zz_dataOut_payload_8_7);
  assign _zz_dataOut_payload_12_3 = (_zz_dataOut_payload_8_14 ? _zz_dataOut_payload_8_7 : _zz_dataOut_payload_8_3);
  assign _zz_dataOut_payload_8_16 = (_zz_dataOut_payload_8_9 < _zz_dataOut_payload_8_13);
  assign _zz_dataOut_payload_8_17 = (_zz_dataOut_payload_8_16 ? _zz_dataOut_payload_8_9 : _zz_dataOut_payload_8_13);
  assign _zz_dataOut_payload_10 = (_zz_dataOut_payload_8_16 ? _zz_dataOut_payload_8_13 : _zz_dataOut_payload_8_9);
  assign _zz_dataOut_payload_8_18 = (_zz_dataOut_payload_8_11 < _zz_dataOut_payload_8_15);
  assign _zz_dataOut_payload_8_19 = (_zz_dataOut_payload_8_18 ? _zz_dataOut_payload_8_11 : _zz_dataOut_payload_8_15);
  assign _zz_dataOut_payload_10_1 = (_zz_dataOut_payload_8_18 ? _zz_dataOut_payload_8_15 : _zz_dataOut_payload_8_11);
  assign _zz_dataOut_payload_8_20 = (_zz_dataOut_payload_8_17 < _zz_dataOut_payload_8_19);
  assign _zz_dataOut_payload_10_2 = (_zz_dataOut_payload_10 < _zz_dataOut_payload_10_1);
  assign _zz_dataOut_payload_12_4 = (_zz_dataOut_payload_12 < _zz_dataOut_payload_12_2);
  assign _zz_dataOut_payload_12_5 = (_zz_dataOut_payload_12_4 ? _zz_dataOut_payload_12 : _zz_dataOut_payload_12_2);
  assign _zz_dataOut_payload_14 = (_zz_dataOut_payload_12_4 ? _zz_dataOut_payload_12_2 : _zz_dataOut_payload_12);
  assign _zz_dataOut_payload_12_6 = (_zz_dataOut_payload_12_1 < _zz_dataOut_payload_12_3);
  assign _zz_dataOut_payload_12_7 = (_zz_dataOut_payload_12_6 ? _zz_dataOut_payload_12_1 : _zz_dataOut_payload_12_3);
  assign _zz_dataOut_payload_14_1 = (_zz_dataOut_payload_12_6 ? _zz_dataOut_payload_12_3 : _zz_dataOut_payload_12_1);
  assign _zz_dataOut_payload_12_8 = (_zz_dataOut_payload_12_5 < _zz_dataOut_payload_12_7);
  assign _zz_dataOut_payload_14_2 = (_zz_dataOut_payload_14 < _zz_dataOut_payload_14_1);
  assign _zz_dataOut_payload_16_16 = (_zz_dataOut_payload_16 < _zz_dataOut_payload_16_8);
  assign _zz_dataOut_payload_16_17 = (_zz_dataOut_payload_16_16 ? _zz_dataOut_payload_16 : _zz_dataOut_payload_16_8);
  assign _zz_dataOut_payload_24 = (_zz_dataOut_payload_16_16 ? _zz_dataOut_payload_16_8 : _zz_dataOut_payload_16);
  assign _zz_dataOut_payload_16_18 = (_zz_dataOut_payload_16_1 < _zz_dataOut_payload_16_9);
  assign _zz_dataOut_payload_16_19 = (_zz_dataOut_payload_16_18 ? _zz_dataOut_payload_16_1 : _zz_dataOut_payload_16_9);
  assign _zz_dataOut_payload_24_1 = (_zz_dataOut_payload_16_18 ? _zz_dataOut_payload_16_9 : _zz_dataOut_payload_16_1);
  assign _zz_dataOut_payload_16_20 = (_zz_dataOut_payload_16_2 < _zz_dataOut_payload_16_10);
  assign _zz_dataOut_payload_16_21 = (_zz_dataOut_payload_16_20 ? _zz_dataOut_payload_16_2 : _zz_dataOut_payload_16_10);
  assign _zz_dataOut_payload_24_2 = (_zz_dataOut_payload_16_20 ? _zz_dataOut_payload_16_10 : _zz_dataOut_payload_16_2);
  assign _zz_dataOut_payload_16_22 = (_zz_dataOut_payload_16_3 < _zz_dataOut_payload_16_11);
  assign _zz_dataOut_payload_16_23 = (_zz_dataOut_payload_16_22 ? _zz_dataOut_payload_16_3 : _zz_dataOut_payload_16_11);
  assign _zz_dataOut_payload_24_3 = (_zz_dataOut_payload_16_22 ? _zz_dataOut_payload_16_11 : _zz_dataOut_payload_16_3);
  assign _zz_dataOut_payload_16_24 = (_zz_dataOut_payload_16_4 < _zz_dataOut_payload_16_12);
  assign _zz_dataOut_payload_16_25 = (_zz_dataOut_payload_16_24 ? _zz_dataOut_payload_16_4 : _zz_dataOut_payload_16_12);
  assign _zz_dataOut_payload_24_4 = (_zz_dataOut_payload_16_24 ? _zz_dataOut_payload_16_12 : _zz_dataOut_payload_16_4);
  assign _zz_dataOut_payload_16_26 = (_zz_dataOut_payload_16_5 < _zz_dataOut_payload_16_13);
  assign _zz_dataOut_payload_16_27 = (_zz_dataOut_payload_16_26 ? _zz_dataOut_payload_16_5 : _zz_dataOut_payload_16_13);
  assign _zz_dataOut_payload_24_5 = (_zz_dataOut_payload_16_26 ? _zz_dataOut_payload_16_13 : _zz_dataOut_payload_16_5);
  assign _zz_dataOut_payload_16_28 = (_zz_dataOut_payload_16_6 < _zz_dataOut_payload_16_14);
  assign _zz_dataOut_payload_16_29 = (_zz_dataOut_payload_16_28 ? _zz_dataOut_payload_16_6 : _zz_dataOut_payload_16_14);
  assign _zz_dataOut_payload_24_6 = (_zz_dataOut_payload_16_28 ? _zz_dataOut_payload_16_14 : _zz_dataOut_payload_16_6);
  assign _zz_dataOut_payload_16_30 = (_zz_dataOut_payload_16_7 < _zz_dataOut_payload_16_15);
  assign _zz_dataOut_payload_16_31 = (_zz_dataOut_payload_16_30 ? _zz_dataOut_payload_16_7 : _zz_dataOut_payload_16_15);
  assign _zz_dataOut_payload_24_7 = (_zz_dataOut_payload_16_30 ? _zz_dataOut_payload_16_15 : _zz_dataOut_payload_16_7);
  assign _zz_dataOut_payload_16_32 = (_zz_dataOut_payload_16_17 < _zz_dataOut_payload_16_25);
  assign _zz_dataOut_payload_16_33 = (_zz_dataOut_payload_16_32 ? _zz_dataOut_payload_16_17 : _zz_dataOut_payload_16_25);
  assign _zz_dataOut_payload_20 = (_zz_dataOut_payload_16_32 ? _zz_dataOut_payload_16_25 : _zz_dataOut_payload_16_17);
  assign _zz_dataOut_payload_16_34 = (_zz_dataOut_payload_16_19 < _zz_dataOut_payload_16_27);
  assign _zz_dataOut_payload_16_35 = (_zz_dataOut_payload_16_34 ? _zz_dataOut_payload_16_19 : _zz_dataOut_payload_16_27);
  assign _zz_dataOut_payload_20_1 = (_zz_dataOut_payload_16_34 ? _zz_dataOut_payload_16_27 : _zz_dataOut_payload_16_19);
  assign _zz_dataOut_payload_16_36 = (_zz_dataOut_payload_16_21 < _zz_dataOut_payload_16_29);
  assign _zz_dataOut_payload_16_37 = (_zz_dataOut_payload_16_36 ? _zz_dataOut_payload_16_21 : _zz_dataOut_payload_16_29);
  assign _zz_dataOut_payload_20_2 = (_zz_dataOut_payload_16_36 ? _zz_dataOut_payload_16_29 : _zz_dataOut_payload_16_21);
  assign _zz_dataOut_payload_16_38 = (_zz_dataOut_payload_16_23 < _zz_dataOut_payload_16_31);
  assign _zz_dataOut_payload_16_39 = (_zz_dataOut_payload_16_38 ? _zz_dataOut_payload_16_23 : _zz_dataOut_payload_16_31);
  assign _zz_dataOut_payload_20_3 = (_zz_dataOut_payload_16_38 ? _zz_dataOut_payload_16_31 : _zz_dataOut_payload_16_23);
  assign _zz_dataOut_payload_16_40 = (_zz_dataOut_payload_16_33 < _zz_dataOut_payload_16_37);
  assign _zz_dataOut_payload_16_41 = (_zz_dataOut_payload_16_40 ? _zz_dataOut_payload_16_33 : _zz_dataOut_payload_16_37);
  assign _zz_dataOut_payload_18 = (_zz_dataOut_payload_16_40 ? _zz_dataOut_payload_16_37 : _zz_dataOut_payload_16_33);
  assign _zz_dataOut_payload_16_42 = (_zz_dataOut_payload_16_35 < _zz_dataOut_payload_16_39);
  assign _zz_dataOut_payload_16_43 = (_zz_dataOut_payload_16_42 ? _zz_dataOut_payload_16_35 : _zz_dataOut_payload_16_39);
  assign _zz_dataOut_payload_18_1 = (_zz_dataOut_payload_16_42 ? _zz_dataOut_payload_16_39 : _zz_dataOut_payload_16_35);
  assign _zz_dataOut_payload_16_44 = (_zz_dataOut_payload_16_41 < _zz_dataOut_payload_16_43);
  assign _zz_dataOut_payload_18_2 = (_zz_dataOut_payload_18 < _zz_dataOut_payload_18_1);
  assign _zz_dataOut_payload_20_4 = (_zz_dataOut_payload_20 < _zz_dataOut_payload_20_2);
  assign _zz_dataOut_payload_20_5 = (_zz_dataOut_payload_20_4 ? _zz_dataOut_payload_20 : _zz_dataOut_payload_20_2);
  assign _zz_dataOut_payload_22 = (_zz_dataOut_payload_20_4 ? _zz_dataOut_payload_20_2 : _zz_dataOut_payload_20);
  assign _zz_dataOut_payload_20_6 = (_zz_dataOut_payload_20_1 < _zz_dataOut_payload_20_3);
  assign _zz_dataOut_payload_20_7 = (_zz_dataOut_payload_20_6 ? _zz_dataOut_payload_20_1 : _zz_dataOut_payload_20_3);
  assign _zz_dataOut_payload_22_1 = (_zz_dataOut_payload_20_6 ? _zz_dataOut_payload_20_3 : _zz_dataOut_payload_20_1);
  assign _zz_dataOut_payload_20_8 = (_zz_dataOut_payload_20_5 < _zz_dataOut_payload_20_7);
  assign _zz_dataOut_payload_22_2 = (_zz_dataOut_payload_22 < _zz_dataOut_payload_22_1);
  assign _zz_dataOut_payload_24_8 = (_zz_dataOut_payload_24 < _zz_dataOut_payload_24_4);
  assign _zz_dataOut_payload_24_9 = (_zz_dataOut_payload_24_8 ? _zz_dataOut_payload_24 : _zz_dataOut_payload_24_4);
  assign _zz_dataOut_payload_28 = (_zz_dataOut_payload_24_8 ? _zz_dataOut_payload_24_4 : _zz_dataOut_payload_24);
  assign _zz_dataOut_payload_24_10 = (_zz_dataOut_payload_24_1 < _zz_dataOut_payload_24_5);
  assign _zz_dataOut_payload_24_11 = (_zz_dataOut_payload_24_10 ? _zz_dataOut_payload_24_1 : _zz_dataOut_payload_24_5);
  assign _zz_dataOut_payload_28_1 = (_zz_dataOut_payload_24_10 ? _zz_dataOut_payload_24_5 : _zz_dataOut_payload_24_1);
  assign _zz_dataOut_payload_24_12 = (_zz_dataOut_payload_24_2 < _zz_dataOut_payload_24_6);
  assign _zz_dataOut_payload_24_13 = (_zz_dataOut_payload_24_12 ? _zz_dataOut_payload_24_2 : _zz_dataOut_payload_24_6);
  assign _zz_dataOut_payload_28_2 = (_zz_dataOut_payload_24_12 ? _zz_dataOut_payload_24_6 : _zz_dataOut_payload_24_2);
  assign _zz_dataOut_payload_24_14 = (_zz_dataOut_payload_24_3 < _zz_dataOut_payload_24_7);
  assign _zz_dataOut_payload_24_15 = (_zz_dataOut_payload_24_14 ? _zz_dataOut_payload_24_3 : _zz_dataOut_payload_24_7);
  assign _zz_dataOut_payload_28_3 = (_zz_dataOut_payload_24_14 ? _zz_dataOut_payload_24_7 : _zz_dataOut_payload_24_3);
  assign _zz_dataOut_payload_24_16 = (_zz_dataOut_payload_24_9 < _zz_dataOut_payload_24_13);
  assign _zz_dataOut_payload_24_17 = (_zz_dataOut_payload_24_16 ? _zz_dataOut_payload_24_9 : _zz_dataOut_payload_24_13);
  assign _zz_dataOut_payload_26 = (_zz_dataOut_payload_24_16 ? _zz_dataOut_payload_24_13 : _zz_dataOut_payload_24_9);
  assign _zz_dataOut_payload_24_18 = (_zz_dataOut_payload_24_11 < _zz_dataOut_payload_24_15);
  assign _zz_dataOut_payload_24_19 = (_zz_dataOut_payload_24_18 ? _zz_dataOut_payload_24_11 : _zz_dataOut_payload_24_15);
  assign _zz_dataOut_payload_26_1 = (_zz_dataOut_payload_24_18 ? _zz_dataOut_payload_24_15 : _zz_dataOut_payload_24_11);
  assign _zz_dataOut_payload_24_20 = (_zz_dataOut_payload_24_17 < _zz_dataOut_payload_24_19);
  assign _zz_dataOut_payload_26_2 = (_zz_dataOut_payload_26 < _zz_dataOut_payload_26_1);
  assign _zz_dataOut_payload_28_4 = (_zz_dataOut_payload_28 < _zz_dataOut_payload_28_2);
  assign _zz_dataOut_payload_28_5 = (_zz_dataOut_payload_28_4 ? _zz_dataOut_payload_28 : _zz_dataOut_payload_28_2);
  assign _zz_dataOut_payload_30 = (_zz_dataOut_payload_28_4 ? _zz_dataOut_payload_28_2 : _zz_dataOut_payload_28);
  assign _zz_dataOut_payload_28_6 = (_zz_dataOut_payload_28_1 < _zz_dataOut_payload_28_3);
  assign _zz_dataOut_payload_28_7 = (_zz_dataOut_payload_28_6 ? _zz_dataOut_payload_28_1 : _zz_dataOut_payload_28_3);
  assign _zz_dataOut_payload_30_1 = (_zz_dataOut_payload_28_6 ? _zz_dataOut_payload_28_3 : _zz_dataOut_payload_28_1);
  assign _zz_dataOut_payload_28_8 = (_zz_dataOut_payload_28_5 < _zz_dataOut_payload_28_7);
  assign _zz_dataOut_payload_30_2 = (_zz_dataOut_payload_30 < _zz_dataOut_payload_30_1);
  assign _zz_dataOut_payload_32_32 = (_zz_dataOut_payload_32 < _zz_dataOut_payload_32_16);
  assign _zz_dataOut_payload_32_33 = (_zz_dataOut_payload_32_32 ? _zz_dataOut_payload_32 : _zz_dataOut_payload_32_16);
  assign _zz_dataOut_payload_48 = (_zz_dataOut_payload_32_32 ? _zz_dataOut_payload_32_16 : _zz_dataOut_payload_32);
  assign _zz_dataOut_payload_32_34 = (_zz_dataOut_payload_32_1 < _zz_dataOut_payload_32_17);
  assign _zz_dataOut_payload_32_35 = (_zz_dataOut_payload_32_34 ? _zz_dataOut_payload_32_1 : _zz_dataOut_payload_32_17);
  assign _zz_dataOut_payload_48_1 = (_zz_dataOut_payload_32_34 ? _zz_dataOut_payload_32_17 : _zz_dataOut_payload_32_1);
  assign _zz_dataOut_payload_32_36 = (_zz_dataOut_payload_32_2 < _zz_dataOut_payload_32_18);
  assign _zz_dataOut_payload_32_37 = (_zz_dataOut_payload_32_36 ? _zz_dataOut_payload_32_2 : _zz_dataOut_payload_32_18);
  assign _zz_dataOut_payload_48_2 = (_zz_dataOut_payload_32_36 ? _zz_dataOut_payload_32_18 : _zz_dataOut_payload_32_2);
  assign _zz_dataOut_payload_32_38 = (_zz_dataOut_payload_32_3 < _zz_dataOut_payload_32_19);
  assign _zz_dataOut_payload_32_39 = (_zz_dataOut_payload_32_38 ? _zz_dataOut_payload_32_3 : _zz_dataOut_payload_32_19);
  assign _zz_dataOut_payload_48_3 = (_zz_dataOut_payload_32_38 ? _zz_dataOut_payload_32_19 : _zz_dataOut_payload_32_3);
  assign _zz_dataOut_payload_32_40 = (_zz_dataOut_payload_32_4 < _zz_dataOut_payload_32_20);
  assign _zz_dataOut_payload_32_41 = (_zz_dataOut_payload_32_40 ? _zz_dataOut_payload_32_4 : _zz_dataOut_payload_32_20);
  assign _zz_dataOut_payload_48_4 = (_zz_dataOut_payload_32_40 ? _zz_dataOut_payload_32_20 : _zz_dataOut_payload_32_4);
  assign _zz_dataOut_payload_32_42 = (_zz_dataOut_payload_32_5 < _zz_dataOut_payload_32_21);
  assign _zz_dataOut_payload_32_43 = (_zz_dataOut_payload_32_42 ? _zz_dataOut_payload_32_5 : _zz_dataOut_payload_32_21);
  assign _zz_dataOut_payload_48_5 = (_zz_dataOut_payload_32_42 ? _zz_dataOut_payload_32_21 : _zz_dataOut_payload_32_5);
  assign _zz_dataOut_payload_32_44 = (_zz_dataOut_payload_32_6 < _zz_dataOut_payload_32_22);
  assign _zz_dataOut_payload_32_45 = (_zz_dataOut_payload_32_44 ? _zz_dataOut_payload_32_6 : _zz_dataOut_payload_32_22);
  assign _zz_dataOut_payload_48_6 = (_zz_dataOut_payload_32_44 ? _zz_dataOut_payload_32_22 : _zz_dataOut_payload_32_6);
  assign _zz_dataOut_payload_32_46 = (_zz_dataOut_payload_32_7 < _zz_dataOut_payload_32_23);
  assign _zz_dataOut_payload_32_47 = (_zz_dataOut_payload_32_46 ? _zz_dataOut_payload_32_7 : _zz_dataOut_payload_32_23);
  assign _zz_dataOut_payload_48_7 = (_zz_dataOut_payload_32_46 ? _zz_dataOut_payload_32_23 : _zz_dataOut_payload_32_7);
  assign _zz_dataOut_payload_32_48 = (_zz_dataOut_payload_32_8 < _zz_dataOut_payload_32_24);
  assign _zz_dataOut_payload_32_49 = (_zz_dataOut_payload_32_48 ? _zz_dataOut_payload_32_8 : _zz_dataOut_payload_32_24);
  assign _zz_dataOut_payload_48_8 = (_zz_dataOut_payload_32_48 ? _zz_dataOut_payload_32_24 : _zz_dataOut_payload_32_8);
  assign _zz_dataOut_payload_32_50 = (_zz_dataOut_payload_32_9 < _zz_dataOut_payload_32_25);
  assign _zz_dataOut_payload_32_51 = (_zz_dataOut_payload_32_50 ? _zz_dataOut_payload_32_9 : _zz_dataOut_payload_32_25);
  assign _zz_dataOut_payload_48_9 = (_zz_dataOut_payload_32_50 ? _zz_dataOut_payload_32_25 : _zz_dataOut_payload_32_9);
  assign _zz_dataOut_payload_32_52 = (_zz_dataOut_payload_32_10 < _zz_dataOut_payload_32_26);
  assign _zz_dataOut_payload_32_53 = (_zz_dataOut_payload_32_52 ? _zz_dataOut_payload_32_10 : _zz_dataOut_payload_32_26);
  assign _zz_dataOut_payload_48_10 = (_zz_dataOut_payload_32_52 ? _zz_dataOut_payload_32_26 : _zz_dataOut_payload_32_10);
  assign _zz_dataOut_payload_32_54 = (_zz_dataOut_payload_32_11 < _zz_dataOut_payload_32_27);
  assign _zz_dataOut_payload_32_55 = (_zz_dataOut_payload_32_54 ? _zz_dataOut_payload_32_11 : _zz_dataOut_payload_32_27);
  assign _zz_dataOut_payload_48_11 = (_zz_dataOut_payload_32_54 ? _zz_dataOut_payload_32_27 : _zz_dataOut_payload_32_11);
  assign _zz_dataOut_payload_32_56 = (_zz_dataOut_payload_32_12 < _zz_dataOut_payload_32_28);
  assign _zz_dataOut_payload_32_57 = (_zz_dataOut_payload_32_56 ? _zz_dataOut_payload_32_12 : _zz_dataOut_payload_32_28);
  assign _zz_dataOut_payload_48_12 = (_zz_dataOut_payload_32_56 ? _zz_dataOut_payload_32_28 : _zz_dataOut_payload_32_12);
  assign _zz_dataOut_payload_32_58 = (_zz_dataOut_payload_32_13 < _zz_dataOut_payload_32_29);
  assign _zz_dataOut_payload_32_59 = (_zz_dataOut_payload_32_58 ? _zz_dataOut_payload_32_13 : _zz_dataOut_payload_32_29);
  assign _zz_dataOut_payload_48_13 = (_zz_dataOut_payload_32_58 ? _zz_dataOut_payload_32_29 : _zz_dataOut_payload_32_13);
  assign _zz_dataOut_payload_32_60 = (_zz_dataOut_payload_32_14 < _zz_dataOut_payload_32_30);
  assign _zz_dataOut_payload_32_61 = (_zz_dataOut_payload_32_60 ? _zz_dataOut_payload_32_14 : _zz_dataOut_payload_32_30);
  assign _zz_dataOut_payload_48_14 = (_zz_dataOut_payload_32_60 ? _zz_dataOut_payload_32_30 : _zz_dataOut_payload_32_14);
  assign _zz_dataOut_payload_32_62 = (_zz_dataOut_payload_32_15 < _zz_dataOut_payload_32_31);
  assign _zz_dataOut_payload_32_63 = (_zz_dataOut_payload_32_62 ? _zz_dataOut_payload_32_15 : _zz_dataOut_payload_32_31);
  assign _zz_dataOut_payload_48_15 = (_zz_dataOut_payload_32_62 ? _zz_dataOut_payload_32_31 : _zz_dataOut_payload_32_15);
  assign _zz_dataOut_payload_32_64 = (_zz_dataOut_payload_32_33 < _zz_dataOut_payload_32_49);
  assign _zz_dataOut_payload_32_65 = (_zz_dataOut_payload_32_64 ? _zz_dataOut_payload_32_33 : _zz_dataOut_payload_32_49);
  assign _zz_dataOut_payload_40 = (_zz_dataOut_payload_32_64 ? _zz_dataOut_payload_32_49 : _zz_dataOut_payload_32_33);
  assign _zz_dataOut_payload_32_66 = (_zz_dataOut_payload_32_35 < _zz_dataOut_payload_32_51);
  assign _zz_dataOut_payload_32_67 = (_zz_dataOut_payload_32_66 ? _zz_dataOut_payload_32_35 : _zz_dataOut_payload_32_51);
  assign _zz_dataOut_payload_40_1 = (_zz_dataOut_payload_32_66 ? _zz_dataOut_payload_32_51 : _zz_dataOut_payload_32_35);
  assign _zz_dataOut_payload_32_68 = (_zz_dataOut_payload_32_37 < _zz_dataOut_payload_32_53);
  assign _zz_dataOut_payload_32_69 = (_zz_dataOut_payload_32_68 ? _zz_dataOut_payload_32_37 : _zz_dataOut_payload_32_53);
  assign _zz_dataOut_payload_40_2 = (_zz_dataOut_payload_32_68 ? _zz_dataOut_payload_32_53 : _zz_dataOut_payload_32_37);
  assign _zz_dataOut_payload_32_70 = (_zz_dataOut_payload_32_39 < _zz_dataOut_payload_32_55);
  assign _zz_dataOut_payload_32_71 = (_zz_dataOut_payload_32_70 ? _zz_dataOut_payload_32_39 : _zz_dataOut_payload_32_55);
  assign _zz_dataOut_payload_40_3 = (_zz_dataOut_payload_32_70 ? _zz_dataOut_payload_32_55 : _zz_dataOut_payload_32_39);
  assign _zz_dataOut_payload_32_72 = (_zz_dataOut_payload_32_41 < _zz_dataOut_payload_32_57);
  assign _zz_dataOut_payload_32_73 = (_zz_dataOut_payload_32_72 ? _zz_dataOut_payload_32_41 : _zz_dataOut_payload_32_57);
  assign _zz_dataOut_payload_40_4 = (_zz_dataOut_payload_32_72 ? _zz_dataOut_payload_32_57 : _zz_dataOut_payload_32_41);
  assign _zz_dataOut_payload_32_74 = (_zz_dataOut_payload_32_43 < _zz_dataOut_payload_32_59);
  assign _zz_dataOut_payload_32_75 = (_zz_dataOut_payload_32_74 ? _zz_dataOut_payload_32_43 : _zz_dataOut_payload_32_59);
  assign _zz_dataOut_payload_40_5 = (_zz_dataOut_payload_32_74 ? _zz_dataOut_payload_32_59 : _zz_dataOut_payload_32_43);
  assign _zz_dataOut_payload_32_76 = (_zz_dataOut_payload_32_45 < _zz_dataOut_payload_32_61);
  assign _zz_dataOut_payload_32_77 = (_zz_dataOut_payload_32_76 ? _zz_dataOut_payload_32_45 : _zz_dataOut_payload_32_61);
  assign _zz_dataOut_payload_40_6 = (_zz_dataOut_payload_32_76 ? _zz_dataOut_payload_32_61 : _zz_dataOut_payload_32_45);
  assign _zz_dataOut_payload_32_78 = (_zz_dataOut_payload_32_47 < _zz_dataOut_payload_32_63);
  assign _zz_dataOut_payload_32_79 = (_zz_dataOut_payload_32_78 ? _zz_dataOut_payload_32_47 : _zz_dataOut_payload_32_63);
  assign _zz_dataOut_payload_40_7 = (_zz_dataOut_payload_32_78 ? _zz_dataOut_payload_32_63 : _zz_dataOut_payload_32_47);
  assign _zz_dataOut_payload_32_80 = (_zz_dataOut_payload_32_65 < _zz_dataOut_payload_32_73);
  assign _zz_dataOut_payload_32_81 = (_zz_dataOut_payload_32_80 ? _zz_dataOut_payload_32_65 : _zz_dataOut_payload_32_73);
  assign _zz_dataOut_payload_36 = (_zz_dataOut_payload_32_80 ? _zz_dataOut_payload_32_73 : _zz_dataOut_payload_32_65);
  assign _zz_dataOut_payload_32_82 = (_zz_dataOut_payload_32_67 < _zz_dataOut_payload_32_75);
  assign _zz_dataOut_payload_32_83 = (_zz_dataOut_payload_32_82 ? _zz_dataOut_payload_32_67 : _zz_dataOut_payload_32_75);
  assign _zz_dataOut_payload_36_1 = (_zz_dataOut_payload_32_82 ? _zz_dataOut_payload_32_75 : _zz_dataOut_payload_32_67);
  assign _zz_dataOut_payload_32_84 = (_zz_dataOut_payload_32_69 < _zz_dataOut_payload_32_77);
  assign _zz_dataOut_payload_32_85 = (_zz_dataOut_payload_32_84 ? _zz_dataOut_payload_32_69 : _zz_dataOut_payload_32_77);
  assign _zz_dataOut_payload_36_2 = (_zz_dataOut_payload_32_84 ? _zz_dataOut_payload_32_77 : _zz_dataOut_payload_32_69);
  assign _zz_dataOut_payload_32_86 = (_zz_dataOut_payload_32_71 < _zz_dataOut_payload_32_79);
  assign _zz_dataOut_payload_32_87 = (_zz_dataOut_payload_32_86 ? _zz_dataOut_payload_32_71 : _zz_dataOut_payload_32_79);
  assign _zz_dataOut_payload_36_3 = (_zz_dataOut_payload_32_86 ? _zz_dataOut_payload_32_79 : _zz_dataOut_payload_32_71);
  assign _zz_dataOut_payload_32_88 = (_zz_dataOut_payload_32_81 < _zz_dataOut_payload_32_85);
  assign _zz_dataOut_payload_32_89 = (_zz_dataOut_payload_32_88 ? _zz_dataOut_payload_32_81 : _zz_dataOut_payload_32_85);
  assign _zz_dataOut_payload_34 = (_zz_dataOut_payload_32_88 ? _zz_dataOut_payload_32_85 : _zz_dataOut_payload_32_81);
  assign _zz_dataOut_payload_32_90 = (_zz_dataOut_payload_32_83 < _zz_dataOut_payload_32_87);
  assign _zz_dataOut_payload_32_91 = (_zz_dataOut_payload_32_90 ? _zz_dataOut_payload_32_83 : _zz_dataOut_payload_32_87);
  assign _zz_dataOut_payload_34_1 = (_zz_dataOut_payload_32_90 ? _zz_dataOut_payload_32_87 : _zz_dataOut_payload_32_83);
  assign _zz_dataOut_payload_32_92 = (_zz_dataOut_payload_32_89 < _zz_dataOut_payload_32_91);
  assign _zz_dataOut_payload_34_2 = (_zz_dataOut_payload_34 < _zz_dataOut_payload_34_1);
  assign _zz_dataOut_payload_36_4 = (_zz_dataOut_payload_36 < _zz_dataOut_payload_36_2);
  assign _zz_dataOut_payload_36_5 = (_zz_dataOut_payload_36_4 ? _zz_dataOut_payload_36 : _zz_dataOut_payload_36_2);
  assign _zz_dataOut_payload_38 = (_zz_dataOut_payload_36_4 ? _zz_dataOut_payload_36_2 : _zz_dataOut_payload_36);
  assign _zz_dataOut_payload_36_6 = (_zz_dataOut_payload_36_1 < _zz_dataOut_payload_36_3);
  assign _zz_dataOut_payload_36_7 = (_zz_dataOut_payload_36_6 ? _zz_dataOut_payload_36_1 : _zz_dataOut_payload_36_3);
  assign _zz_dataOut_payload_38_1 = (_zz_dataOut_payload_36_6 ? _zz_dataOut_payload_36_3 : _zz_dataOut_payload_36_1);
  assign _zz_dataOut_payload_36_8 = (_zz_dataOut_payload_36_5 < _zz_dataOut_payload_36_7);
  assign _zz_dataOut_payload_38_2 = (_zz_dataOut_payload_38 < _zz_dataOut_payload_38_1);
  assign _zz_dataOut_payload_40_8 = (_zz_dataOut_payload_40 < _zz_dataOut_payload_40_4);
  assign _zz_dataOut_payload_40_9 = (_zz_dataOut_payload_40_8 ? _zz_dataOut_payload_40 : _zz_dataOut_payload_40_4);
  assign _zz_dataOut_payload_44 = (_zz_dataOut_payload_40_8 ? _zz_dataOut_payload_40_4 : _zz_dataOut_payload_40);
  assign _zz_dataOut_payload_40_10 = (_zz_dataOut_payload_40_1 < _zz_dataOut_payload_40_5);
  assign _zz_dataOut_payload_40_11 = (_zz_dataOut_payload_40_10 ? _zz_dataOut_payload_40_1 : _zz_dataOut_payload_40_5);
  assign _zz_dataOut_payload_44_1 = (_zz_dataOut_payload_40_10 ? _zz_dataOut_payload_40_5 : _zz_dataOut_payload_40_1);
  assign _zz_dataOut_payload_40_12 = (_zz_dataOut_payload_40_2 < _zz_dataOut_payload_40_6);
  assign _zz_dataOut_payload_40_13 = (_zz_dataOut_payload_40_12 ? _zz_dataOut_payload_40_2 : _zz_dataOut_payload_40_6);
  assign _zz_dataOut_payload_44_2 = (_zz_dataOut_payload_40_12 ? _zz_dataOut_payload_40_6 : _zz_dataOut_payload_40_2);
  assign _zz_dataOut_payload_40_14 = (_zz_dataOut_payload_40_3 < _zz_dataOut_payload_40_7);
  assign _zz_dataOut_payload_40_15 = (_zz_dataOut_payload_40_14 ? _zz_dataOut_payload_40_3 : _zz_dataOut_payload_40_7);
  assign _zz_dataOut_payload_44_3 = (_zz_dataOut_payload_40_14 ? _zz_dataOut_payload_40_7 : _zz_dataOut_payload_40_3);
  assign _zz_dataOut_payload_40_16 = (_zz_dataOut_payload_40_9 < _zz_dataOut_payload_40_13);
  assign _zz_dataOut_payload_40_17 = (_zz_dataOut_payload_40_16 ? _zz_dataOut_payload_40_9 : _zz_dataOut_payload_40_13);
  assign _zz_dataOut_payload_42 = (_zz_dataOut_payload_40_16 ? _zz_dataOut_payload_40_13 : _zz_dataOut_payload_40_9);
  assign _zz_dataOut_payload_40_18 = (_zz_dataOut_payload_40_11 < _zz_dataOut_payload_40_15);
  assign _zz_dataOut_payload_40_19 = (_zz_dataOut_payload_40_18 ? _zz_dataOut_payload_40_11 : _zz_dataOut_payload_40_15);
  assign _zz_dataOut_payload_42_1 = (_zz_dataOut_payload_40_18 ? _zz_dataOut_payload_40_15 : _zz_dataOut_payload_40_11);
  assign _zz_dataOut_payload_40_20 = (_zz_dataOut_payload_40_17 < _zz_dataOut_payload_40_19);
  assign _zz_dataOut_payload_42_2 = (_zz_dataOut_payload_42 < _zz_dataOut_payload_42_1);
  assign _zz_dataOut_payload_44_4 = (_zz_dataOut_payload_44 < _zz_dataOut_payload_44_2);
  assign _zz_dataOut_payload_44_5 = (_zz_dataOut_payload_44_4 ? _zz_dataOut_payload_44 : _zz_dataOut_payload_44_2);
  assign _zz_dataOut_payload_46 = (_zz_dataOut_payload_44_4 ? _zz_dataOut_payload_44_2 : _zz_dataOut_payload_44);
  assign _zz_dataOut_payload_44_6 = (_zz_dataOut_payload_44_1 < _zz_dataOut_payload_44_3);
  assign _zz_dataOut_payload_44_7 = (_zz_dataOut_payload_44_6 ? _zz_dataOut_payload_44_1 : _zz_dataOut_payload_44_3);
  assign _zz_dataOut_payload_46_1 = (_zz_dataOut_payload_44_6 ? _zz_dataOut_payload_44_3 : _zz_dataOut_payload_44_1);
  assign _zz_dataOut_payload_44_8 = (_zz_dataOut_payload_44_5 < _zz_dataOut_payload_44_7);
  assign _zz_dataOut_payload_46_2 = (_zz_dataOut_payload_46 < _zz_dataOut_payload_46_1);
  assign _zz_dataOut_payload_48_16 = (_zz_dataOut_payload_48 < _zz_dataOut_payload_48_8);
  assign _zz_dataOut_payload_48_17 = (_zz_dataOut_payload_48_16 ? _zz_dataOut_payload_48 : _zz_dataOut_payload_48_8);
  assign _zz_dataOut_payload_56 = (_zz_dataOut_payload_48_16 ? _zz_dataOut_payload_48_8 : _zz_dataOut_payload_48);
  assign _zz_dataOut_payload_48_18 = (_zz_dataOut_payload_48_1 < _zz_dataOut_payload_48_9);
  assign _zz_dataOut_payload_48_19 = (_zz_dataOut_payload_48_18 ? _zz_dataOut_payload_48_1 : _zz_dataOut_payload_48_9);
  assign _zz_dataOut_payload_56_1 = (_zz_dataOut_payload_48_18 ? _zz_dataOut_payload_48_9 : _zz_dataOut_payload_48_1);
  assign _zz_dataOut_payload_48_20 = (_zz_dataOut_payload_48_2 < _zz_dataOut_payload_48_10);
  assign _zz_dataOut_payload_48_21 = (_zz_dataOut_payload_48_20 ? _zz_dataOut_payload_48_2 : _zz_dataOut_payload_48_10);
  assign _zz_dataOut_payload_56_2 = (_zz_dataOut_payload_48_20 ? _zz_dataOut_payload_48_10 : _zz_dataOut_payload_48_2);
  assign _zz_dataOut_payload_48_22 = (_zz_dataOut_payload_48_3 < _zz_dataOut_payload_48_11);
  assign _zz_dataOut_payload_48_23 = (_zz_dataOut_payload_48_22 ? _zz_dataOut_payload_48_3 : _zz_dataOut_payload_48_11);
  assign _zz_dataOut_payload_56_3 = (_zz_dataOut_payload_48_22 ? _zz_dataOut_payload_48_11 : _zz_dataOut_payload_48_3);
  assign _zz_dataOut_payload_48_24 = (_zz_dataOut_payload_48_4 < _zz_dataOut_payload_48_12);
  assign _zz_dataOut_payload_48_25 = (_zz_dataOut_payload_48_24 ? _zz_dataOut_payload_48_4 : _zz_dataOut_payload_48_12);
  assign _zz_dataOut_payload_56_4 = (_zz_dataOut_payload_48_24 ? _zz_dataOut_payload_48_12 : _zz_dataOut_payload_48_4);
  assign _zz_dataOut_payload_48_26 = (_zz_dataOut_payload_48_5 < _zz_dataOut_payload_48_13);
  assign _zz_dataOut_payload_48_27 = (_zz_dataOut_payload_48_26 ? _zz_dataOut_payload_48_5 : _zz_dataOut_payload_48_13);
  assign _zz_dataOut_payload_56_5 = (_zz_dataOut_payload_48_26 ? _zz_dataOut_payload_48_13 : _zz_dataOut_payload_48_5);
  assign _zz_dataOut_payload_48_28 = (_zz_dataOut_payload_48_6 < _zz_dataOut_payload_48_14);
  assign _zz_dataOut_payload_48_29 = (_zz_dataOut_payload_48_28 ? _zz_dataOut_payload_48_6 : _zz_dataOut_payload_48_14);
  assign _zz_dataOut_payload_56_6 = (_zz_dataOut_payload_48_28 ? _zz_dataOut_payload_48_14 : _zz_dataOut_payload_48_6);
  assign _zz_dataOut_payload_48_30 = (_zz_dataOut_payload_48_7 < _zz_dataOut_payload_48_15);
  assign _zz_dataOut_payload_48_31 = (_zz_dataOut_payload_48_30 ? _zz_dataOut_payload_48_7 : _zz_dataOut_payload_48_15);
  assign _zz_dataOut_payload_56_7 = (_zz_dataOut_payload_48_30 ? _zz_dataOut_payload_48_15 : _zz_dataOut_payload_48_7);
  assign _zz_dataOut_payload_48_32 = (_zz_dataOut_payload_48_17 < _zz_dataOut_payload_48_25);
  assign _zz_dataOut_payload_48_33 = (_zz_dataOut_payload_48_32 ? _zz_dataOut_payload_48_17 : _zz_dataOut_payload_48_25);
  assign _zz_dataOut_payload_52 = (_zz_dataOut_payload_48_32 ? _zz_dataOut_payload_48_25 : _zz_dataOut_payload_48_17);
  assign _zz_dataOut_payload_48_34 = (_zz_dataOut_payload_48_19 < _zz_dataOut_payload_48_27);
  assign _zz_dataOut_payload_48_35 = (_zz_dataOut_payload_48_34 ? _zz_dataOut_payload_48_19 : _zz_dataOut_payload_48_27);
  assign _zz_dataOut_payload_52_1 = (_zz_dataOut_payload_48_34 ? _zz_dataOut_payload_48_27 : _zz_dataOut_payload_48_19);
  assign _zz_dataOut_payload_48_36 = (_zz_dataOut_payload_48_21 < _zz_dataOut_payload_48_29);
  assign _zz_dataOut_payload_48_37 = (_zz_dataOut_payload_48_36 ? _zz_dataOut_payload_48_21 : _zz_dataOut_payload_48_29);
  assign _zz_dataOut_payload_52_2 = (_zz_dataOut_payload_48_36 ? _zz_dataOut_payload_48_29 : _zz_dataOut_payload_48_21);
  assign _zz_dataOut_payload_48_38 = (_zz_dataOut_payload_48_23 < _zz_dataOut_payload_48_31);
  assign _zz_dataOut_payload_48_39 = (_zz_dataOut_payload_48_38 ? _zz_dataOut_payload_48_23 : _zz_dataOut_payload_48_31);
  assign _zz_dataOut_payload_52_3 = (_zz_dataOut_payload_48_38 ? _zz_dataOut_payload_48_31 : _zz_dataOut_payload_48_23);
  assign _zz_dataOut_payload_48_40 = (_zz_dataOut_payload_48_33 < _zz_dataOut_payload_48_37);
  assign _zz_dataOut_payload_48_41 = (_zz_dataOut_payload_48_40 ? _zz_dataOut_payload_48_33 : _zz_dataOut_payload_48_37);
  assign _zz_dataOut_payload_50 = (_zz_dataOut_payload_48_40 ? _zz_dataOut_payload_48_37 : _zz_dataOut_payload_48_33);
  assign _zz_dataOut_payload_48_42 = (_zz_dataOut_payload_48_35 < _zz_dataOut_payload_48_39);
  assign _zz_dataOut_payload_48_43 = (_zz_dataOut_payload_48_42 ? _zz_dataOut_payload_48_35 : _zz_dataOut_payload_48_39);
  assign _zz_dataOut_payload_50_1 = (_zz_dataOut_payload_48_42 ? _zz_dataOut_payload_48_39 : _zz_dataOut_payload_48_35);
  assign _zz_dataOut_payload_48_44 = (_zz_dataOut_payload_48_41 < _zz_dataOut_payload_48_43);
  assign _zz_dataOut_payload_50_2 = (_zz_dataOut_payload_50 < _zz_dataOut_payload_50_1);
  assign _zz_dataOut_payload_52_4 = (_zz_dataOut_payload_52 < _zz_dataOut_payload_52_2);
  assign _zz_dataOut_payload_52_5 = (_zz_dataOut_payload_52_4 ? _zz_dataOut_payload_52 : _zz_dataOut_payload_52_2);
  assign _zz_dataOut_payload_54 = (_zz_dataOut_payload_52_4 ? _zz_dataOut_payload_52_2 : _zz_dataOut_payload_52);
  assign _zz_dataOut_payload_52_6 = (_zz_dataOut_payload_52_1 < _zz_dataOut_payload_52_3);
  assign _zz_dataOut_payload_52_7 = (_zz_dataOut_payload_52_6 ? _zz_dataOut_payload_52_1 : _zz_dataOut_payload_52_3);
  assign _zz_dataOut_payload_54_1 = (_zz_dataOut_payload_52_6 ? _zz_dataOut_payload_52_3 : _zz_dataOut_payload_52_1);
  assign _zz_dataOut_payload_52_8 = (_zz_dataOut_payload_52_5 < _zz_dataOut_payload_52_7);
  assign _zz_dataOut_payload_54_2 = (_zz_dataOut_payload_54 < _zz_dataOut_payload_54_1);
  assign _zz_dataOut_payload_56_8 = (_zz_dataOut_payload_56 < _zz_dataOut_payload_56_4);
  assign _zz_dataOut_payload_56_9 = (_zz_dataOut_payload_56_8 ? _zz_dataOut_payload_56 : _zz_dataOut_payload_56_4);
  assign _zz_dataOut_payload_60 = (_zz_dataOut_payload_56_8 ? _zz_dataOut_payload_56_4 : _zz_dataOut_payload_56);
  assign _zz_dataOut_payload_56_10 = (_zz_dataOut_payload_56_1 < _zz_dataOut_payload_56_5);
  assign _zz_dataOut_payload_56_11 = (_zz_dataOut_payload_56_10 ? _zz_dataOut_payload_56_1 : _zz_dataOut_payload_56_5);
  assign _zz_dataOut_payload_60_1 = (_zz_dataOut_payload_56_10 ? _zz_dataOut_payload_56_5 : _zz_dataOut_payload_56_1);
  assign _zz_dataOut_payload_56_12 = (_zz_dataOut_payload_56_2 < _zz_dataOut_payload_56_6);
  assign _zz_dataOut_payload_56_13 = (_zz_dataOut_payload_56_12 ? _zz_dataOut_payload_56_2 : _zz_dataOut_payload_56_6);
  assign _zz_dataOut_payload_60_2 = (_zz_dataOut_payload_56_12 ? _zz_dataOut_payload_56_6 : _zz_dataOut_payload_56_2);
  assign _zz_dataOut_payload_56_14 = (_zz_dataOut_payload_56_3 < _zz_dataOut_payload_56_7);
  assign _zz_dataOut_payload_56_15 = (_zz_dataOut_payload_56_14 ? _zz_dataOut_payload_56_3 : _zz_dataOut_payload_56_7);
  assign _zz_dataOut_payload_60_3 = (_zz_dataOut_payload_56_14 ? _zz_dataOut_payload_56_7 : _zz_dataOut_payload_56_3);
  assign _zz_dataOut_payload_56_16 = (_zz_dataOut_payload_56_9 < _zz_dataOut_payload_56_13);
  assign _zz_dataOut_payload_56_17 = (_zz_dataOut_payload_56_16 ? _zz_dataOut_payload_56_9 : _zz_dataOut_payload_56_13);
  assign _zz_dataOut_payload_58 = (_zz_dataOut_payload_56_16 ? _zz_dataOut_payload_56_13 : _zz_dataOut_payload_56_9);
  assign _zz_dataOut_payload_56_18 = (_zz_dataOut_payload_56_11 < _zz_dataOut_payload_56_15);
  assign _zz_dataOut_payload_56_19 = (_zz_dataOut_payload_56_18 ? _zz_dataOut_payload_56_11 : _zz_dataOut_payload_56_15);
  assign _zz_dataOut_payload_58_1 = (_zz_dataOut_payload_56_18 ? _zz_dataOut_payload_56_15 : _zz_dataOut_payload_56_11);
  assign _zz_dataOut_payload_56_20 = (_zz_dataOut_payload_56_17 < _zz_dataOut_payload_56_19);
  assign _zz_dataOut_payload_58_2 = (_zz_dataOut_payload_58 < _zz_dataOut_payload_58_1);
  assign _zz_dataOut_payload_60_4 = (_zz_dataOut_payload_60 < _zz_dataOut_payload_60_2);
  assign _zz_dataOut_payload_60_5 = (_zz_dataOut_payload_60_4 ? _zz_dataOut_payload_60 : _zz_dataOut_payload_60_2);
  assign _zz_dataOut_payload_62 = (_zz_dataOut_payload_60_4 ? _zz_dataOut_payload_60_2 : _zz_dataOut_payload_60);
  assign _zz_dataOut_payload_60_6 = (_zz_dataOut_payload_60_1 < _zz_dataOut_payload_60_3);
  assign _zz_dataOut_payload_60_7 = (_zz_dataOut_payload_60_6 ? _zz_dataOut_payload_60_1 : _zz_dataOut_payload_60_3);
  assign _zz_dataOut_payload_62_1 = (_zz_dataOut_payload_60_6 ? _zz_dataOut_payload_60_3 : _zz_dataOut_payload_60_1);
  assign _zz_dataOut_payload_60_8 = (_zz_dataOut_payload_60_5 < _zz_dataOut_payload_60_7);
  assign _zz_dataOut_payload_62_2 = (_zz_dataOut_payload_62 < _zz_dataOut_payload_62_1);
  assign _zz_dataOut_payload_64_64 = (_zz_dataOut_payload_64 < _zz_dataOut_payload_64_32);
  assign _zz_dataOut_payload_64_65 = (_zz_dataOut_payload_64_64 ? _zz_dataOut_payload_64 : _zz_dataOut_payload_64_32);
  assign _zz_dataOut_payload_96 = (_zz_dataOut_payload_64_64 ? _zz_dataOut_payload_64_32 : _zz_dataOut_payload_64);
  assign _zz_dataOut_payload_64_66 = (_zz_dataOut_payload_64_1 < _zz_dataOut_payload_64_33);
  assign _zz_dataOut_payload_64_67 = (_zz_dataOut_payload_64_66 ? _zz_dataOut_payload_64_1 : _zz_dataOut_payload_64_33);
  assign _zz_dataOut_payload_96_1 = (_zz_dataOut_payload_64_66 ? _zz_dataOut_payload_64_33 : _zz_dataOut_payload_64_1);
  assign _zz_dataOut_payload_64_68 = (_zz_dataOut_payload_64_2 < _zz_dataOut_payload_64_34);
  assign _zz_dataOut_payload_64_69 = (_zz_dataOut_payload_64_68 ? _zz_dataOut_payload_64_2 : _zz_dataOut_payload_64_34);
  assign _zz_dataOut_payload_96_2 = (_zz_dataOut_payload_64_68 ? _zz_dataOut_payload_64_34 : _zz_dataOut_payload_64_2);
  assign _zz_dataOut_payload_64_70 = (_zz_dataOut_payload_64_3 < _zz_dataOut_payload_64_35);
  assign _zz_dataOut_payload_64_71 = (_zz_dataOut_payload_64_70 ? _zz_dataOut_payload_64_3 : _zz_dataOut_payload_64_35);
  assign _zz_dataOut_payload_96_3 = (_zz_dataOut_payload_64_70 ? _zz_dataOut_payload_64_35 : _zz_dataOut_payload_64_3);
  assign _zz_dataOut_payload_64_72 = (_zz_dataOut_payload_64_4 < _zz_dataOut_payload_64_36);
  assign _zz_dataOut_payload_64_73 = (_zz_dataOut_payload_64_72 ? _zz_dataOut_payload_64_4 : _zz_dataOut_payload_64_36);
  assign _zz_dataOut_payload_96_4 = (_zz_dataOut_payload_64_72 ? _zz_dataOut_payload_64_36 : _zz_dataOut_payload_64_4);
  assign _zz_dataOut_payload_64_74 = (_zz_dataOut_payload_64_5 < _zz_dataOut_payload_64_37);
  assign _zz_dataOut_payload_64_75 = (_zz_dataOut_payload_64_74 ? _zz_dataOut_payload_64_5 : _zz_dataOut_payload_64_37);
  assign _zz_dataOut_payload_96_5 = (_zz_dataOut_payload_64_74 ? _zz_dataOut_payload_64_37 : _zz_dataOut_payload_64_5);
  assign _zz_dataOut_payload_64_76 = (_zz_dataOut_payload_64_6 < _zz_dataOut_payload_64_38);
  assign _zz_dataOut_payload_64_77 = (_zz_dataOut_payload_64_76 ? _zz_dataOut_payload_64_6 : _zz_dataOut_payload_64_38);
  assign _zz_dataOut_payload_96_6 = (_zz_dataOut_payload_64_76 ? _zz_dataOut_payload_64_38 : _zz_dataOut_payload_64_6);
  assign _zz_dataOut_payload_64_78 = (_zz_dataOut_payload_64_7 < _zz_dataOut_payload_64_39);
  assign _zz_dataOut_payload_64_79 = (_zz_dataOut_payload_64_78 ? _zz_dataOut_payload_64_7 : _zz_dataOut_payload_64_39);
  assign _zz_dataOut_payload_96_7 = (_zz_dataOut_payload_64_78 ? _zz_dataOut_payload_64_39 : _zz_dataOut_payload_64_7);
  assign _zz_dataOut_payload_64_80 = (_zz_dataOut_payload_64_8 < _zz_dataOut_payload_64_40);
  assign _zz_dataOut_payload_64_81 = (_zz_dataOut_payload_64_80 ? _zz_dataOut_payload_64_8 : _zz_dataOut_payload_64_40);
  assign _zz_dataOut_payload_96_8 = (_zz_dataOut_payload_64_80 ? _zz_dataOut_payload_64_40 : _zz_dataOut_payload_64_8);
  assign _zz_dataOut_payload_64_82 = (_zz_dataOut_payload_64_9 < _zz_dataOut_payload_64_41);
  assign _zz_dataOut_payload_64_83 = (_zz_dataOut_payload_64_82 ? _zz_dataOut_payload_64_9 : _zz_dataOut_payload_64_41);
  assign _zz_dataOut_payload_96_9 = (_zz_dataOut_payload_64_82 ? _zz_dataOut_payload_64_41 : _zz_dataOut_payload_64_9);
  assign _zz_dataOut_payload_64_84 = (_zz_dataOut_payload_64_10 < _zz_dataOut_payload_64_42);
  assign _zz_dataOut_payload_64_85 = (_zz_dataOut_payload_64_84 ? _zz_dataOut_payload_64_10 : _zz_dataOut_payload_64_42);
  assign _zz_dataOut_payload_96_10 = (_zz_dataOut_payload_64_84 ? _zz_dataOut_payload_64_42 : _zz_dataOut_payload_64_10);
  assign _zz_dataOut_payload_64_86 = (_zz_dataOut_payload_64_11 < _zz_dataOut_payload_64_43);
  assign _zz_dataOut_payload_64_87 = (_zz_dataOut_payload_64_86 ? _zz_dataOut_payload_64_11 : _zz_dataOut_payload_64_43);
  assign _zz_dataOut_payload_96_11 = (_zz_dataOut_payload_64_86 ? _zz_dataOut_payload_64_43 : _zz_dataOut_payload_64_11);
  assign _zz_dataOut_payload_64_88 = (_zz_dataOut_payload_64_12 < _zz_dataOut_payload_64_44);
  assign _zz_dataOut_payload_64_89 = (_zz_dataOut_payload_64_88 ? _zz_dataOut_payload_64_12 : _zz_dataOut_payload_64_44);
  assign _zz_dataOut_payload_96_12 = (_zz_dataOut_payload_64_88 ? _zz_dataOut_payload_64_44 : _zz_dataOut_payload_64_12);
  assign _zz_dataOut_payload_64_90 = (_zz_dataOut_payload_64_13 < _zz_dataOut_payload_64_45);
  assign _zz_dataOut_payload_64_91 = (_zz_dataOut_payload_64_90 ? _zz_dataOut_payload_64_13 : _zz_dataOut_payload_64_45);
  assign _zz_dataOut_payload_96_13 = (_zz_dataOut_payload_64_90 ? _zz_dataOut_payload_64_45 : _zz_dataOut_payload_64_13);
  assign _zz_dataOut_payload_64_92 = (_zz_dataOut_payload_64_14 < _zz_dataOut_payload_64_46);
  assign _zz_dataOut_payload_64_93 = (_zz_dataOut_payload_64_92 ? _zz_dataOut_payload_64_14 : _zz_dataOut_payload_64_46);
  assign _zz_dataOut_payload_96_14 = (_zz_dataOut_payload_64_92 ? _zz_dataOut_payload_64_46 : _zz_dataOut_payload_64_14);
  assign _zz_dataOut_payload_64_94 = (_zz_dataOut_payload_64_15 < _zz_dataOut_payload_64_47);
  assign _zz_dataOut_payload_64_95 = (_zz_dataOut_payload_64_94 ? _zz_dataOut_payload_64_15 : _zz_dataOut_payload_64_47);
  assign _zz_dataOut_payload_96_15 = (_zz_dataOut_payload_64_94 ? _zz_dataOut_payload_64_47 : _zz_dataOut_payload_64_15);
  assign _zz_dataOut_payload_64_96 = (_zz_dataOut_payload_64_16 < _zz_dataOut_payload_64_48);
  assign _zz_dataOut_payload_64_97 = (_zz_dataOut_payload_64_96 ? _zz_dataOut_payload_64_16 : _zz_dataOut_payload_64_48);
  assign _zz_dataOut_payload_96_16 = (_zz_dataOut_payload_64_96 ? _zz_dataOut_payload_64_48 : _zz_dataOut_payload_64_16);
  assign _zz_dataOut_payload_64_98 = (_zz_dataOut_payload_64_17 < _zz_dataOut_payload_64_49);
  assign _zz_dataOut_payload_64_99 = (_zz_dataOut_payload_64_98 ? _zz_dataOut_payload_64_17 : _zz_dataOut_payload_64_49);
  assign _zz_dataOut_payload_96_17 = (_zz_dataOut_payload_64_98 ? _zz_dataOut_payload_64_49 : _zz_dataOut_payload_64_17);
  assign _zz_dataOut_payload_64_100 = (_zz_dataOut_payload_64_18 < _zz_dataOut_payload_64_50);
  assign _zz_dataOut_payload_64_101 = (_zz_dataOut_payload_64_100 ? _zz_dataOut_payload_64_18 : _zz_dataOut_payload_64_50);
  assign _zz_dataOut_payload_96_18 = (_zz_dataOut_payload_64_100 ? _zz_dataOut_payload_64_50 : _zz_dataOut_payload_64_18);
  assign _zz_dataOut_payload_64_102 = (_zz_dataOut_payload_64_19 < _zz_dataOut_payload_64_51);
  assign _zz_dataOut_payload_64_103 = (_zz_dataOut_payload_64_102 ? _zz_dataOut_payload_64_19 : _zz_dataOut_payload_64_51);
  assign _zz_dataOut_payload_96_19 = (_zz_dataOut_payload_64_102 ? _zz_dataOut_payload_64_51 : _zz_dataOut_payload_64_19);
  assign _zz_dataOut_payload_64_104 = (_zz_dataOut_payload_64_20 < _zz_dataOut_payload_64_52);
  assign _zz_dataOut_payload_64_105 = (_zz_dataOut_payload_64_104 ? _zz_dataOut_payload_64_20 : _zz_dataOut_payload_64_52);
  assign _zz_dataOut_payload_96_20 = (_zz_dataOut_payload_64_104 ? _zz_dataOut_payload_64_52 : _zz_dataOut_payload_64_20);
  assign _zz_dataOut_payload_64_106 = (_zz_dataOut_payload_64_21 < _zz_dataOut_payload_64_53);
  assign _zz_dataOut_payload_64_107 = (_zz_dataOut_payload_64_106 ? _zz_dataOut_payload_64_21 : _zz_dataOut_payload_64_53);
  assign _zz_dataOut_payload_96_21 = (_zz_dataOut_payload_64_106 ? _zz_dataOut_payload_64_53 : _zz_dataOut_payload_64_21);
  assign _zz_dataOut_payload_64_108 = (_zz_dataOut_payload_64_22 < _zz_dataOut_payload_64_54);
  assign _zz_dataOut_payload_64_109 = (_zz_dataOut_payload_64_108 ? _zz_dataOut_payload_64_22 : _zz_dataOut_payload_64_54);
  assign _zz_dataOut_payload_96_22 = (_zz_dataOut_payload_64_108 ? _zz_dataOut_payload_64_54 : _zz_dataOut_payload_64_22);
  assign _zz_dataOut_payload_64_110 = (_zz_dataOut_payload_64_23 < _zz_dataOut_payload_64_55);
  assign _zz_dataOut_payload_64_111 = (_zz_dataOut_payload_64_110 ? _zz_dataOut_payload_64_23 : _zz_dataOut_payload_64_55);
  assign _zz_dataOut_payload_96_23 = (_zz_dataOut_payload_64_110 ? _zz_dataOut_payload_64_55 : _zz_dataOut_payload_64_23);
  assign _zz_dataOut_payload_64_112 = (_zz_dataOut_payload_64_24 < _zz_dataOut_payload_64_56);
  assign _zz_dataOut_payload_64_113 = (_zz_dataOut_payload_64_112 ? _zz_dataOut_payload_64_24 : _zz_dataOut_payload_64_56);
  assign _zz_dataOut_payload_96_24 = (_zz_dataOut_payload_64_112 ? _zz_dataOut_payload_64_56 : _zz_dataOut_payload_64_24);
  assign _zz_dataOut_payload_64_114 = (_zz_dataOut_payload_64_25 < _zz_dataOut_payload_64_57);
  assign _zz_dataOut_payload_64_115 = (_zz_dataOut_payload_64_114 ? _zz_dataOut_payload_64_25 : _zz_dataOut_payload_64_57);
  assign _zz_dataOut_payload_96_25 = (_zz_dataOut_payload_64_114 ? _zz_dataOut_payload_64_57 : _zz_dataOut_payload_64_25);
  assign _zz_dataOut_payload_64_116 = (_zz_dataOut_payload_64_26 < _zz_dataOut_payload_64_58);
  assign _zz_dataOut_payload_64_117 = (_zz_dataOut_payload_64_116 ? _zz_dataOut_payload_64_26 : _zz_dataOut_payload_64_58);
  assign _zz_dataOut_payload_96_26 = (_zz_dataOut_payload_64_116 ? _zz_dataOut_payload_64_58 : _zz_dataOut_payload_64_26);
  assign _zz_dataOut_payload_64_118 = (_zz_dataOut_payload_64_27 < _zz_dataOut_payload_64_59);
  assign _zz_dataOut_payload_64_119 = (_zz_dataOut_payload_64_118 ? _zz_dataOut_payload_64_27 : _zz_dataOut_payload_64_59);
  assign _zz_dataOut_payload_96_27 = (_zz_dataOut_payload_64_118 ? _zz_dataOut_payload_64_59 : _zz_dataOut_payload_64_27);
  assign _zz_dataOut_payload_64_120 = (_zz_dataOut_payload_64_28 < _zz_dataOut_payload_64_60);
  assign _zz_dataOut_payload_64_121 = (_zz_dataOut_payload_64_120 ? _zz_dataOut_payload_64_28 : _zz_dataOut_payload_64_60);
  assign _zz_dataOut_payload_96_28 = (_zz_dataOut_payload_64_120 ? _zz_dataOut_payload_64_60 : _zz_dataOut_payload_64_28);
  assign _zz_dataOut_payload_64_122 = (_zz_dataOut_payload_64_29 < _zz_dataOut_payload_64_61);
  assign _zz_dataOut_payload_64_123 = (_zz_dataOut_payload_64_122 ? _zz_dataOut_payload_64_29 : _zz_dataOut_payload_64_61);
  assign _zz_dataOut_payload_96_29 = (_zz_dataOut_payload_64_122 ? _zz_dataOut_payload_64_61 : _zz_dataOut_payload_64_29);
  assign _zz_dataOut_payload_64_124 = (_zz_dataOut_payload_64_30 < _zz_dataOut_payload_64_62);
  assign _zz_dataOut_payload_64_125 = (_zz_dataOut_payload_64_124 ? _zz_dataOut_payload_64_30 : _zz_dataOut_payload_64_62);
  assign _zz_dataOut_payload_96_30 = (_zz_dataOut_payload_64_124 ? _zz_dataOut_payload_64_62 : _zz_dataOut_payload_64_30);
  assign _zz_dataOut_payload_64_126 = (_zz_dataOut_payload_64_31 < _zz_dataOut_payload_64_63);
  assign _zz_dataOut_payload_64_127 = (_zz_dataOut_payload_64_126 ? _zz_dataOut_payload_64_31 : _zz_dataOut_payload_64_63);
  assign _zz_dataOut_payload_96_31 = (_zz_dataOut_payload_64_126 ? _zz_dataOut_payload_64_63 : _zz_dataOut_payload_64_31);
  assign _zz_dataOut_payload_64_128 = (_zz_dataOut_payload_64_65 < _zz_dataOut_payload_64_97);
  assign _zz_dataOut_payload_64_129 = (_zz_dataOut_payload_64_128 ? _zz_dataOut_payload_64_65 : _zz_dataOut_payload_64_97);
  assign _zz_dataOut_payload_80 = (_zz_dataOut_payload_64_128 ? _zz_dataOut_payload_64_97 : _zz_dataOut_payload_64_65);
  assign _zz_dataOut_payload_64_130 = (_zz_dataOut_payload_64_67 < _zz_dataOut_payload_64_99);
  assign _zz_dataOut_payload_64_131 = (_zz_dataOut_payload_64_130 ? _zz_dataOut_payload_64_67 : _zz_dataOut_payload_64_99);
  assign _zz_dataOut_payload_80_1 = (_zz_dataOut_payload_64_130 ? _zz_dataOut_payload_64_99 : _zz_dataOut_payload_64_67);
  assign _zz_dataOut_payload_64_132 = (_zz_dataOut_payload_64_69 < _zz_dataOut_payload_64_101);
  assign _zz_dataOut_payload_64_133 = (_zz_dataOut_payload_64_132 ? _zz_dataOut_payload_64_69 : _zz_dataOut_payload_64_101);
  assign _zz_dataOut_payload_80_2 = (_zz_dataOut_payload_64_132 ? _zz_dataOut_payload_64_101 : _zz_dataOut_payload_64_69);
  assign _zz_dataOut_payload_64_134 = (_zz_dataOut_payload_64_71 < _zz_dataOut_payload_64_103);
  assign _zz_dataOut_payload_64_135 = (_zz_dataOut_payload_64_134 ? _zz_dataOut_payload_64_71 : _zz_dataOut_payload_64_103);
  assign _zz_dataOut_payload_80_3 = (_zz_dataOut_payload_64_134 ? _zz_dataOut_payload_64_103 : _zz_dataOut_payload_64_71);
  assign _zz_dataOut_payload_64_136 = (_zz_dataOut_payload_64_73 < _zz_dataOut_payload_64_105);
  assign _zz_dataOut_payload_64_137 = (_zz_dataOut_payload_64_136 ? _zz_dataOut_payload_64_73 : _zz_dataOut_payload_64_105);
  assign _zz_dataOut_payload_80_4 = (_zz_dataOut_payload_64_136 ? _zz_dataOut_payload_64_105 : _zz_dataOut_payload_64_73);
  assign _zz_dataOut_payload_64_138 = (_zz_dataOut_payload_64_75 < _zz_dataOut_payload_64_107);
  assign _zz_dataOut_payload_64_139 = (_zz_dataOut_payload_64_138 ? _zz_dataOut_payload_64_75 : _zz_dataOut_payload_64_107);
  assign _zz_dataOut_payload_80_5 = (_zz_dataOut_payload_64_138 ? _zz_dataOut_payload_64_107 : _zz_dataOut_payload_64_75);
  assign _zz_dataOut_payload_64_140 = (_zz_dataOut_payload_64_77 < _zz_dataOut_payload_64_109);
  assign _zz_dataOut_payload_64_141 = (_zz_dataOut_payload_64_140 ? _zz_dataOut_payload_64_77 : _zz_dataOut_payload_64_109);
  assign _zz_dataOut_payload_80_6 = (_zz_dataOut_payload_64_140 ? _zz_dataOut_payload_64_109 : _zz_dataOut_payload_64_77);
  assign _zz_dataOut_payload_64_142 = (_zz_dataOut_payload_64_79 < _zz_dataOut_payload_64_111);
  assign _zz_dataOut_payload_64_143 = (_zz_dataOut_payload_64_142 ? _zz_dataOut_payload_64_79 : _zz_dataOut_payload_64_111);
  assign _zz_dataOut_payload_80_7 = (_zz_dataOut_payload_64_142 ? _zz_dataOut_payload_64_111 : _zz_dataOut_payload_64_79);
  assign _zz_dataOut_payload_64_144 = (_zz_dataOut_payload_64_81 < _zz_dataOut_payload_64_113);
  assign _zz_dataOut_payload_64_145 = (_zz_dataOut_payload_64_144 ? _zz_dataOut_payload_64_81 : _zz_dataOut_payload_64_113);
  assign _zz_dataOut_payload_80_8 = (_zz_dataOut_payload_64_144 ? _zz_dataOut_payload_64_113 : _zz_dataOut_payload_64_81);
  assign _zz_dataOut_payload_64_146 = (_zz_dataOut_payload_64_83 < _zz_dataOut_payload_64_115);
  assign _zz_dataOut_payload_64_147 = (_zz_dataOut_payload_64_146 ? _zz_dataOut_payload_64_83 : _zz_dataOut_payload_64_115);
  assign _zz_dataOut_payload_80_9 = (_zz_dataOut_payload_64_146 ? _zz_dataOut_payload_64_115 : _zz_dataOut_payload_64_83);
  assign _zz_dataOut_payload_64_148 = (_zz_dataOut_payload_64_85 < _zz_dataOut_payload_64_117);
  assign _zz_dataOut_payload_64_149 = (_zz_dataOut_payload_64_148 ? _zz_dataOut_payload_64_85 : _zz_dataOut_payload_64_117);
  assign _zz_dataOut_payload_80_10 = (_zz_dataOut_payload_64_148 ? _zz_dataOut_payload_64_117 : _zz_dataOut_payload_64_85);
  assign _zz_dataOut_payload_64_150 = (_zz_dataOut_payload_64_87 < _zz_dataOut_payload_64_119);
  assign _zz_dataOut_payload_64_151 = (_zz_dataOut_payload_64_150 ? _zz_dataOut_payload_64_87 : _zz_dataOut_payload_64_119);
  assign _zz_dataOut_payload_80_11 = (_zz_dataOut_payload_64_150 ? _zz_dataOut_payload_64_119 : _zz_dataOut_payload_64_87);
  assign _zz_dataOut_payload_64_152 = (_zz_dataOut_payload_64_89 < _zz_dataOut_payload_64_121);
  assign _zz_dataOut_payload_64_153 = (_zz_dataOut_payload_64_152 ? _zz_dataOut_payload_64_89 : _zz_dataOut_payload_64_121);
  assign _zz_dataOut_payload_80_12 = (_zz_dataOut_payload_64_152 ? _zz_dataOut_payload_64_121 : _zz_dataOut_payload_64_89);
  assign _zz_dataOut_payload_64_154 = (_zz_dataOut_payload_64_91 < _zz_dataOut_payload_64_123);
  assign _zz_dataOut_payload_64_155 = (_zz_dataOut_payload_64_154 ? _zz_dataOut_payload_64_91 : _zz_dataOut_payload_64_123);
  assign _zz_dataOut_payload_80_13 = (_zz_dataOut_payload_64_154 ? _zz_dataOut_payload_64_123 : _zz_dataOut_payload_64_91);
  assign _zz_dataOut_payload_64_156 = (_zz_dataOut_payload_64_93 < _zz_dataOut_payload_64_125);
  assign _zz_dataOut_payload_64_157 = (_zz_dataOut_payload_64_156 ? _zz_dataOut_payload_64_93 : _zz_dataOut_payload_64_125);
  assign _zz_dataOut_payload_80_14 = (_zz_dataOut_payload_64_156 ? _zz_dataOut_payload_64_125 : _zz_dataOut_payload_64_93);
  assign _zz_dataOut_payload_64_158 = (_zz_dataOut_payload_64_95 < _zz_dataOut_payload_64_127);
  assign _zz_dataOut_payload_64_159 = (_zz_dataOut_payload_64_158 ? _zz_dataOut_payload_64_95 : _zz_dataOut_payload_64_127);
  assign _zz_dataOut_payload_80_15 = (_zz_dataOut_payload_64_158 ? _zz_dataOut_payload_64_127 : _zz_dataOut_payload_64_95);
  assign _zz_dataOut_payload_64_160 = (_zz_dataOut_payload_64_129 < _zz_dataOut_payload_64_145);
  assign _zz_dataOut_payload_64_161 = (_zz_dataOut_payload_64_160 ? _zz_dataOut_payload_64_129 : _zz_dataOut_payload_64_145);
  assign _zz_dataOut_payload_72 = (_zz_dataOut_payload_64_160 ? _zz_dataOut_payload_64_145 : _zz_dataOut_payload_64_129);
  assign _zz_dataOut_payload_64_162 = (_zz_dataOut_payload_64_131 < _zz_dataOut_payload_64_147);
  assign _zz_dataOut_payload_64_163 = (_zz_dataOut_payload_64_162 ? _zz_dataOut_payload_64_131 : _zz_dataOut_payload_64_147);
  assign _zz_dataOut_payload_72_1 = (_zz_dataOut_payload_64_162 ? _zz_dataOut_payload_64_147 : _zz_dataOut_payload_64_131);
  assign _zz_dataOut_payload_64_164 = (_zz_dataOut_payload_64_133 < _zz_dataOut_payload_64_149);
  assign _zz_dataOut_payload_64_165 = (_zz_dataOut_payload_64_164 ? _zz_dataOut_payload_64_133 : _zz_dataOut_payload_64_149);
  assign _zz_dataOut_payload_72_2 = (_zz_dataOut_payload_64_164 ? _zz_dataOut_payload_64_149 : _zz_dataOut_payload_64_133);
  assign _zz_dataOut_payload_64_166 = (_zz_dataOut_payload_64_135 < _zz_dataOut_payload_64_151);
  assign _zz_dataOut_payload_64_167 = (_zz_dataOut_payload_64_166 ? _zz_dataOut_payload_64_135 : _zz_dataOut_payload_64_151);
  assign _zz_dataOut_payload_72_3 = (_zz_dataOut_payload_64_166 ? _zz_dataOut_payload_64_151 : _zz_dataOut_payload_64_135);
  assign _zz_dataOut_payload_64_168 = (_zz_dataOut_payload_64_137 < _zz_dataOut_payload_64_153);
  assign _zz_dataOut_payload_64_169 = (_zz_dataOut_payload_64_168 ? _zz_dataOut_payload_64_137 : _zz_dataOut_payload_64_153);
  assign _zz_dataOut_payload_72_4 = (_zz_dataOut_payload_64_168 ? _zz_dataOut_payload_64_153 : _zz_dataOut_payload_64_137);
  assign _zz_dataOut_payload_64_170 = (_zz_dataOut_payload_64_139 < _zz_dataOut_payload_64_155);
  assign _zz_dataOut_payload_64_171 = (_zz_dataOut_payload_64_170 ? _zz_dataOut_payload_64_139 : _zz_dataOut_payload_64_155);
  assign _zz_dataOut_payload_72_5 = (_zz_dataOut_payload_64_170 ? _zz_dataOut_payload_64_155 : _zz_dataOut_payload_64_139);
  assign _zz_dataOut_payload_64_172 = (_zz_dataOut_payload_64_141 < _zz_dataOut_payload_64_157);
  assign _zz_dataOut_payload_64_173 = (_zz_dataOut_payload_64_172 ? _zz_dataOut_payload_64_141 : _zz_dataOut_payload_64_157);
  assign _zz_dataOut_payload_72_6 = (_zz_dataOut_payload_64_172 ? _zz_dataOut_payload_64_157 : _zz_dataOut_payload_64_141);
  assign _zz_dataOut_payload_64_174 = (_zz_dataOut_payload_64_143 < _zz_dataOut_payload_64_159);
  assign _zz_dataOut_payload_64_175 = (_zz_dataOut_payload_64_174 ? _zz_dataOut_payload_64_143 : _zz_dataOut_payload_64_159);
  assign _zz_dataOut_payload_72_7 = (_zz_dataOut_payload_64_174 ? _zz_dataOut_payload_64_159 : _zz_dataOut_payload_64_143);
  assign _zz_dataOut_payload_64_176 = (_zz_dataOut_payload_64_161 < _zz_dataOut_payload_64_169);
  assign _zz_dataOut_payload_64_177 = (_zz_dataOut_payload_64_176 ? _zz_dataOut_payload_64_161 : _zz_dataOut_payload_64_169);
  assign _zz_dataOut_payload_68 = (_zz_dataOut_payload_64_176 ? _zz_dataOut_payload_64_169 : _zz_dataOut_payload_64_161);
  assign _zz_dataOut_payload_64_178 = (_zz_dataOut_payload_64_163 < _zz_dataOut_payload_64_171);
  assign _zz_dataOut_payload_64_179 = (_zz_dataOut_payload_64_178 ? _zz_dataOut_payload_64_163 : _zz_dataOut_payload_64_171);
  assign _zz_dataOut_payload_68_1 = (_zz_dataOut_payload_64_178 ? _zz_dataOut_payload_64_171 : _zz_dataOut_payload_64_163);
  assign _zz_dataOut_payload_64_180 = (_zz_dataOut_payload_64_165 < _zz_dataOut_payload_64_173);
  assign _zz_dataOut_payload_64_181 = (_zz_dataOut_payload_64_180 ? _zz_dataOut_payload_64_165 : _zz_dataOut_payload_64_173);
  assign _zz_dataOut_payload_68_2 = (_zz_dataOut_payload_64_180 ? _zz_dataOut_payload_64_173 : _zz_dataOut_payload_64_165);
  assign _zz_dataOut_payload_64_182 = (_zz_dataOut_payload_64_167 < _zz_dataOut_payload_64_175);
  assign _zz_dataOut_payload_64_183 = (_zz_dataOut_payload_64_182 ? _zz_dataOut_payload_64_167 : _zz_dataOut_payload_64_175);
  assign _zz_dataOut_payload_68_3 = (_zz_dataOut_payload_64_182 ? _zz_dataOut_payload_64_175 : _zz_dataOut_payload_64_167);
  assign _zz_dataOut_payload_64_184 = (_zz_dataOut_payload_64_177 < _zz_dataOut_payload_64_181);
  assign _zz_dataOut_payload_64_185 = (_zz_dataOut_payload_64_184 ? _zz_dataOut_payload_64_177 : _zz_dataOut_payload_64_181);
  assign _zz_dataOut_payload_66 = (_zz_dataOut_payload_64_184 ? _zz_dataOut_payload_64_181 : _zz_dataOut_payload_64_177);
  assign _zz_dataOut_payload_64_186 = (_zz_dataOut_payload_64_179 < _zz_dataOut_payload_64_183);
  assign _zz_dataOut_payload_64_187 = (_zz_dataOut_payload_64_186 ? _zz_dataOut_payload_64_179 : _zz_dataOut_payload_64_183);
  assign _zz_dataOut_payload_66_1 = (_zz_dataOut_payload_64_186 ? _zz_dataOut_payload_64_183 : _zz_dataOut_payload_64_179);
  assign _zz_dataOut_payload_64_188 = (_zz_dataOut_payload_64_185 < _zz_dataOut_payload_64_187);
  assign _zz_dataOut_payload_66_2 = (_zz_dataOut_payload_66 < _zz_dataOut_payload_66_1);
  assign _zz_dataOut_payload_68_4 = (_zz_dataOut_payload_68 < _zz_dataOut_payload_68_2);
  assign _zz_dataOut_payload_68_5 = (_zz_dataOut_payload_68_4 ? _zz_dataOut_payload_68 : _zz_dataOut_payload_68_2);
  assign _zz_dataOut_payload_70 = (_zz_dataOut_payload_68_4 ? _zz_dataOut_payload_68_2 : _zz_dataOut_payload_68);
  assign _zz_dataOut_payload_68_6 = (_zz_dataOut_payload_68_1 < _zz_dataOut_payload_68_3);
  assign _zz_dataOut_payload_68_7 = (_zz_dataOut_payload_68_6 ? _zz_dataOut_payload_68_1 : _zz_dataOut_payload_68_3);
  assign _zz_dataOut_payload_70_1 = (_zz_dataOut_payload_68_6 ? _zz_dataOut_payload_68_3 : _zz_dataOut_payload_68_1);
  assign _zz_dataOut_payload_68_8 = (_zz_dataOut_payload_68_5 < _zz_dataOut_payload_68_7);
  assign _zz_dataOut_payload_70_2 = (_zz_dataOut_payload_70 < _zz_dataOut_payload_70_1);
  assign _zz_dataOut_payload_72_8 = (_zz_dataOut_payload_72 < _zz_dataOut_payload_72_4);
  assign _zz_dataOut_payload_72_9 = (_zz_dataOut_payload_72_8 ? _zz_dataOut_payload_72 : _zz_dataOut_payload_72_4);
  assign _zz_dataOut_payload_76 = (_zz_dataOut_payload_72_8 ? _zz_dataOut_payload_72_4 : _zz_dataOut_payload_72);
  assign _zz_dataOut_payload_72_10 = (_zz_dataOut_payload_72_1 < _zz_dataOut_payload_72_5);
  assign _zz_dataOut_payload_72_11 = (_zz_dataOut_payload_72_10 ? _zz_dataOut_payload_72_1 : _zz_dataOut_payload_72_5);
  assign _zz_dataOut_payload_76_1 = (_zz_dataOut_payload_72_10 ? _zz_dataOut_payload_72_5 : _zz_dataOut_payload_72_1);
  assign _zz_dataOut_payload_72_12 = (_zz_dataOut_payload_72_2 < _zz_dataOut_payload_72_6);
  assign _zz_dataOut_payload_72_13 = (_zz_dataOut_payload_72_12 ? _zz_dataOut_payload_72_2 : _zz_dataOut_payload_72_6);
  assign _zz_dataOut_payload_76_2 = (_zz_dataOut_payload_72_12 ? _zz_dataOut_payload_72_6 : _zz_dataOut_payload_72_2);
  assign _zz_dataOut_payload_72_14 = (_zz_dataOut_payload_72_3 < _zz_dataOut_payload_72_7);
  assign _zz_dataOut_payload_72_15 = (_zz_dataOut_payload_72_14 ? _zz_dataOut_payload_72_3 : _zz_dataOut_payload_72_7);
  assign _zz_dataOut_payload_76_3 = (_zz_dataOut_payload_72_14 ? _zz_dataOut_payload_72_7 : _zz_dataOut_payload_72_3);
  assign _zz_dataOut_payload_72_16 = (_zz_dataOut_payload_72_9 < _zz_dataOut_payload_72_13);
  assign _zz_dataOut_payload_72_17 = (_zz_dataOut_payload_72_16 ? _zz_dataOut_payload_72_9 : _zz_dataOut_payload_72_13);
  assign _zz_dataOut_payload_74 = (_zz_dataOut_payload_72_16 ? _zz_dataOut_payload_72_13 : _zz_dataOut_payload_72_9);
  assign _zz_dataOut_payload_72_18 = (_zz_dataOut_payload_72_11 < _zz_dataOut_payload_72_15);
  assign _zz_dataOut_payload_72_19 = (_zz_dataOut_payload_72_18 ? _zz_dataOut_payload_72_11 : _zz_dataOut_payload_72_15);
  assign _zz_dataOut_payload_74_1 = (_zz_dataOut_payload_72_18 ? _zz_dataOut_payload_72_15 : _zz_dataOut_payload_72_11);
  assign _zz_dataOut_payload_72_20 = (_zz_dataOut_payload_72_17 < _zz_dataOut_payload_72_19);
  assign _zz_dataOut_payload_74_2 = (_zz_dataOut_payload_74 < _zz_dataOut_payload_74_1);
  assign _zz_dataOut_payload_76_4 = (_zz_dataOut_payload_76 < _zz_dataOut_payload_76_2);
  assign _zz_dataOut_payload_76_5 = (_zz_dataOut_payload_76_4 ? _zz_dataOut_payload_76 : _zz_dataOut_payload_76_2);
  assign _zz_dataOut_payload_78 = (_zz_dataOut_payload_76_4 ? _zz_dataOut_payload_76_2 : _zz_dataOut_payload_76);
  assign _zz_dataOut_payload_76_6 = (_zz_dataOut_payload_76_1 < _zz_dataOut_payload_76_3);
  assign _zz_dataOut_payload_76_7 = (_zz_dataOut_payload_76_6 ? _zz_dataOut_payload_76_1 : _zz_dataOut_payload_76_3);
  assign _zz_dataOut_payload_78_1 = (_zz_dataOut_payload_76_6 ? _zz_dataOut_payload_76_3 : _zz_dataOut_payload_76_1);
  assign _zz_dataOut_payload_76_8 = (_zz_dataOut_payload_76_5 < _zz_dataOut_payload_76_7);
  assign _zz_dataOut_payload_78_2 = (_zz_dataOut_payload_78 < _zz_dataOut_payload_78_1);
  assign _zz_dataOut_payload_80_16 = (_zz_dataOut_payload_80 < _zz_dataOut_payload_80_8);
  assign _zz_dataOut_payload_80_17 = (_zz_dataOut_payload_80_16 ? _zz_dataOut_payload_80 : _zz_dataOut_payload_80_8);
  assign _zz_dataOut_payload_88 = (_zz_dataOut_payload_80_16 ? _zz_dataOut_payload_80_8 : _zz_dataOut_payload_80);
  assign _zz_dataOut_payload_80_18 = (_zz_dataOut_payload_80_1 < _zz_dataOut_payload_80_9);
  assign _zz_dataOut_payload_80_19 = (_zz_dataOut_payload_80_18 ? _zz_dataOut_payload_80_1 : _zz_dataOut_payload_80_9);
  assign _zz_dataOut_payload_88_1 = (_zz_dataOut_payload_80_18 ? _zz_dataOut_payload_80_9 : _zz_dataOut_payload_80_1);
  assign _zz_dataOut_payload_80_20 = (_zz_dataOut_payload_80_2 < _zz_dataOut_payload_80_10);
  assign _zz_dataOut_payload_80_21 = (_zz_dataOut_payload_80_20 ? _zz_dataOut_payload_80_2 : _zz_dataOut_payload_80_10);
  assign _zz_dataOut_payload_88_2 = (_zz_dataOut_payload_80_20 ? _zz_dataOut_payload_80_10 : _zz_dataOut_payload_80_2);
  assign _zz_dataOut_payload_80_22 = (_zz_dataOut_payload_80_3 < _zz_dataOut_payload_80_11);
  assign _zz_dataOut_payload_80_23 = (_zz_dataOut_payload_80_22 ? _zz_dataOut_payload_80_3 : _zz_dataOut_payload_80_11);
  assign _zz_dataOut_payload_88_3 = (_zz_dataOut_payload_80_22 ? _zz_dataOut_payload_80_11 : _zz_dataOut_payload_80_3);
  assign _zz_dataOut_payload_80_24 = (_zz_dataOut_payload_80_4 < _zz_dataOut_payload_80_12);
  assign _zz_dataOut_payload_80_25 = (_zz_dataOut_payload_80_24 ? _zz_dataOut_payload_80_4 : _zz_dataOut_payload_80_12);
  assign _zz_dataOut_payload_88_4 = (_zz_dataOut_payload_80_24 ? _zz_dataOut_payload_80_12 : _zz_dataOut_payload_80_4);
  assign _zz_dataOut_payload_80_26 = (_zz_dataOut_payload_80_5 < _zz_dataOut_payload_80_13);
  assign _zz_dataOut_payload_80_27 = (_zz_dataOut_payload_80_26 ? _zz_dataOut_payload_80_5 : _zz_dataOut_payload_80_13);
  assign _zz_dataOut_payload_88_5 = (_zz_dataOut_payload_80_26 ? _zz_dataOut_payload_80_13 : _zz_dataOut_payload_80_5);
  assign _zz_dataOut_payload_80_28 = (_zz_dataOut_payload_80_6 < _zz_dataOut_payload_80_14);
  assign _zz_dataOut_payload_80_29 = (_zz_dataOut_payload_80_28 ? _zz_dataOut_payload_80_6 : _zz_dataOut_payload_80_14);
  assign _zz_dataOut_payload_88_6 = (_zz_dataOut_payload_80_28 ? _zz_dataOut_payload_80_14 : _zz_dataOut_payload_80_6);
  assign _zz_dataOut_payload_80_30 = (_zz_dataOut_payload_80_7 < _zz_dataOut_payload_80_15);
  assign _zz_dataOut_payload_80_31 = (_zz_dataOut_payload_80_30 ? _zz_dataOut_payload_80_7 : _zz_dataOut_payload_80_15);
  assign _zz_dataOut_payload_88_7 = (_zz_dataOut_payload_80_30 ? _zz_dataOut_payload_80_15 : _zz_dataOut_payload_80_7);
  assign _zz_dataOut_payload_80_32 = (_zz_dataOut_payload_80_17 < _zz_dataOut_payload_80_25);
  assign _zz_dataOut_payload_80_33 = (_zz_dataOut_payload_80_32 ? _zz_dataOut_payload_80_17 : _zz_dataOut_payload_80_25);
  assign _zz_dataOut_payload_84 = (_zz_dataOut_payload_80_32 ? _zz_dataOut_payload_80_25 : _zz_dataOut_payload_80_17);
  assign _zz_dataOut_payload_80_34 = (_zz_dataOut_payload_80_19 < _zz_dataOut_payload_80_27);
  assign _zz_dataOut_payload_80_35 = (_zz_dataOut_payload_80_34 ? _zz_dataOut_payload_80_19 : _zz_dataOut_payload_80_27);
  assign _zz_dataOut_payload_84_1 = (_zz_dataOut_payload_80_34 ? _zz_dataOut_payload_80_27 : _zz_dataOut_payload_80_19);
  assign _zz_dataOut_payload_80_36 = (_zz_dataOut_payload_80_21 < _zz_dataOut_payload_80_29);
  assign _zz_dataOut_payload_80_37 = (_zz_dataOut_payload_80_36 ? _zz_dataOut_payload_80_21 : _zz_dataOut_payload_80_29);
  assign _zz_dataOut_payload_84_2 = (_zz_dataOut_payload_80_36 ? _zz_dataOut_payload_80_29 : _zz_dataOut_payload_80_21);
  assign _zz_dataOut_payload_80_38 = (_zz_dataOut_payload_80_23 < _zz_dataOut_payload_80_31);
  assign _zz_dataOut_payload_80_39 = (_zz_dataOut_payload_80_38 ? _zz_dataOut_payload_80_23 : _zz_dataOut_payload_80_31);
  assign _zz_dataOut_payload_84_3 = (_zz_dataOut_payload_80_38 ? _zz_dataOut_payload_80_31 : _zz_dataOut_payload_80_23);
  assign _zz_dataOut_payload_80_40 = (_zz_dataOut_payload_80_33 < _zz_dataOut_payload_80_37);
  assign _zz_dataOut_payload_80_41 = (_zz_dataOut_payload_80_40 ? _zz_dataOut_payload_80_33 : _zz_dataOut_payload_80_37);
  assign _zz_dataOut_payload_82 = (_zz_dataOut_payload_80_40 ? _zz_dataOut_payload_80_37 : _zz_dataOut_payload_80_33);
  assign _zz_dataOut_payload_80_42 = (_zz_dataOut_payload_80_35 < _zz_dataOut_payload_80_39);
  assign _zz_dataOut_payload_80_43 = (_zz_dataOut_payload_80_42 ? _zz_dataOut_payload_80_35 : _zz_dataOut_payload_80_39);
  assign _zz_dataOut_payload_82_1 = (_zz_dataOut_payload_80_42 ? _zz_dataOut_payload_80_39 : _zz_dataOut_payload_80_35);
  assign _zz_dataOut_payload_80_44 = (_zz_dataOut_payload_80_41 < _zz_dataOut_payload_80_43);
  assign _zz_dataOut_payload_82_2 = (_zz_dataOut_payload_82 < _zz_dataOut_payload_82_1);
  assign _zz_dataOut_payload_84_4 = (_zz_dataOut_payload_84 < _zz_dataOut_payload_84_2);
  assign _zz_dataOut_payload_84_5 = (_zz_dataOut_payload_84_4 ? _zz_dataOut_payload_84 : _zz_dataOut_payload_84_2);
  assign _zz_dataOut_payload_86 = (_zz_dataOut_payload_84_4 ? _zz_dataOut_payload_84_2 : _zz_dataOut_payload_84);
  assign _zz_dataOut_payload_84_6 = (_zz_dataOut_payload_84_1 < _zz_dataOut_payload_84_3);
  assign _zz_dataOut_payload_84_7 = (_zz_dataOut_payload_84_6 ? _zz_dataOut_payload_84_1 : _zz_dataOut_payload_84_3);
  assign _zz_dataOut_payload_86_1 = (_zz_dataOut_payload_84_6 ? _zz_dataOut_payload_84_3 : _zz_dataOut_payload_84_1);
  assign _zz_dataOut_payload_84_8 = (_zz_dataOut_payload_84_5 < _zz_dataOut_payload_84_7);
  assign _zz_dataOut_payload_86_2 = (_zz_dataOut_payload_86 < _zz_dataOut_payload_86_1);
  assign _zz_dataOut_payload_88_8 = (_zz_dataOut_payload_88 < _zz_dataOut_payload_88_4);
  assign _zz_dataOut_payload_88_9 = (_zz_dataOut_payload_88_8 ? _zz_dataOut_payload_88 : _zz_dataOut_payload_88_4);
  assign _zz_dataOut_payload_92 = (_zz_dataOut_payload_88_8 ? _zz_dataOut_payload_88_4 : _zz_dataOut_payload_88);
  assign _zz_dataOut_payload_88_10 = (_zz_dataOut_payload_88_1 < _zz_dataOut_payload_88_5);
  assign _zz_dataOut_payload_88_11 = (_zz_dataOut_payload_88_10 ? _zz_dataOut_payload_88_1 : _zz_dataOut_payload_88_5);
  assign _zz_dataOut_payload_92_1 = (_zz_dataOut_payload_88_10 ? _zz_dataOut_payload_88_5 : _zz_dataOut_payload_88_1);
  assign _zz_dataOut_payload_88_12 = (_zz_dataOut_payload_88_2 < _zz_dataOut_payload_88_6);
  assign _zz_dataOut_payload_88_13 = (_zz_dataOut_payload_88_12 ? _zz_dataOut_payload_88_2 : _zz_dataOut_payload_88_6);
  assign _zz_dataOut_payload_92_2 = (_zz_dataOut_payload_88_12 ? _zz_dataOut_payload_88_6 : _zz_dataOut_payload_88_2);
  assign _zz_dataOut_payload_88_14 = (_zz_dataOut_payload_88_3 < _zz_dataOut_payload_88_7);
  assign _zz_dataOut_payload_88_15 = (_zz_dataOut_payload_88_14 ? _zz_dataOut_payload_88_3 : _zz_dataOut_payload_88_7);
  assign _zz_dataOut_payload_92_3 = (_zz_dataOut_payload_88_14 ? _zz_dataOut_payload_88_7 : _zz_dataOut_payload_88_3);
  assign _zz_dataOut_payload_88_16 = (_zz_dataOut_payload_88_9 < _zz_dataOut_payload_88_13);
  assign _zz_dataOut_payload_88_17 = (_zz_dataOut_payload_88_16 ? _zz_dataOut_payload_88_9 : _zz_dataOut_payload_88_13);
  assign _zz_dataOut_payload_90 = (_zz_dataOut_payload_88_16 ? _zz_dataOut_payload_88_13 : _zz_dataOut_payload_88_9);
  assign _zz_dataOut_payload_88_18 = (_zz_dataOut_payload_88_11 < _zz_dataOut_payload_88_15);
  assign _zz_dataOut_payload_88_19 = (_zz_dataOut_payload_88_18 ? _zz_dataOut_payload_88_11 : _zz_dataOut_payload_88_15);
  assign _zz_dataOut_payload_90_1 = (_zz_dataOut_payload_88_18 ? _zz_dataOut_payload_88_15 : _zz_dataOut_payload_88_11);
  assign _zz_dataOut_payload_88_20 = (_zz_dataOut_payload_88_17 < _zz_dataOut_payload_88_19);
  assign _zz_dataOut_payload_90_2 = (_zz_dataOut_payload_90 < _zz_dataOut_payload_90_1);
  assign _zz_dataOut_payload_92_4 = (_zz_dataOut_payload_92 < _zz_dataOut_payload_92_2);
  assign _zz_dataOut_payload_92_5 = (_zz_dataOut_payload_92_4 ? _zz_dataOut_payload_92 : _zz_dataOut_payload_92_2);
  assign _zz_dataOut_payload_94 = (_zz_dataOut_payload_92_4 ? _zz_dataOut_payload_92_2 : _zz_dataOut_payload_92);
  assign _zz_dataOut_payload_92_6 = (_zz_dataOut_payload_92_1 < _zz_dataOut_payload_92_3);
  assign _zz_dataOut_payload_92_7 = (_zz_dataOut_payload_92_6 ? _zz_dataOut_payload_92_1 : _zz_dataOut_payload_92_3);
  assign _zz_dataOut_payload_94_1 = (_zz_dataOut_payload_92_6 ? _zz_dataOut_payload_92_3 : _zz_dataOut_payload_92_1);
  assign _zz_dataOut_payload_92_8 = (_zz_dataOut_payload_92_5 < _zz_dataOut_payload_92_7);
  assign _zz_dataOut_payload_94_2 = (_zz_dataOut_payload_94 < _zz_dataOut_payload_94_1);
  assign _zz_dataOut_payload_96_32 = (_zz_dataOut_payload_96 < _zz_dataOut_payload_96_16);
  assign _zz_dataOut_payload_96_33 = (_zz_dataOut_payload_96_32 ? _zz_dataOut_payload_96 : _zz_dataOut_payload_96_16);
  assign _zz_dataOut_payload_112 = (_zz_dataOut_payload_96_32 ? _zz_dataOut_payload_96_16 : _zz_dataOut_payload_96);
  assign _zz_dataOut_payload_96_34 = (_zz_dataOut_payload_96_1 < _zz_dataOut_payload_96_17);
  assign _zz_dataOut_payload_96_35 = (_zz_dataOut_payload_96_34 ? _zz_dataOut_payload_96_1 : _zz_dataOut_payload_96_17);
  assign _zz_dataOut_payload_112_1 = (_zz_dataOut_payload_96_34 ? _zz_dataOut_payload_96_17 : _zz_dataOut_payload_96_1);
  assign _zz_dataOut_payload_96_36 = (_zz_dataOut_payload_96_2 < _zz_dataOut_payload_96_18);
  assign _zz_dataOut_payload_96_37 = (_zz_dataOut_payload_96_36 ? _zz_dataOut_payload_96_2 : _zz_dataOut_payload_96_18);
  assign _zz_dataOut_payload_112_2 = (_zz_dataOut_payload_96_36 ? _zz_dataOut_payload_96_18 : _zz_dataOut_payload_96_2);
  assign _zz_dataOut_payload_96_38 = (_zz_dataOut_payload_96_3 < _zz_dataOut_payload_96_19);
  assign _zz_dataOut_payload_96_39 = (_zz_dataOut_payload_96_38 ? _zz_dataOut_payload_96_3 : _zz_dataOut_payload_96_19);
  assign _zz_dataOut_payload_112_3 = (_zz_dataOut_payload_96_38 ? _zz_dataOut_payload_96_19 : _zz_dataOut_payload_96_3);
  assign _zz_dataOut_payload_96_40 = (_zz_dataOut_payload_96_4 < _zz_dataOut_payload_96_20);
  assign _zz_dataOut_payload_96_41 = (_zz_dataOut_payload_96_40 ? _zz_dataOut_payload_96_4 : _zz_dataOut_payload_96_20);
  assign _zz_dataOut_payload_112_4 = (_zz_dataOut_payload_96_40 ? _zz_dataOut_payload_96_20 : _zz_dataOut_payload_96_4);
  assign _zz_dataOut_payload_96_42 = (_zz_dataOut_payload_96_5 < _zz_dataOut_payload_96_21);
  assign _zz_dataOut_payload_96_43 = (_zz_dataOut_payload_96_42 ? _zz_dataOut_payload_96_5 : _zz_dataOut_payload_96_21);
  assign _zz_dataOut_payload_112_5 = (_zz_dataOut_payload_96_42 ? _zz_dataOut_payload_96_21 : _zz_dataOut_payload_96_5);
  assign _zz_dataOut_payload_96_44 = (_zz_dataOut_payload_96_6 < _zz_dataOut_payload_96_22);
  assign _zz_dataOut_payload_96_45 = (_zz_dataOut_payload_96_44 ? _zz_dataOut_payload_96_6 : _zz_dataOut_payload_96_22);
  assign _zz_dataOut_payload_112_6 = (_zz_dataOut_payload_96_44 ? _zz_dataOut_payload_96_22 : _zz_dataOut_payload_96_6);
  assign _zz_dataOut_payload_96_46 = (_zz_dataOut_payload_96_7 < _zz_dataOut_payload_96_23);
  assign _zz_dataOut_payload_96_47 = (_zz_dataOut_payload_96_46 ? _zz_dataOut_payload_96_7 : _zz_dataOut_payload_96_23);
  assign _zz_dataOut_payload_112_7 = (_zz_dataOut_payload_96_46 ? _zz_dataOut_payload_96_23 : _zz_dataOut_payload_96_7);
  assign _zz_dataOut_payload_96_48 = (_zz_dataOut_payload_96_8 < _zz_dataOut_payload_96_24);
  assign _zz_dataOut_payload_96_49 = (_zz_dataOut_payload_96_48 ? _zz_dataOut_payload_96_8 : _zz_dataOut_payload_96_24);
  assign _zz_dataOut_payload_112_8 = (_zz_dataOut_payload_96_48 ? _zz_dataOut_payload_96_24 : _zz_dataOut_payload_96_8);
  assign _zz_dataOut_payload_96_50 = (_zz_dataOut_payload_96_9 < _zz_dataOut_payload_96_25);
  assign _zz_dataOut_payload_96_51 = (_zz_dataOut_payload_96_50 ? _zz_dataOut_payload_96_9 : _zz_dataOut_payload_96_25);
  assign _zz_dataOut_payload_112_9 = (_zz_dataOut_payload_96_50 ? _zz_dataOut_payload_96_25 : _zz_dataOut_payload_96_9);
  assign _zz_dataOut_payload_96_52 = (_zz_dataOut_payload_96_10 < _zz_dataOut_payload_96_26);
  assign _zz_dataOut_payload_96_53 = (_zz_dataOut_payload_96_52 ? _zz_dataOut_payload_96_10 : _zz_dataOut_payload_96_26);
  assign _zz_dataOut_payload_112_10 = (_zz_dataOut_payload_96_52 ? _zz_dataOut_payload_96_26 : _zz_dataOut_payload_96_10);
  assign _zz_dataOut_payload_96_54 = (_zz_dataOut_payload_96_11 < _zz_dataOut_payload_96_27);
  assign _zz_dataOut_payload_96_55 = (_zz_dataOut_payload_96_54 ? _zz_dataOut_payload_96_11 : _zz_dataOut_payload_96_27);
  assign _zz_dataOut_payload_112_11 = (_zz_dataOut_payload_96_54 ? _zz_dataOut_payload_96_27 : _zz_dataOut_payload_96_11);
  assign _zz_dataOut_payload_96_56 = (_zz_dataOut_payload_96_12 < _zz_dataOut_payload_96_28);
  assign _zz_dataOut_payload_96_57 = (_zz_dataOut_payload_96_56 ? _zz_dataOut_payload_96_12 : _zz_dataOut_payload_96_28);
  assign _zz_dataOut_payload_112_12 = (_zz_dataOut_payload_96_56 ? _zz_dataOut_payload_96_28 : _zz_dataOut_payload_96_12);
  assign _zz_dataOut_payload_96_58 = (_zz_dataOut_payload_96_13 < _zz_dataOut_payload_96_29);
  assign _zz_dataOut_payload_96_59 = (_zz_dataOut_payload_96_58 ? _zz_dataOut_payload_96_13 : _zz_dataOut_payload_96_29);
  assign _zz_dataOut_payload_112_13 = (_zz_dataOut_payload_96_58 ? _zz_dataOut_payload_96_29 : _zz_dataOut_payload_96_13);
  assign _zz_dataOut_payload_96_60 = (_zz_dataOut_payload_96_14 < _zz_dataOut_payload_96_30);
  assign _zz_dataOut_payload_96_61 = (_zz_dataOut_payload_96_60 ? _zz_dataOut_payload_96_14 : _zz_dataOut_payload_96_30);
  assign _zz_dataOut_payload_112_14 = (_zz_dataOut_payload_96_60 ? _zz_dataOut_payload_96_30 : _zz_dataOut_payload_96_14);
  assign _zz_dataOut_payload_96_62 = (_zz_dataOut_payload_96_15 < _zz_dataOut_payload_96_31);
  assign _zz_dataOut_payload_96_63 = (_zz_dataOut_payload_96_62 ? _zz_dataOut_payload_96_15 : _zz_dataOut_payload_96_31);
  assign _zz_dataOut_payload_112_15 = (_zz_dataOut_payload_96_62 ? _zz_dataOut_payload_96_31 : _zz_dataOut_payload_96_15);
  assign _zz_dataOut_payload_96_64 = (_zz_dataOut_payload_96_33 < _zz_dataOut_payload_96_49);
  assign _zz_dataOut_payload_96_65 = (_zz_dataOut_payload_96_64 ? _zz_dataOut_payload_96_33 : _zz_dataOut_payload_96_49);
  assign _zz_dataOut_payload_104 = (_zz_dataOut_payload_96_64 ? _zz_dataOut_payload_96_49 : _zz_dataOut_payload_96_33);
  assign _zz_dataOut_payload_96_66 = (_zz_dataOut_payload_96_35 < _zz_dataOut_payload_96_51);
  assign _zz_dataOut_payload_96_67 = (_zz_dataOut_payload_96_66 ? _zz_dataOut_payload_96_35 : _zz_dataOut_payload_96_51);
  assign _zz_dataOut_payload_104_1 = (_zz_dataOut_payload_96_66 ? _zz_dataOut_payload_96_51 : _zz_dataOut_payload_96_35);
  assign _zz_dataOut_payload_96_68 = (_zz_dataOut_payload_96_37 < _zz_dataOut_payload_96_53);
  assign _zz_dataOut_payload_96_69 = (_zz_dataOut_payload_96_68 ? _zz_dataOut_payload_96_37 : _zz_dataOut_payload_96_53);
  assign _zz_dataOut_payload_104_2 = (_zz_dataOut_payload_96_68 ? _zz_dataOut_payload_96_53 : _zz_dataOut_payload_96_37);
  assign _zz_dataOut_payload_96_70 = (_zz_dataOut_payload_96_39 < _zz_dataOut_payload_96_55);
  assign _zz_dataOut_payload_96_71 = (_zz_dataOut_payload_96_70 ? _zz_dataOut_payload_96_39 : _zz_dataOut_payload_96_55);
  assign _zz_dataOut_payload_104_3 = (_zz_dataOut_payload_96_70 ? _zz_dataOut_payload_96_55 : _zz_dataOut_payload_96_39);
  assign _zz_dataOut_payload_96_72 = (_zz_dataOut_payload_96_41 < _zz_dataOut_payload_96_57);
  assign _zz_dataOut_payload_96_73 = (_zz_dataOut_payload_96_72 ? _zz_dataOut_payload_96_41 : _zz_dataOut_payload_96_57);
  assign _zz_dataOut_payload_104_4 = (_zz_dataOut_payload_96_72 ? _zz_dataOut_payload_96_57 : _zz_dataOut_payload_96_41);
  assign _zz_dataOut_payload_96_74 = (_zz_dataOut_payload_96_43 < _zz_dataOut_payload_96_59);
  assign _zz_dataOut_payload_96_75 = (_zz_dataOut_payload_96_74 ? _zz_dataOut_payload_96_43 : _zz_dataOut_payload_96_59);
  assign _zz_dataOut_payload_104_5 = (_zz_dataOut_payload_96_74 ? _zz_dataOut_payload_96_59 : _zz_dataOut_payload_96_43);
  assign _zz_dataOut_payload_96_76 = (_zz_dataOut_payload_96_45 < _zz_dataOut_payload_96_61);
  assign _zz_dataOut_payload_96_77 = (_zz_dataOut_payload_96_76 ? _zz_dataOut_payload_96_45 : _zz_dataOut_payload_96_61);
  assign _zz_dataOut_payload_104_6 = (_zz_dataOut_payload_96_76 ? _zz_dataOut_payload_96_61 : _zz_dataOut_payload_96_45);
  assign _zz_dataOut_payload_96_78 = (_zz_dataOut_payload_96_47 < _zz_dataOut_payload_96_63);
  assign _zz_dataOut_payload_96_79 = (_zz_dataOut_payload_96_78 ? _zz_dataOut_payload_96_47 : _zz_dataOut_payload_96_63);
  assign _zz_dataOut_payload_104_7 = (_zz_dataOut_payload_96_78 ? _zz_dataOut_payload_96_63 : _zz_dataOut_payload_96_47);
  assign _zz_dataOut_payload_96_80 = (_zz_dataOut_payload_96_65 < _zz_dataOut_payload_96_73);
  assign _zz_dataOut_payload_96_81 = (_zz_dataOut_payload_96_80 ? _zz_dataOut_payload_96_65 : _zz_dataOut_payload_96_73);
  assign _zz_dataOut_payload_100 = (_zz_dataOut_payload_96_80 ? _zz_dataOut_payload_96_73 : _zz_dataOut_payload_96_65);
  assign _zz_dataOut_payload_96_82 = (_zz_dataOut_payload_96_67 < _zz_dataOut_payload_96_75);
  assign _zz_dataOut_payload_96_83 = (_zz_dataOut_payload_96_82 ? _zz_dataOut_payload_96_67 : _zz_dataOut_payload_96_75);
  assign _zz_dataOut_payload_100_1 = (_zz_dataOut_payload_96_82 ? _zz_dataOut_payload_96_75 : _zz_dataOut_payload_96_67);
  assign _zz_dataOut_payload_96_84 = (_zz_dataOut_payload_96_69 < _zz_dataOut_payload_96_77);
  assign _zz_dataOut_payload_96_85 = (_zz_dataOut_payload_96_84 ? _zz_dataOut_payload_96_69 : _zz_dataOut_payload_96_77);
  assign _zz_dataOut_payload_100_2 = (_zz_dataOut_payload_96_84 ? _zz_dataOut_payload_96_77 : _zz_dataOut_payload_96_69);
  assign _zz_dataOut_payload_96_86 = (_zz_dataOut_payload_96_71 < _zz_dataOut_payload_96_79);
  assign _zz_dataOut_payload_96_87 = (_zz_dataOut_payload_96_86 ? _zz_dataOut_payload_96_71 : _zz_dataOut_payload_96_79);
  assign _zz_dataOut_payload_100_3 = (_zz_dataOut_payload_96_86 ? _zz_dataOut_payload_96_79 : _zz_dataOut_payload_96_71);
  assign _zz_dataOut_payload_96_88 = (_zz_dataOut_payload_96_81 < _zz_dataOut_payload_96_85);
  assign _zz_dataOut_payload_96_89 = (_zz_dataOut_payload_96_88 ? _zz_dataOut_payload_96_81 : _zz_dataOut_payload_96_85);
  assign _zz_dataOut_payload_98 = (_zz_dataOut_payload_96_88 ? _zz_dataOut_payload_96_85 : _zz_dataOut_payload_96_81);
  assign _zz_dataOut_payload_96_90 = (_zz_dataOut_payload_96_83 < _zz_dataOut_payload_96_87);
  assign _zz_dataOut_payload_96_91 = (_zz_dataOut_payload_96_90 ? _zz_dataOut_payload_96_83 : _zz_dataOut_payload_96_87);
  assign _zz_dataOut_payload_98_1 = (_zz_dataOut_payload_96_90 ? _zz_dataOut_payload_96_87 : _zz_dataOut_payload_96_83);
  assign _zz_dataOut_payload_96_92 = (_zz_dataOut_payload_96_89 < _zz_dataOut_payload_96_91);
  assign _zz_dataOut_payload_98_2 = (_zz_dataOut_payload_98 < _zz_dataOut_payload_98_1);
  assign _zz_dataOut_payload_100_4 = (_zz_dataOut_payload_100 < _zz_dataOut_payload_100_2);
  assign _zz_dataOut_payload_100_5 = (_zz_dataOut_payload_100_4 ? _zz_dataOut_payload_100 : _zz_dataOut_payload_100_2);
  assign _zz_dataOut_payload_102 = (_zz_dataOut_payload_100_4 ? _zz_dataOut_payload_100_2 : _zz_dataOut_payload_100);
  assign _zz_dataOut_payload_100_6 = (_zz_dataOut_payload_100_1 < _zz_dataOut_payload_100_3);
  assign _zz_dataOut_payload_100_7 = (_zz_dataOut_payload_100_6 ? _zz_dataOut_payload_100_1 : _zz_dataOut_payload_100_3);
  assign _zz_dataOut_payload_102_1 = (_zz_dataOut_payload_100_6 ? _zz_dataOut_payload_100_3 : _zz_dataOut_payload_100_1);
  assign _zz_dataOut_payload_100_8 = (_zz_dataOut_payload_100_5 < _zz_dataOut_payload_100_7);
  assign _zz_dataOut_payload_102_2 = (_zz_dataOut_payload_102 < _zz_dataOut_payload_102_1);
  assign _zz_dataOut_payload_104_8 = (_zz_dataOut_payload_104 < _zz_dataOut_payload_104_4);
  assign _zz_dataOut_payload_104_9 = (_zz_dataOut_payload_104_8 ? _zz_dataOut_payload_104 : _zz_dataOut_payload_104_4);
  assign _zz_dataOut_payload_108 = (_zz_dataOut_payload_104_8 ? _zz_dataOut_payload_104_4 : _zz_dataOut_payload_104);
  assign _zz_dataOut_payload_104_10 = (_zz_dataOut_payload_104_1 < _zz_dataOut_payload_104_5);
  assign _zz_dataOut_payload_104_11 = (_zz_dataOut_payload_104_10 ? _zz_dataOut_payload_104_1 : _zz_dataOut_payload_104_5);
  assign _zz_dataOut_payload_108_1 = (_zz_dataOut_payload_104_10 ? _zz_dataOut_payload_104_5 : _zz_dataOut_payload_104_1);
  assign _zz_dataOut_payload_104_12 = (_zz_dataOut_payload_104_2 < _zz_dataOut_payload_104_6);
  assign _zz_dataOut_payload_104_13 = (_zz_dataOut_payload_104_12 ? _zz_dataOut_payload_104_2 : _zz_dataOut_payload_104_6);
  assign _zz_dataOut_payload_108_2 = (_zz_dataOut_payload_104_12 ? _zz_dataOut_payload_104_6 : _zz_dataOut_payload_104_2);
  assign _zz_dataOut_payload_104_14 = (_zz_dataOut_payload_104_3 < _zz_dataOut_payload_104_7);
  assign _zz_dataOut_payload_104_15 = (_zz_dataOut_payload_104_14 ? _zz_dataOut_payload_104_3 : _zz_dataOut_payload_104_7);
  assign _zz_dataOut_payload_108_3 = (_zz_dataOut_payload_104_14 ? _zz_dataOut_payload_104_7 : _zz_dataOut_payload_104_3);
  assign _zz_dataOut_payload_104_16 = (_zz_dataOut_payload_104_9 < _zz_dataOut_payload_104_13);
  assign _zz_dataOut_payload_104_17 = (_zz_dataOut_payload_104_16 ? _zz_dataOut_payload_104_9 : _zz_dataOut_payload_104_13);
  assign _zz_dataOut_payload_106 = (_zz_dataOut_payload_104_16 ? _zz_dataOut_payload_104_13 : _zz_dataOut_payload_104_9);
  assign _zz_dataOut_payload_104_18 = (_zz_dataOut_payload_104_11 < _zz_dataOut_payload_104_15);
  assign _zz_dataOut_payload_104_19 = (_zz_dataOut_payload_104_18 ? _zz_dataOut_payload_104_11 : _zz_dataOut_payload_104_15);
  assign _zz_dataOut_payload_106_1 = (_zz_dataOut_payload_104_18 ? _zz_dataOut_payload_104_15 : _zz_dataOut_payload_104_11);
  assign _zz_dataOut_payload_104_20 = (_zz_dataOut_payload_104_17 < _zz_dataOut_payload_104_19);
  assign _zz_dataOut_payload_106_2 = (_zz_dataOut_payload_106 < _zz_dataOut_payload_106_1);
  assign _zz_dataOut_payload_108_4 = (_zz_dataOut_payload_108 < _zz_dataOut_payload_108_2);
  assign _zz_dataOut_payload_108_5 = (_zz_dataOut_payload_108_4 ? _zz_dataOut_payload_108 : _zz_dataOut_payload_108_2);
  assign _zz_dataOut_payload_110 = (_zz_dataOut_payload_108_4 ? _zz_dataOut_payload_108_2 : _zz_dataOut_payload_108);
  assign _zz_dataOut_payload_108_6 = (_zz_dataOut_payload_108_1 < _zz_dataOut_payload_108_3);
  assign _zz_dataOut_payload_108_7 = (_zz_dataOut_payload_108_6 ? _zz_dataOut_payload_108_1 : _zz_dataOut_payload_108_3);
  assign _zz_dataOut_payload_110_1 = (_zz_dataOut_payload_108_6 ? _zz_dataOut_payload_108_3 : _zz_dataOut_payload_108_1);
  assign _zz_dataOut_payload_108_8 = (_zz_dataOut_payload_108_5 < _zz_dataOut_payload_108_7);
  assign _zz_dataOut_payload_110_2 = (_zz_dataOut_payload_110 < _zz_dataOut_payload_110_1);
  assign _zz_dataOut_payload_112_16 = (_zz_dataOut_payload_112 < _zz_dataOut_payload_112_8);
  assign _zz_dataOut_payload_112_17 = (_zz_dataOut_payload_112_16 ? _zz_dataOut_payload_112 : _zz_dataOut_payload_112_8);
  assign _zz_dataOut_payload_120 = (_zz_dataOut_payload_112_16 ? _zz_dataOut_payload_112_8 : _zz_dataOut_payload_112);
  assign _zz_dataOut_payload_112_18 = (_zz_dataOut_payload_112_1 < _zz_dataOut_payload_112_9);
  assign _zz_dataOut_payload_112_19 = (_zz_dataOut_payload_112_18 ? _zz_dataOut_payload_112_1 : _zz_dataOut_payload_112_9);
  assign _zz_dataOut_payload_120_1 = (_zz_dataOut_payload_112_18 ? _zz_dataOut_payload_112_9 : _zz_dataOut_payload_112_1);
  assign _zz_dataOut_payload_112_20 = (_zz_dataOut_payload_112_2 < _zz_dataOut_payload_112_10);
  assign _zz_dataOut_payload_112_21 = (_zz_dataOut_payload_112_20 ? _zz_dataOut_payload_112_2 : _zz_dataOut_payload_112_10);
  assign _zz_dataOut_payload_120_2 = (_zz_dataOut_payload_112_20 ? _zz_dataOut_payload_112_10 : _zz_dataOut_payload_112_2);
  assign _zz_dataOut_payload_112_22 = (_zz_dataOut_payload_112_3 < _zz_dataOut_payload_112_11);
  assign _zz_dataOut_payload_112_23 = (_zz_dataOut_payload_112_22 ? _zz_dataOut_payload_112_3 : _zz_dataOut_payload_112_11);
  assign _zz_dataOut_payload_120_3 = (_zz_dataOut_payload_112_22 ? _zz_dataOut_payload_112_11 : _zz_dataOut_payload_112_3);
  assign _zz_dataOut_payload_112_24 = (_zz_dataOut_payload_112_4 < _zz_dataOut_payload_112_12);
  assign _zz_dataOut_payload_112_25 = (_zz_dataOut_payload_112_24 ? _zz_dataOut_payload_112_4 : _zz_dataOut_payload_112_12);
  assign _zz_dataOut_payload_120_4 = (_zz_dataOut_payload_112_24 ? _zz_dataOut_payload_112_12 : _zz_dataOut_payload_112_4);
  assign _zz_dataOut_payload_112_26 = (_zz_dataOut_payload_112_5 < _zz_dataOut_payload_112_13);
  assign _zz_dataOut_payload_112_27 = (_zz_dataOut_payload_112_26 ? _zz_dataOut_payload_112_5 : _zz_dataOut_payload_112_13);
  assign _zz_dataOut_payload_120_5 = (_zz_dataOut_payload_112_26 ? _zz_dataOut_payload_112_13 : _zz_dataOut_payload_112_5);
  assign _zz_dataOut_payload_112_28 = (_zz_dataOut_payload_112_6 < _zz_dataOut_payload_112_14);
  assign _zz_dataOut_payload_112_29 = (_zz_dataOut_payload_112_28 ? _zz_dataOut_payload_112_6 : _zz_dataOut_payload_112_14);
  assign _zz_dataOut_payload_120_6 = (_zz_dataOut_payload_112_28 ? _zz_dataOut_payload_112_14 : _zz_dataOut_payload_112_6);
  assign _zz_dataOut_payload_112_30 = (_zz_dataOut_payload_112_7 < _zz_dataOut_payload_112_15);
  assign _zz_dataOut_payload_112_31 = (_zz_dataOut_payload_112_30 ? _zz_dataOut_payload_112_7 : _zz_dataOut_payload_112_15);
  assign _zz_dataOut_payload_120_7 = (_zz_dataOut_payload_112_30 ? _zz_dataOut_payload_112_15 : _zz_dataOut_payload_112_7);
  assign _zz_dataOut_payload_112_32 = (_zz_dataOut_payload_112_17 < _zz_dataOut_payload_112_25);
  assign _zz_dataOut_payload_112_33 = (_zz_dataOut_payload_112_32 ? _zz_dataOut_payload_112_17 : _zz_dataOut_payload_112_25);
  assign _zz_dataOut_payload_116 = (_zz_dataOut_payload_112_32 ? _zz_dataOut_payload_112_25 : _zz_dataOut_payload_112_17);
  assign _zz_dataOut_payload_112_34 = (_zz_dataOut_payload_112_19 < _zz_dataOut_payload_112_27);
  assign _zz_dataOut_payload_112_35 = (_zz_dataOut_payload_112_34 ? _zz_dataOut_payload_112_19 : _zz_dataOut_payload_112_27);
  assign _zz_dataOut_payload_116_1 = (_zz_dataOut_payload_112_34 ? _zz_dataOut_payload_112_27 : _zz_dataOut_payload_112_19);
  assign _zz_dataOut_payload_112_36 = (_zz_dataOut_payload_112_21 < _zz_dataOut_payload_112_29);
  assign _zz_dataOut_payload_112_37 = (_zz_dataOut_payload_112_36 ? _zz_dataOut_payload_112_21 : _zz_dataOut_payload_112_29);
  assign _zz_dataOut_payload_116_2 = (_zz_dataOut_payload_112_36 ? _zz_dataOut_payload_112_29 : _zz_dataOut_payload_112_21);
  assign _zz_dataOut_payload_112_38 = (_zz_dataOut_payload_112_23 < _zz_dataOut_payload_112_31);
  assign _zz_dataOut_payload_112_39 = (_zz_dataOut_payload_112_38 ? _zz_dataOut_payload_112_23 : _zz_dataOut_payload_112_31);
  assign _zz_dataOut_payload_116_3 = (_zz_dataOut_payload_112_38 ? _zz_dataOut_payload_112_31 : _zz_dataOut_payload_112_23);
  assign _zz_dataOut_payload_112_40 = (_zz_dataOut_payload_112_33 < _zz_dataOut_payload_112_37);
  assign _zz_dataOut_payload_112_41 = (_zz_dataOut_payload_112_40 ? _zz_dataOut_payload_112_33 : _zz_dataOut_payload_112_37);
  assign _zz_dataOut_payload_114 = (_zz_dataOut_payload_112_40 ? _zz_dataOut_payload_112_37 : _zz_dataOut_payload_112_33);
  assign _zz_dataOut_payload_112_42 = (_zz_dataOut_payload_112_35 < _zz_dataOut_payload_112_39);
  assign _zz_dataOut_payload_112_43 = (_zz_dataOut_payload_112_42 ? _zz_dataOut_payload_112_35 : _zz_dataOut_payload_112_39);
  assign _zz_dataOut_payload_114_1 = (_zz_dataOut_payload_112_42 ? _zz_dataOut_payload_112_39 : _zz_dataOut_payload_112_35);
  assign _zz_dataOut_payload_112_44 = (_zz_dataOut_payload_112_41 < _zz_dataOut_payload_112_43);
  assign _zz_dataOut_payload_114_2 = (_zz_dataOut_payload_114 < _zz_dataOut_payload_114_1);
  assign _zz_dataOut_payload_116_4 = (_zz_dataOut_payload_116 < _zz_dataOut_payload_116_2);
  assign _zz_dataOut_payload_116_5 = (_zz_dataOut_payload_116_4 ? _zz_dataOut_payload_116 : _zz_dataOut_payload_116_2);
  assign _zz_dataOut_payload_118 = (_zz_dataOut_payload_116_4 ? _zz_dataOut_payload_116_2 : _zz_dataOut_payload_116);
  assign _zz_dataOut_payload_116_6 = (_zz_dataOut_payload_116_1 < _zz_dataOut_payload_116_3);
  assign _zz_dataOut_payload_116_7 = (_zz_dataOut_payload_116_6 ? _zz_dataOut_payload_116_1 : _zz_dataOut_payload_116_3);
  assign _zz_dataOut_payload_118_1 = (_zz_dataOut_payload_116_6 ? _zz_dataOut_payload_116_3 : _zz_dataOut_payload_116_1);
  assign _zz_dataOut_payload_116_8 = (_zz_dataOut_payload_116_5 < _zz_dataOut_payload_116_7);
  assign _zz_dataOut_payload_118_2 = (_zz_dataOut_payload_118 < _zz_dataOut_payload_118_1);
  assign _zz_dataOut_payload_120_8 = (_zz_dataOut_payload_120 < _zz_dataOut_payload_120_4);
  assign _zz_dataOut_payload_120_9 = (_zz_dataOut_payload_120_8 ? _zz_dataOut_payload_120 : _zz_dataOut_payload_120_4);
  assign _zz_dataOut_payload_124 = (_zz_dataOut_payload_120_8 ? _zz_dataOut_payload_120_4 : _zz_dataOut_payload_120);
  assign _zz_dataOut_payload_120_10 = (_zz_dataOut_payload_120_1 < _zz_dataOut_payload_120_5);
  assign _zz_dataOut_payload_120_11 = (_zz_dataOut_payload_120_10 ? _zz_dataOut_payload_120_1 : _zz_dataOut_payload_120_5);
  assign _zz_dataOut_payload_124_1 = (_zz_dataOut_payload_120_10 ? _zz_dataOut_payload_120_5 : _zz_dataOut_payload_120_1);
  assign _zz_dataOut_payload_120_12 = (_zz_dataOut_payload_120_2 < _zz_dataOut_payload_120_6);
  assign _zz_dataOut_payload_120_13 = (_zz_dataOut_payload_120_12 ? _zz_dataOut_payload_120_2 : _zz_dataOut_payload_120_6);
  assign _zz_dataOut_payload_124_2 = (_zz_dataOut_payload_120_12 ? _zz_dataOut_payload_120_6 : _zz_dataOut_payload_120_2);
  assign _zz_dataOut_payload_120_14 = (_zz_dataOut_payload_120_3 < _zz_dataOut_payload_120_7);
  assign _zz_dataOut_payload_120_15 = (_zz_dataOut_payload_120_14 ? _zz_dataOut_payload_120_3 : _zz_dataOut_payload_120_7);
  assign _zz_dataOut_payload_124_3 = (_zz_dataOut_payload_120_14 ? _zz_dataOut_payload_120_7 : _zz_dataOut_payload_120_3);
  assign _zz_dataOut_payload_120_16 = (_zz_dataOut_payload_120_9 < _zz_dataOut_payload_120_13);
  assign _zz_dataOut_payload_120_17 = (_zz_dataOut_payload_120_16 ? _zz_dataOut_payload_120_9 : _zz_dataOut_payload_120_13);
  assign _zz_dataOut_payload_122 = (_zz_dataOut_payload_120_16 ? _zz_dataOut_payload_120_13 : _zz_dataOut_payload_120_9);
  assign _zz_dataOut_payload_120_18 = (_zz_dataOut_payload_120_11 < _zz_dataOut_payload_120_15);
  assign _zz_dataOut_payload_120_19 = (_zz_dataOut_payload_120_18 ? _zz_dataOut_payload_120_11 : _zz_dataOut_payload_120_15);
  assign _zz_dataOut_payload_122_1 = (_zz_dataOut_payload_120_18 ? _zz_dataOut_payload_120_15 : _zz_dataOut_payload_120_11);
  assign _zz_dataOut_payload_120_20 = (_zz_dataOut_payload_120_17 < _zz_dataOut_payload_120_19);
  assign _zz_dataOut_payload_122_2 = (_zz_dataOut_payload_122 < _zz_dataOut_payload_122_1);
  assign _zz_dataOut_payload_124_4 = (_zz_dataOut_payload_124 < _zz_dataOut_payload_124_2);
  assign _zz_dataOut_payload_124_5 = (_zz_dataOut_payload_124_4 ? _zz_dataOut_payload_124 : _zz_dataOut_payload_124_2);
  assign _zz_dataOut_payload_126 = (_zz_dataOut_payload_124_4 ? _zz_dataOut_payload_124_2 : _zz_dataOut_payload_124);
  assign _zz_dataOut_payload_124_6 = (_zz_dataOut_payload_124_1 < _zz_dataOut_payload_124_3);
  assign _zz_dataOut_payload_124_7 = (_zz_dataOut_payload_124_6 ? _zz_dataOut_payload_124_1 : _zz_dataOut_payload_124_3);
  assign _zz_dataOut_payload_126_1 = (_zz_dataOut_payload_124_6 ? _zz_dataOut_payload_124_3 : _zz_dataOut_payload_124_1);
  assign _zz_dataOut_payload_124_8 = (_zz_dataOut_payload_124_5 < _zz_dataOut_payload_124_7);
  assign _zz_dataOut_payload_126_2 = (_zz_dataOut_payload_126 < _zz_dataOut_payload_126_1);
  assign _zz_dataOut_payload_128_128 = (_zz_dataOut_payload_128_127 < _zz_dataOut_payload_128_63);
  assign _zz_dataOut_payload_128_129 = (_zz_dataOut_payload_128_128 ? _zz_dataOut_payload_128_127 : _zz_dataOut_payload_128_63);
  assign _zz_dataOut_payload_192 = (_zz_dataOut_payload_128_128 ? _zz_dataOut_payload_128_63 : _zz_dataOut_payload_128_127);
  assign _zz_dataOut_payload_128_130 = (_zz_dataOut_payload_128_126 < _zz_dataOut_payload_128_62);
  assign _zz_dataOut_payload_128_131 = (_zz_dataOut_payload_128_130 ? _zz_dataOut_payload_128_126 : _zz_dataOut_payload_128_62);
  assign _zz_dataOut_payload_192_1 = (_zz_dataOut_payload_128_130 ? _zz_dataOut_payload_128_62 : _zz_dataOut_payload_128_126);
  assign _zz_dataOut_payload_128_132 = (_zz_dataOut_payload_128_125 < _zz_dataOut_payload_128_61);
  assign _zz_dataOut_payload_128_133 = (_zz_dataOut_payload_128_132 ? _zz_dataOut_payload_128_125 : _zz_dataOut_payload_128_61);
  assign _zz_dataOut_payload_192_2 = (_zz_dataOut_payload_128_132 ? _zz_dataOut_payload_128_61 : _zz_dataOut_payload_128_125);
  assign _zz_dataOut_payload_128_134 = (_zz_dataOut_payload_128_124 < _zz_dataOut_payload_128_60);
  assign _zz_dataOut_payload_128_135 = (_zz_dataOut_payload_128_134 ? _zz_dataOut_payload_128_124 : _zz_dataOut_payload_128_60);
  assign _zz_dataOut_payload_192_3 = (_zz_dataOut_payload_128_134 ? _zz_dataOut_payload_128_60 : _zz_dataOut_payload_128_124);
  assign _zz_dataOut_payload_128_136 = (_zz_dataOut_payload_128_123 < _zz_dataOut_payload_128_59);
  assign _zz_dataOut_payload_128_137 = (_zz_dataOut_payload_128_136 ? _zz_dataOut_payload_128_123 : _zz_dataOut_payload_128_59);
  assign _zz_dataOut_payload_192_4 = (_zz_dataOut_payload_128_136 ? _zz_dataOut_payload_128_59 : _zz_dataOut_payload_128_123);
  assign _zz_dataOut_payload_128_138 = (_zz_dataOut_payload_128_122 < _zz_dataOut_payload_128_58);
  assign _zz_dataOut_payload_128_139 = (_zz_dataOut_payload_128_138 ? _zz_dataOut_payload_128_122 : _zz_dataOut_payload_128_58);
  assign _zz_dataOut_payload_192_5 = (_zz_dataOut_payload_128_138 ? _zz_dataOut_payload_128_58 : _zz_dataOut_payload_128_122);
  assign _zz_dataOut_payload_128_140 = (_zz_dataOut_payload_128_121 < _zz_dataOut_payload_128_57);
  assign _zz_dataOut_payload_128_141 = (_zz_dataOut_payload_128_140 ? _zz_dataOut_payload_128_121 : _zz_dataOut_payload_128_57);
  assign _zz_dataOut_payload_192_6 = (_zz_dataOut_payload_128_140 ? _zz_dataOut_payload_128_57 : _zz_dataOut_payload_128_121);
  assign _zz_dataOut_payload_128_142 = (_zz_dataOut_payload_128_120 < _zz_dataOut_payload_128_56);
  assign _zz_dataOut_payload_128_143 = (_zz_dataOut_payload_128_142 ? _zz_dataOut_payload_128_120 : _zz_dataOut_payload_128_56);
  assign _zz_dataOut_payload_192_7 = (_zz_dataOut_payload_128_142 ? _zz_dataOut_payload_128_56 : _zz_dataOut_payload_128_120);
  assign _zz_dataOut_payload_128_144 = (_zz_dataOut_payload_128_119 < _zz_dataOut_payload_128_55);
  assign _zz_dataOut_payload_128_145 = (_zz_dataOut_payload_128_144 ? _zz_dataOut_payload_128_119 : _zz_dataOut_payload_128_55);
  assign _zz_dataOut_payload_192_8 = (_zz_dataOut_payload_128_144 ? _zz_dataOut_payload_128_55 : _zz_dataOut_payload_128_119);
  assign _zz_dataOut_payload_128_146 = (_zz_dataOut_payload_128_118 < _zz_dataOut_payload_128_54);
  assign _zz_dataOut_payload_128_147 = (_zz_dataOut_payload_128_146 ? _zz_dataOut_payload_128_118 : _zz_dataOut_payload_128_54);
  assign _zz_dataOut_payload_192_9 = (_zz_dataOut_payload_128_146 ? _zz_dataOut_payload_128_54 : _zz_dataOut_payload_128_118);
  assign _zz_dataOut_payload_128_148 = (_zz_dataOut_payload_128_117 < _zz_dataOut_payload_128_53);
  assign _zz_dataOut_payload_128_149 = (_zz_dataOut_payload_128_148 ? _zz_dataOut_payload_128_117 : _zz_dataOut_payload_128_53);
  assign _zz_dataOut_payload_192_10 = (_zz_dataOut_payload_128_148 ? _zz_dataOut_payload_128_53 : _zz_dataOut_payload_128_117);
  assign _zz_dataOut_payload_128_150 = (_zz_dataOut_payload_128_116 < _zz_dataOut_payload_128_52);
  assign _zz_dataOut_payload_128_151 = (_zz_dataOut_payload_128_150 ? _zz_dataOut_payload_128_116 : _zz_dataOut_payload_128_52);
  assign _zz_dataOut_payload_192_11 = (_zz_dataOut_payload_128_150 ? _zz_dataOut_payload_128_52 : _zz_dataOut_payload_128_116);
  assign _zz_dataOut_payload_128_152 = (_zz_dataOut_payload_128_115 < _zz_dataOut_payload_128_51);
  assign _zz_dataOut_payload_128_153 = (_zz_dataOut_payload_128_152 ? _zz_dataOut_payload_128_115 : _zz_dataOut_payload_128_51);
  assign _zz_dataOut_payload_192_12 = (_zz_dataOut_payload_128_152 ? _zz_dataOut_payload_128_51 : _zz_dataOut_payload_128_115);
  assign _zz_dataOut_payload_128_154 = (_zz_dataOut_payload_128_114 < _zz_dataOut_payload_128_50);
  assign _zz_dataOut_payload_128_155 = (_zz_dataOut_payload_128_154 ? _zz_dataOut_payload_128_114 : _zz_dataOut_payload_128_50);
  assign _zz_dataOut_payload_192_13 = (_zz_dataOut_payload_128_154 ? _zz_dataOut_payload_128_50 : _zz_dataOut_payload_128_114);
  assign _zz_dataOut_payload_128_156 = (_zz_dataOut_payload_128_113 < _zz_dataOut_payload_128_49);
  assign _zz_dataOut_payload_128_157 = (_zz_dataOut_payload_128_156 ? _zz_dataOut_payload_128_113 : _zz_dataOut_payload_128_49);
  assign _zz_dataOut_payload_192_14 = (_zz_dataOut_payload_128_156 ? _zz_dataOut_payload_128_49 : _zz_dataOut_payload_128_113);
  assign _zz_dataOut_payload_128_158 = (_zz_dataOut_payload_128_112 < _zz_dataOut_payload_128_48);
  assign _zz_dataOut_payload_128_159 = (_zz_dataOut_payload_128_158 ? _zz_dataOut_payload_128_112 : _zz_dataOut_payload_128_48);
  assign _zz_dataOut_payload_192_15 = (_zz_dataOut_payload_128_158 ? _zz_dataOut_payload_128_48 : _zz_dataOut_payload_128_112);
  assign _zz_dataOut_payload_128_160 = (_zz_dataOut_payload_128_111 < _zz_dataOut_payload_128_47);
  assign _zz_dataOut_payload_128_161 = (_zz_dataOut_payload_128_160 ? _zz_dataOut_payload_128_111 : _zz_dataOut_payload_128_47);
  assign _zz_dataOut_payload_192_16 = (_zz_dataOut_payload_128_160 ? _zz_dataOut_payload_128_47 : _zz_dataOut_payload_128_111);
  assign _zz_dataOut_payload_128_162 = (_zz_dataOut_payload_128_110 < _zz_dataOut_payload_128_46);
  assign _zz_dataOut_payload_128_163 = (_zz_dataOut_payload_128_162 ? _zz_dataOut_payload_128_110 : _zz_dataOut_payload_128_46);
  assign _zz_dataOut_payload_192_17 = (_zz_dataOut_payload_128_162 ? _zz_dataOut_payload_128_46 : _zz_dataOut_payload_128_110);
  assign _zz_dataOut_payload_128_164 = (_zz_dataOut_payload_128_109 < _zz_dataOut_payload_128_45);
  assign _zz_dataOut_payload_128_165 = (_zz_dataOut_payload_128_164 ? _zz_dataOut_payload_128_109 : _zz_dataOut_payload_128_45);
  assign _zz_dataOut_payload_192_18 = (_zz_dataOut_payload_128_164 ? _zz_dataOut_payload_128_45 : _zz_dataOut_payload_128_109);
  assign _zz_dataOut_payload_128_166 = (_zz_dataOut_payload_128_108 < _zz_dataOut_payload_128_44);
  assign _zz_dataOut_payload_128_167 = (_zz_dataOut_payload_128_166 ? _zz_dataOut_payload_128_108 : _zz_dataOut_payload_128_44);
  assign _zz_dataOut_payload_192_19 = (_zz_dataOut_payload_128_166 ? _zz_dataOut_payload_128_44 : _zz_dataOut_payload_128_108);
  assign _zz_dataOut_payload_128_168 = (_zz_dataOut_payload_128_107 < _zz_dataOut_payload_128_43);
  assign _zz_dataOut_payload_128_169 = (_zz_dataOut_payload_128_168 ? _zz_dataOut_payload_128_107 : _zz_dataOut_payload_128_43);
  assign _zz_dataOut_payload_192_20 = (_zz_dataOut_payload_128_168 ? _zz_dataOut_payload_128_43 : _zz_dataOut_payload_128_107);
  assign _zz_dataOut_payload_128_170 = (_zz_dataOut_payload_128_106 < _zz_dataOut_payload_128_42);
  assign _zz_dataOut_payload_128_171 = (_zz_dataOut_payload_128_170 ? _zz_dataOut_payload_128_106 : _zz_dataOut_payload_128_42);
  assign _zz_dataOut_payload_192_21 = (_zz_dataOut_payload_128_170 ? _zz_dataOut_payload_128_42 : _zz_dataOut_payload_128_106);
  assign _zz_dataOut_payload_128_172 = (_zz_dataOut_payload_128_105 < _zz_dataOut_payload_128_41);
  assign _zz_dataOut_payload_128_173 = (_zz_dataOut_payload_128_172 ? _zz_dataOut_payload_128_105 : _zz_dataOut_payload_128_41);
  assign _zz_dataOut_payload_192_22 = (_zz_dataOut_payload_128_172 ? _zz_dataOut_payload_128_41 : _zz_dataOut_payload_128_105);
  assign _zz_dataOut_payload_128_174 = (_zz_dataOut_payload_128_104 < _zz_dataOut_payload_128_40);
  assign _zz_dataOut_payload_128_175 = (_zz_dataOut_payload_128_174 ? _zz_dataOut_payload_128_104 : _zz_dataOut_payload_128_40);
  assign _zz_dataOut_payload_192_23 = (_zz_dataOut_payload_128_174 ? _zz_dataOut_payload_128_40 : _zz_dataOut_payload_128_104);
  assign _zz_dataOut_payload_128_176 = (_zz_dataOut_payload_128_103 < _zz_dataOut_payload_128_39);
  assign _zz_dataOut_payload_128_177 = (_zz_dataOut_payload_128_176 ? _zz_dataOut_payload_128_103 : _zz_dataOut_payload_128_39);
  assign _zz_dataOut_payload_192_24 = (_zz_dataOut_payload_128_176 ? _zz_dataOut_payload_128_39 : _zz_dataOut_payload_128_103);
  assign _zz_dataOut_payload_128_178 = (_zz_dataOut_payload_128_102 < _zz_dataOut_payload_128_38);
  assign _zz_dataOut_payload_128_179 = (_zz_dataOut_payload_128_178 ? _zz_dataOut_payload_128_102 : _zz_dataOut_payload_128_38);
  assign _zz_dataOut_payload_192_25 = (_zz_dataOut_payload_128_178 ? _zz_dataOut_payload_128_38 : _zz_dataOut_payload_128_102);
  assign _zz_dataOut_payload_128_180 = (_zz_dataOut_payload_128_101 < _zz_dataOut_payload_128_37);
  assign _zz_dataOut_payload_128_181 = (_zz_dataOut_payload_128_180 ? _zz_dataOut_payload_128_101 : _zz_dataOut_payload_128_37);
  assign _zz_dataOut_payload_192_26 = (_zz_dataOut_payload_128_180 ? _zz_dataOut_payload_128_37 : _zz_dataOut_payload_128_101);
  assign _zz_dataOut_payload_128_182 = (_zz_dataOut_payload_128_100 < _zz_dataOut_payload_128_36);
  assign _zz_dataOut_payload_128_183 = (_zz_dataOut_payload_128_182 ? _zz_dataOut_payload_128_100 : _zz_dataOut_payload_128_36);
  assign _zz_dataOut_payload_192_27 = (_zz_dataOut_payload_128_182 ? _zz_dataOut_payload_128_36 : _zz_dataOut_payload_128_100);
  assign _zz_dataOut_payload_128_184 = (_zz_dataOut_payload_128_99 < _zz_dataOut_payload_128_35);
  assign _zz_dataOut_payload_128_185 = (_zz_dataOut_payload_128_184 ? _zz_dataOut_payload_128_99 : _zz_dataOut_payload_128_35);
  assign _zz_dataOut_payload_192_28 = (_zz_dataOut_payload_128_184 ? _zz_dataOut_payload_128_35 : _zz_dataOut_payload_128_99);
  assign _zz_dataOut_payload_128_186 = (_zz_dataOut_payload_128_98 < _zz_dataOut_payload_128_34);
  assign _zz_dataOut_payload_128_187 = (_zz_dataOut_payload_128_186 ? _zz_dataOut_payload_128_98 : _zz_dataOut_payload_128_34);
  assign _zz_dataOut_payload_192_29 = (_zz_dataOut_payload_128_186 ? _zz_dataOut_payload_128_34 : _zz_dataOut_payload_128_98);
  assign _zz_dataOut_payload_128_188 = (_zz_dataOut_payload_128_97 < _zz_dataOut_payload_128_33);
  assign _zz_dataOut_payload_128_189 = (_zz_dataOut_payload_128_188 ? _zz_dataOut_payload_128_97 : _zz_dataOut_payload_128_33);
  assign _zz_dataOut_payload_192_30 = (_zz_dataOut_payload_128_188 ? _zz_dataOut_payload_128_33 : _zz_dataOut_payload_128_97);
  assign _zz_dataOut_payload_128_190 = (_zz_dataOut_payload_128_96 < _zz_dataOut_payload_128_32);
  assign _zz_dataOut_payload_128_191 = (_zz_dataOut_payload_128_190 ? _zz_dataOut_payload_128_96 : _zz_dataOut_payload_128_32);
  assign _zz_dataOut_payload_192_31 = (_zz_dataOut_payload_128_190 ? _zz_dataOut_payload_128_32 : _zz_dataOut_payload_128_96);
  assign _zz_dataOut_payload_128_192 = (_zz_dataOut_payload_128_95 < _zz_dataOut_payload_128_31);
  assign _zz_dataOut_payload_128_193 = (_zz_dataOut_payload_128_192 ? _zz_dataOut_payload_128_95 : _zz_dataOut_payload_128_31);
  assign _zz_dataOut_payload_192_32 = (_zz_dataOut_payload_128_192 ? _zz_dataOut_payload_128_31 : _zz_dataOut_payload_128_95);
  assign _zz_dataOut_payload_128_194 = (_zz_dataOut_payload_128_94 < _zz_dataOut_payload_128_30);
  assign _zz_dataOut_payload_128_195 = (_zz_dataOut_payload_128_194 ? _zz_dataOut_payload_128_94 : _zz_dataOut_payload_128_30);
  assign _zz_dataOut_payload_192_33 = (_zz_dataOut_payload_128_194 ? _zz_dataOut_payload_128_30 : _zz_dataOut_payload_128_94);
  assign _zz_dataOut_payload_128_196 = (_zz_dataOut_payload_128_93 < _zz_dataOut_payload_128_29);
  assign _zz_dataOut_payload_128_197 = (_zz_dataOut_payload_128_196 ? _zz_dataOut_payload_128_93 : _zz_dataOut_payload_128_29);
  assign _zz_dataOut_payload_192_34 = (_zz_dataOut_payload_128_196 ? _zz_dataOut_payload_128_29 : _zz_dataOut_payload_128_93);
  assign _zz_dataOut_payload_128_198 = (_zz_dataOut_payload_128_92 < _zz_dataOut_payload_128_28);
  assign _zz_dataOut_payload_128_199 = (_zz_dataOut_payload_128_198 ? _zz_dataOut_payload_128_92 : _zz_dataOut_payload_128_28);
  assign _zz_dataOut_payload_192_35 = (_zz_dataOut_payload_128_198 ? _zz_dataOut_payload_128_28 : _zz_dataOut_payload_128_92);
  assign _zz_dataOut_payload_128_200 = (_zz_dataOut_payload_128_91 < _zz_dataOut_payload_128_27);
  assign _zz_dataOut_payload_128_201 = (_zz_dataOut_payload_128_200 ? _zz_dataOut_payload_128_91 : _zz_dataOut_payload_128_27);
  assign _zz_dataOut_payload_192_36 = (_zz_dataOut_payload_128_200 ? _zz_dataOut_payload_128_27 : _zz_dataOut_payload_128_91);
  assign _zz_dataOut_payload_128_202 = (_zz_dataOut_payload_128_90 < _zz_dataOut_payload_128_26);
  assign _zz_dataOut_payload_128_203 = (_zz_dataOut_payload_128_202 ? _zz_dataOut_payload_128_90 : _zz_dataOut_payload_128_26);
  assign _zz_dataOut_payload_192_37 = (_zz_dataOut_payload_128_202 ? _zz_dataOut_payload_128_26 : _zz_dataOut_payload_128_90);
  assign _zz_dataOut_payload_128_204 = (_zz_dataOut_payload_128_89 < _zz_dataOut_payload_128_25);
  assign _zz_dataOut_payload_128_205 = (_zz_dataOut_payload_128_204 ? _zz_dataOut_payload_128_89 : _zz_dataOut_payload_128_25);
  assign _zz_dataOut_payload_192_38 = (_zz_dataOut_payload_128_204 ? _zz_dataOut_payload_128_25 : _zz_dataOut_payload_128_89);
  assign _zz_dataOut_payload_128_206 = (_zz_dataOut_payload_128_88 < _zz_dataOut_payload_128_24);
  assign _zz_dataOut_payload_128_207 = (_zz_dataOut_payload_128_206 ? _zz_dataOut_payload_128_88 : _zz_dataOut_payload_128_24);
  assign _zz_dataOut_payload_192_39 = (_zz_dataOut_payload_128_206 ? _zz_dataOut_payload_128_24 : _zz_dataOut_payload_128_88);
  assign _zz_dataOut_payload_128_208 = (_zz_dataOut_payload_128_87 < _zz_dataOut_payload_128_23);
  assign _zz_dataOut_payload_128_209 = (_zz_dataOut_payload_128_208 ? _zz_dataOut_payload_128_87 : _zz_dataOut_payload_128_23);
  assign _zz_dataOut_payload_192_40 = (_zz_dataOut_payload_128_208 ? _zz_dataOut_payload_128_23 : _zz_dataOut_payload_128_87);
  assign _zz_dataOut_payload_128_210 = (_zz_dataOut_payload_128_86 < _zz_dataOut_payload_128_22);
  assign _zz_dataOut_payload_128_211 = (_zz_dataOut_payload_128_210 ? _zz_dataOut_payload_128_86 : _zz_dataOut_payload_128_22);
  assign _zz_dataOut_payload_192_41 = (_zz_dataOut_payload_128_210 ? _zz_dataOut_payload_128_22 : _zz_dataOut_payload_128_86);
  assign _zz_dataOut_payload_128_212 = (_zz_dataOut_payload_128_85 < _zz_dataOut_payload_128_21);
  assign _zz_dataOut_payload_128_213 = (_zz_dataOut_payload_128_212 ? _zz_dataOut_payload_128_85 : _zz_dataOut_payload_128_21);
  assign _zz_dataOut_payload_192_42 = (_zz_dataOut_payload_128_212 ? _zz_dataOut_payload_128_21 : _zz_dataOut_payload_128_85);
  assign _zz_dataOut_payload_128_214 = (_zz_dataOut_payload_128_84 < _zz_dataOut_payload_128_20);
  assign _zz_dataOut_payload_128_215 = (_zz_dataOut_payload_128_214 ? _zz_dataOut_payload_128_84 : _zz_dataOut_payload_128_20);
  assign _zz_dataOut_payload_192_43 = (_zz_dataOut_payload_128_214 ? _zz_dataOut_payload_128_20 : _zz_dataOut_payload_128_84);
  assign _zz_dataOut_payload_128_216 = (_zz_dataOut_payload_128_83 < _zz_dataOut_payload_128_19);
  assign _zz_dataOut_payload_128_217 = (_zz_dataOut_payload_128_216 ? _zz_dataOut_payload_128_83 : _zz_dataOut_payload_128_19);
  assign _zz_dataOut_payload_192_44 = (_zz_dataOut_payload_128_216 ? _zz_dataOut_payload_128_19 : _zz_dataOut_payload_128_83);
  assign _zz_dataOut_payload_128_218 = (_zz_dataOut_payload_128_82 < _zz_dataOut_payload_128_18);
  assign _zz_dataOut_payload_128_219 = (_zz_dataOut_payload_128_218 ? _zz_dataOut_payload_128_82 : _zz_dataOut_payload_128_18);
  assign _zz_dataOut_payload_192_45 = (_zz_dataOut_payload_128_218 ? _zz_dataOut_payload_128_18 : _zz_dataOut_payload_128_82);
  assign _zz_dataOut_payload_128_220 = (_zz_dataOut_payload_128_81 < _zz_dataOut_payload_128_17);
  assign _zz_dataOut_payload_128_221 = (_zz_dataOut_payload_128_220 ? _zz_dataOut_payload_128_81 : _zz_dataOut_payload_128_17);
  assign _zz_dataOut_payload_192_46 = (_zz_dataOut_payload_128_220 ? _zz_dataOut_payload_128_17 : _zz_dataOut_payload_128_81);
  assign _zz_dataOut_payload_128_222 = (_zz_dataOut_payload_128_80 < _zz_dataOut_payload_128_16);
  assign _zz_dataOut_payload_128_223 = (_zz_dataOut_payload_128_222 ? _zz_dataOut_payload_128_80 : _zz_dataOut_payload_128_16);
  assign _zz_dataOut_payload_192_47 = (_zz_dataOut_payload_128_222 ? _zz_dataOut_payload_128_16 : _zz_dataOut_payload_128_80);
  assign _zz_dataOut_payload_128_224 = (_zz_dataOut_payload_128_79 < _zz_dataOut_payload_128_15);
  assign _zz_dataOut_payload_128_225 = (_zz_dataOut_payload_128_224 ? _zz_dataOut_payload_128_79 : _zz_dataOut_payload_128_15);
  assign _zz_dataOut_payload_192_48 = (_zz_dataOut_payload_128_224 ? _zz_dataOut_payload_128_15 : _zz_dataOut_payload_128_79);
  assign _zz_dataOut_payload_128_226 = (_zz_dataOut_payload_128_78 < _zz_dataOut_payload_128_14);
  assign _zz_dataOut_payload_128_227 = (_zz_dataOut_payload_128_226 ? _zz_dataOut_payload_128_78 : _zz_dataOut_payload_128_14);
  assign _zz_dataOut_payload_192_49 = (_zz_dataOut_payload_128_226 ? _zz_dataOut_payload_128_14 : _zz_dataOut_payload_128_78);
  assign _zz_dataOut_payload_128_228 = (_zz_dataOut_payload_128_77 < _zz_dataOut_payload_128_13);
  assign _zz_dataOut_payload_128_229 = (_zz_dataOut_payload_128_228 ? _zz_dataOut_payload_128_77 : _zz_dataOut_payload_128_13);
  assign _zz_dataOut_payload_192_50 = (_zz_dataOut_payload_128_228 ? _zz_dataOut_payload_128_13 : _zz_dataOut_payload_128_77);
  assign _zz_dataOut_payload_128_230 = (_zz_dataOut_payload_128_76 < _zz_dataOut_payload_128_12);
  assign _zz_dataOut_payload_128_231 = (_zz_dataOut_payload_128_230 ? _zz_dataOut_payload_128_76 : _zz_dataOut_payload_128_12);
  assign _zz_dataOut_payload_192_51 = (_zz_dataOut_payload_128_230 ? _zz_dataOut_payload_128_12 : _zz_dataOut_payload_128_76);
  assign _zz_dataOut_payload_128_232 = (_zz_dataOut_payload_128_75 < _zz_dataOut_payload_128_11);
  assign _zz_dataOut_payload_128_233 = (_zz_dataOut_payload_128_232 ? _zz_dataOut_payload_128_75 : _zz_dataOut_payload_128_11);
  assign _zz_dataOut_payload_192_52 = (_zz_dataOut_payload_128_232 ? _zz_dataOut_payload_128_11 : _zz_dataOut_payload_128_75);
  assign _zz_dataOut_payload_128_234 = (_zz_dataOut_payload_128_74 < _zz_dataOut_payload_128_10);
  assign _zz_dataOut_payload_128_235 = (_zz_dataOut_payload_128_234 ? _zz_dataOut_payload_128_74 : _zz_dataOut_payload_128_10);
  assign _zz_dataOut_payload_192_53 = (_zz_dataOut_payload_128_234 ? _zz_dataOut_payload_128_10 : _zz_dataOut_payload_128_74);
  assign _zz_dataOut_payload_128_236 = (_zz_dataOut_payload_128_73 < _zz_dataOut_payload_128_9);
  assign _zz_dataOut_payload_128_237 = (_zz_dataOut_payload_128_236 ? _zz_dataOut_payload_128_73 : _zz_dataOut_payload_128_9);
  assign _zz_dataOut_payload_192_54 = (_zz_dataOut_payload_128_236 ? _zz_dataOut_payload_128_9 : _zz_dataOut_payload_128_73);
  assign _zz_dataOut_payload_128_238 = (_zz_dataOut_payload_128_72 < _zz_dataOut_payload_128_8);
  assign _zz_dataOut_payload_128_239 = (_zz_dataOut_payload_128_238 ? _zz_dataOut_payload_128_72 : _zz_dataOut_payload_128_8);
  assign _zz_dataOut_payload_192_55 = (_zz_dataOut_payload_128_238 ? _zz_dataOut_payload_128_8 : _zz_dataOut_payload_128_72);
  assign _zz_dataOut_payload_128_240 = (_zz_dataOut_payload_128_71 < _zz_dataOut_payload_128_7);
  assign _zz_dataOut_payload_128_241 = (_zz_dataOut_payload_128_240 ? _zz_dataOut_payload_128_71 : _zz_dataOut_payload_128_7);
  assign _zz_dataOut_payload_192_56 = (_zz_dataOut_payload_128_240 ? _zz_dataOut_payload_128_7 : _zz_dataOut_payload_128_71);
  assign _zz_dataOut_payload_128_242 = (_zz_dataOut_payload_128_70 < _zz_dataOut_payload_128_6);
  assign _zz_dataOut_payload_128_243 = (_zz_dataOut_payload_128_242 ? _zz_dataOut_payload_128_70 : _zz_dataOut_payload_128_6);
  assign _zz_dataOut_payload_192_57 = (_zz_dataOut_payload_128_242 ? _zz_dataOut_payload_128_6 : _zz_dataOut_payload_128_70);
  assign _zz_dataOut_payload_128_244 = (_zz_dataOut_payload_128_69 < _zz_dataOut_payload_128_5);
  assign _zz_dataOut_payload_128_245 = (_zz_dataOut_payload_128_244 ? _zz_dataOut_payload_128_69 : _zz_dataOut_payload_128_5);
  assign _zz_dataOut_payload_192_58 = (_zz_dataOut_payload_128_244 ? _zz_dataOut_payload_128_5 : _zz_dataOut_payload_128_69);
  assign _zz_dataOut_payload_128_246 = (_zz_dataOut_payload_128_68 < _zz_dataOut_payload_128_4);
  assign _zz_dataOut_payload_128_247 = (_zz_dataOut_payload_128_246 ? _zz_dataOut_payload_128_68 : _zz_dataOut_payload_128_4);
  assign _zz_dataOut_payload_192_59 = (_zz_dataOut_payload_128_246 ? _zz_dataOut_payload_128_4 : _zz_dataOut_payload_128_68);
  assign _zz_dataOut_payload_128_248 = (_zz_dataOut_payload_128_67 < _zz_dataOut_payload_128_3);
  assign _zz_dataOut_payload_128_249 = (_zz_dataOut_payload_128_248 ? _zz_dataOut_payload_128_67 : _zz_dataOut_payload_128_3);
  assign _zz_dataOut_payload_192_60 = (_zz_dataOut_payload_128_248 ? _zz_dataOut_payload_128_3 : _zz_dataOut_payload_128_67);
  assign _zz_dataOut_payload_128_250 = (_zz_dataOut_payload_128_66 < _zz_dataOut_payload_128_2);
  assign _zz_dataOut_payload_128_251 = (_zz_dataOut_payload_128_250 ? _zz_dataOut_payload_128_66 : _zz_dataOut_payload_128_2);
  assign _zz_dataOut_payload_192_61 = (_zz_dataOut_payload_128_250 ? _zz_dataOut_payload_128_2 : _zz_dataOut_payload_128_66);
  assign _zz_dataOut_payload_128_252 = (_zz_dataOut_payload_128_65 < _zz_dataOut_payload_128_1);
  assign _zz_dataOut_payload_128_253 = (_zz_dataOut_payload_128_252 ? _zz_dataOut_payload_128_65 : _zz_dataOut_payload_128_1);
  assign _zz_dataOut_payload_192_62 = (_zz_dataOut_payload_128_252 ? _zz_dataOut_payload_128_1 : _zz_dataOut_payload_128_65);
  assign _zz_dataOut_payload_128_254 = (_zz_dataOut_payload_128_64 < _zz_dataOut_payload_128);
  assign _zz_dataOut_payload_128_255 = (_zz_dataOut_payload_128_254 ? _zz_dataOut_payload_128_64 : _zz_dataOut_payload_128);
  assign _zz_dataOut_payload_192_63 = (_zz_dataOut_payload_128_254 ? _zz_dataOut_payload_128 : _zz_dataOut_payload_128_64);
  assign _zz_dataOut_payload_128_256 = (_zz_dataOut_payload_128_129 < _zz_dataOut_payload_128_193);
  assign _zz_dataOut_payload_128_257 = (_zz_dataOut_payload_128_256 ? _zz_dataOut_payload_128_129 : _zz_dataOut_payload_128_193);
  assign _zz_dataOut_payload_160 = (_zz_dataOut_payload_128_256 ? _zz_dataOut_payload_128_193 : _zz_dataOut_payload_128_129);
  assign _zz_dataOut_payload_128_258 = (_zz_dataOut_payload_128_131 < _zz_dataOut_payload_128_195);
  assign _zz_dataOut_payload_128_259 = (_zz_dataOut_payload_128_258 ? _zz_dataOut_payload_128_131 : _zz_dataOut_payload_128_195);
  assign _zz_dataOut_payload_160_1 = (_zz_dataOut_payload_128_258 ? _zz_dataOut_payload_128_195 : _zz_dataOut_payload_128_131);
  assign _zz_dataOut_payload_128_260 = (_zz_dataOut_payload_128_133 < _zz_dataOut_payload_128_197);
  assign _zz_dataOut_payload_128_261 = (_zz_dataOut_payload_128_260 ? _zz_dataOut_payload_128_133 : _zz_dataOut_payload_128_197);
  assign _zz_dataOut_payload_160_2 = (_zz_dataOut_payload_128_260 ? _zz_dataOut_payload_128_197 : _zz_dataOut_payload_128_133);
  assign _zz_dataOut_payload_128_262 = (_zz_dataOut_payload_128_135 < _zz_dataOut_payload_128_199);
  assign _zz_dataOut_payload_128_263 = (_zz_dataOut_payload_128_262 ? _zz_dataOut_payload_128_135 : _zz_dataOut_payload_128_199);
  assign _zz_dataOut_payload_160_3 = (_zz_dataOut_payload_128_262 ? _zz_dataOut_payload_128_199 : _zz_dataOut_payload_128_135);
  assign _zz_dataOut_payload_128_264 = (_zz_dataOut_payload_128_137 < _zz_dataOut_payload_128_201);
  assign _zz_dataOut_payload_128_265 = (_zz_dataOut_payload_128_264 ? _zz_dataOut_payload_128_137 : _zz_dataOut_payload_128_201);
  assign _zz_dataOut_payload_160_4 = (_zz_dataOut_payload_128_264 ? _zz_dataOut_payload_128_201 : _zz_dataOut_payload_128_137);
  assign _zz_dataOut_payload_128_266 = (_zz_dataOut_payload_128_139 < _zz_dataOut_payload_128_203);
  assign _zz_dataOut_payload_128_267 = (_zz_dataOut_payload_128_266 ? _zz_dataOut_payload_128_139 : _zz_dataOut_payload_128_203);
  assign _zz_dataOut_payload_160_5 = (_zz_dataOut_payload_128_266 ? _zz_dataOut_payload_128_203 : _zz_dataOut_payload_128_139);
  assign _zz_dataOut_payload_128_268 = (_zz_dataOut_payload_128_141 < _zz_dataOut_payload_128_205);
  assign _zz_dataOut_payload_128_269 = (_zz_dataOut_payload_128_268 ? _zz_dataOut_payload_128_141 : _zz_dataOut_payload_128_205);
  assign _zz_dataOut_payload_160_6 = (_zz_dataOut_payload_128_268 ? _zz_dataOut_payload_128_205 : _zz_dataOut_payload_128_141);
  assign _zz_dataOut_payload_128_270 = (_zz_dataOut_payload_128_143 < _zz_dataOut_payload_128_207);
  assign _zz_dataOut_payload_128_271 = (_zz_dataOut_payload_128_270 ? _zz_dataOut_payload_128_143 : _zz_dataOut_payload_128_207);
  assign _zz_dataOut_payload_160_7 = (_zz_dataOut_payload_128_270 ? _zz_dataOut_payload_128_207 : _zz_dataOut_payload_128_143);
  assign _zz_dataOut_payload_128_272 = (_zz_dataOut_payload_128_145 < _zz_dataOut_payload_128_209);
  assign _zz_dataOut_payload_128_273 = (_zz_dataOut_payload_128_272 ? _zz_dataOut_payload_128_145 : _zz_dataOut_payload_128_209);
  assign _zz_dataOut_payload_160_8 = (_zz_dataOut_payload_128_272 ? _zz_dataOut_payload_128_209 : _zz_dataOut_payload_128_145);
  assign _zz_dataOut_payload_128_274 = (_zz_dataOut_payload_128_147 < _zz_dataOut_payload_128_211);
  assign _zz_dataOut_payload_128_275 = (_zz_dataOut_payload_128_274 ? _zz_dataOut_payload_128_147 : _zz_dataOut_payload_128_211);
  assign _zz_dataOut_payload_160_9 = (_zz_dataOut_payload_128_274 ? _zz_dataOut_payload_128_211 : _zz_dataOut_payload_128_147);
  assign _zz_dataOut_payload_128_276 = (_zz_dataOut_payload_128_149 < _zz_dataOut_payload_128_213);
  assign _zz_dataOut_payload_128_277 = (_zz_dataOut_payload_128_276 ? _zz_dataOut_payload_128_149 : _zz_dataOut_payload_128_213);
  assign _zz_dataOut_payload_160_10 = (_zz_dataOut_payload_128_276 ? _zz_dataOut_payload_128_213 : _zz_dataOut_payload_128_149);
  assign _zz_dataOut_payload_128_278 = (_zz_dataOut_payload_128_151 < _zz_dataOut_payload_128_215);
  assign _zz_dataOut_payload_128_279 = (_zz_dataOut_payload_128_278 ? _zz_dataOut_payload_128_151 : _zz_dataOut_payload_128_215);
  assign _zz_dataOut_payload_160_11 = (_zz_dataOut_payload_128_278 ? _zz_dataOut_payload_128_215 : _zz_dataOut_payload_128_151);
  assign _zz_dataOut_payload_128_280 = (_zz_dataOut_payload_128_153 < _zz_dataOut_payload_128_217);
  assign _zz_dataOut_payload_128_281 = (_zz_dataOut_payload_128_280 ? _zz_dataOut_payload_128_153 : _zz_dataOut_payload_128_217);
  assign _zz_dataOut_payload_160_12 = (_zz_dataOut_payload_128_280 ? _zz_dataOut_payload_128_217 : _zz_dataOut_payload_128_153);
  assign _zz_dataOut_payload_128_282 = (_zz_dataOut_payload_128_155 < _zz_dataOut_payload_128_219);
  assign _zz_dataOut_payload_128_283 = (_zz_dataOut_payload_128_282 ? _zz_dataOut_payload_128_155 : _zz_dataOut_payload_128_219);
  assign _zz_dataOut_payload_160_13 = (_zz_dataOut_payload_128_282 ? _zz_dataOut_payload_128_219 : _zz_dataOut_payload_128_155);
  assign _zz_dataOut_payload_128_284 = (_zz_dataOut_payload_128_157 < _zz_dataOut_payload_128_221);
  assign _zz_dataOut_payload_128_285 = (_zz_dataOut_payload_128_284 ? _zz_dataOut_payload_128_157 : _zz_dataOut_payload_128_221);
  assign _zz_dataOut_payload_160_14 = (_zz_dataOut_payload_128_284 ? _zz_dataOut_payload_128_221 : _zz_dataOut_payload_128_157);
  assign _zz_dataOut_payload_128_286 = (_zz_dataOut_payload_128_159 < _zz_dataOut_payload_128_223);
  assign _zz_dataOut_payload_128_287 = (_zz_dataOut_payload_128_286 ? _zz_dataOut_payload_128_159 : _zz_dataOut_payload_128_223);
  assign _zz_dataOut_payload_160_15 = (_zz_dataOut_payload_128_286 ? _zz_dataOut_payload_128_223 : _zz_dataOut_payload_128_159);
  assign _zz_dataOut_payload_128_288 = (_zz_dataOut_payload_128_161 < _zz_dataOut_payload_128_225);
  assign _zz_dataOut_payload_128_289 = (_zz_dataOut_payload_128_288 ? _zz_dataOut_payload_128_161 : _zz_dataOut_payload_128_225);
  assign _zz_dataOut_payload_160_16 = (_zz_dataOut_payload_128_288 ? _zz_dataOut_payload_128_225 : _zz_dataOut_payload_128_161);
  assign _zz_dataOut_payload_128_290 = (_zz_dataOut_payload_128_163 < _zz_dataOut_payload_128_227);
  assign _zz_dataOut_payload_128_291 = (_zz_dataOut_payload_128_290 ? _zz_dataOut_payload_128_163 : _zz_dataOut_payload_128_227);
  assign _zz_dataOut_payload_160_17 = (_zz_dataOut_payload_128_290 ? _zz_dataOut_payload_128_227 : _zz_dataOut_payload_128_163);
  assign _zz_dataOut_payload_128_292 = (_zz_dataOut_payload_128_165 < _zz_dataOut_payload_128_229);
  assign _zz_dataOut_payload_128_293 = (_zz_dataOut_payload_128_292 ? _zz_dataOut_payload_128_165 : _zz_dataOut_payload_128_229);
  assign _zz_dataOut_payload_160_18 = (_zz_dataOut_payload_128_292 ? _zz_dataOut_payload_128_229 : _zz_dataOut_payload_128_165);
  assign _zz_dataOut_payload_128_294 = (_zz_dataOut_payload_128_167 < _zz_dataOut_payload_128_231);
  assign _zz_dataOut_payload_128_295 = (_zz_dataOut_payload_128_294 ? _zz_dataOut_payload_128_167 : _zz_dataOut_payload_128_231);
  assign _zz_dataOut_payload_160_19 = (_zz_dataOut_payload_128_294 ? _zz_dataOut_payload_128_231 : _zz_dataOut_payload_128_167);
  assign _zz_dataOut_payload_128_296 = (_zz_dataOut_payload_128_169 < _zz_dataOut_payload_128_233);
  assign _zz_dataOut_payload_128_297 = (_zz_dataOut_payload_128_296 ? _zz_dataOut_payload_128_169 : _zz_dataOut_payload_128_233);
  assign _zz_dataOut_payload_160_20 = (_zz_dataOut_payload_128_296 ? _zz_dataOut_payload_128_233 : _zz_dataOut_payload_128_169);
  assign _zz_dataOut_payload_128_298 = (_zz_dataOut_payload_128_171 < _zz_dataOut_payload_128_235);
  assign _zz_dataOut_payload_128_299 = (_zz_dataOut_payload_128_298 ? _zz_dataOut_payload_128_171 : _zz_dataOut_payload_128_235);
  assign _zz_dataOut_payload_160_21 = (_zz_dataOut_payload_128_298 ? _zz_dataOut_payload_128_235 : _zz_dataOut_payload_128_171);
  assign _zz_dataOut_payload_128_300 = (_zz_dataOut_payload_128_173 < _zz_dataOut_payload_128_237);
  assign _zz_dataOut_payload_128_301 = (_zz_dataOut_payload_128_300 ? _zz_dataOut_payload_128_173 : _zz_dataOut_payload_128_237);
  assign _zz_dataOut_payload_160_22 = (_zz_dataOut_payload_128_300 ? _zz_dataOut_payload_128_237 : _zz_dataOut_payload_128_173);
  assign _zz_dataOut_payload_128_302 = (_zz_dataOut_payload_128_175 < _zz_dataOut_payload_128_239);
  assign _zz_dataOut_payload_128_303 = (_zz_dataOut_payload_128_302 ? _zz_dataOut_payload_128_175 : _zz_dataOut_payload_128_239);
  assign _zz_dataOut_payload_160_23 = (_zz_dataOut_payload_128_302 ? _zz_dataOut_payload_128_239 : _zz_dataOut_payload_128_175);
  assign _zz_dataOut_payload_128_304 = (_zz_dataOut_payload_128_177 < _zz_dataOut_payload_128_241);
  assign _zz_dataOut_payload_128_305 = (_zz_dataOut_payload_128_304 ? _zz_dataOut_payload_128_177 : _zz_dataOut_payload_128_241);
  assign _zz_dataOut_payload_160_24 = (_zz_dataOut_payload_128_304 ? _zz_dataOut_payload_128_241 : _zz_dataOut_payload_128_177);
  assign _zz_dataOut_payload_128_306 = (_zz_dataOut_payload_128_179 < _zz_dataOut_payload_128_243);
  assign _zz_dataOut_payload_128_307 = (_zz_dataOut_payload_128_306 ? _zz_dataOut_payload_128_179 : _zz_dataOut_payload_128_243);
  assign _zz_dataOut_payload_160_25 = (_zz_dataOut_payload_128_306 ? _zz_dataOut_payload_128_243 : _zz_dataOut_payload_128_179);
  assign _zz_dataOut_payload_128_308 = (_zz_dataOut_payload_128_181 < _zz_dataOut_payload_128_245);
  assign _zz_dataOut_payload_128_309 = (_zz_dataOut_payload_128_308 ? _zz_dataOut_payload_128_181 : _zz_dataOut_payload_128_245);
  assign _zz_dataOut_payload_160_26 = (_zz_dataOut_payload_128_308 ? _zz_dataOut_payload_128_245 : _zz_dataOut_payload_128_181);
  assign _zz_dataOut_payload_128_310 = (_zz_dataOut_payload_128_183 < _zz_dataOut_payload_128_247);
  assign _zz_dataOut_payload_128_311 = (_zz_dataOut_payload_128_310 ? _zz_dataOut_payload_128_183 : _zz_dataOut_payload_128_247);
  assign _zz_dataOut_payload_160_27 = (_zz_dataOut_payload_128_310 ? _zz_dataOut_payload_128_247 : _zz_dataOut_payload_128_183);
  assign _zz_dataOut_payload_128_312 = (_zz_dataOut_payload_128_185 < _zz_dataOut_payload_128_249);
  assign _zz_dataOut_payload_128_313 = (_zz_dataOut_payload_128_312 ? _zz_dataOut_payload_128_185 : _zz_dataOut_payload_128_249);
  assign _zz_dataOut_payload_160_28 = (_zz_dataOut_payload_128_312 ? _zz_dataOut_payload_128_249 : _zz_dataOut_payload_128_185);
  assign _zz_dataOut_payload_128_314 = (_zz_dataOut_payload_128_187 < _zz_dataOut_payload_128_251);
  assign _zz_dataOut_payload_128_315 = (_zz_dataOut_payload_128_314 ? _zz_dataOut_payload_128_187 : _zz_dataOut_payload_128_251);
  assign _zz_dataOut_payload_160_29 = (_zz_dataOut_payload_128_314 ? _zz_dataOut_payload_128_251 : _zz_dataOut_payload_128_187);
  assign _zz_dataOut_payload_128_316 = (_zz_dataOut_payload_128_189 < _zz_dataOut_payload_128_253);
  assign _zz_dataOut_payload_128_317 = (_zz_dataOut_payload_128_316 ? _zz_dataOut_payload_128_189 : _zz_dataOut_payload_128_253);
  assign _zz_dataOut_payload_160_30 = (_zz_dataOut_payload_128_316 ? _zz_dataOut_payload_128_253 : _zz_dataOut_payload_128_189);
  assign _zz_dataOut_payload_128_318 = (_zz_dataOut_payload_128_191 < _zz_dataOut_payload_128_255);
  assign _zz_dataOut_payload_128_319 = (_zz_dataOut_payload_128_318 ? _zz_dataOut_payload_128_191 : _zz_dataOut_payload_128_255);
  assign _zz_dataOut_payload_160_31 = (_zz_dataOut_payload_128_318 ? _zz_dataOut_payload_128_255 : _zz_dataOut_payload_128_191);
  assign _zz_dataOut_payload_128_320 = (_zz_dataOut_payload_128_257 < _zz_dataOut_payload_128_289);
  assign _zz_dataOut_payload_128_321 = (_zz_dataOut_payload_128_320 ? _zz_dataOut_payload_128_257 : _zz_dataOut_payload_128_289);
  assign _zz_dataOut_payload_144 = (_zz_dataOut_payload_128_320 ? _zz_dataOut_payload_128_289 : _zz_dataOut_payload_128_257);
  assign _zz_dataOut_payload_128_322 = (_zz_dataOut_payload_128_259 < _zz_dataOut_payload_128_291);
  assign _zz_dataOut_payload_128_323 = (_zz_dataOut_payload_128_322 ? _zz_dataOut_payload_128_259 : _zz_dataOut_payload_128_291);
  assign _zz_dataOut_payload_144_1 = (_zz_dataOut_payload_128_322 ? _zz_dataOut_payload_128_291 : _zz_dataOut_payload_128_259);
  assign _zz_dataOut_payload_128_324 = (_zz_dataOut_payload_128_261 < _zz_dataOut_payload_128_293);
  assign _zz_dataOut_payload_128_325 = (_zz_dataOut_payload_128_324 ? _zz_dataOut_payload_128_261 : _zz_dataOut_payload_128_293);
  assign _zz_dataOut_payload_144_2 = (_zz_dataOut_payload_128_324 ? _zz_dataOut_payload_128_293 : _zz_dataOut_payload_128_261);
  assign _zz_dataOut_payload_128_326 = (_zz_dataOut_payload_128_263 < _zz_dataOut_payload_128_295);
  assign _zz_dataOut_payload_128_327 = (_zz_dataOut_payload_128_326 ? _zz_dataOut_payload_128_263 : _zz_dataOut_payload_128_295);
  assign _zz_dataOut_payload_144_3 = (_zz_dataOut_payload_128_326 ? _zz_dataOut_payload_128_295 : _zz_dataOut_payload_128_263);
  assign _zz_dataOut_payload_128_328 = (_zz_dataOut_payload_128_265 < _zz_dataOut_payload_128_297);
  assign _zz_dataOut_payload_128_329 = (_zz_dataOut_payload_128_328 ? _zz_dataOut_payload_128_265 : _zz_dataOut_payload_128_297);
  assign _zz_dataOut_payload_144_4 = (_zz_dataOut_payload_128_328 ? _zz_dataOut_payload_128_297 : _zz_dataOut_payload_128_265);
  assign _zz_dataOut_payload_128_330 = (_zz_dataOut_payload_128_267 < _zz_dataOut_payload_128_299);
  assign _zz_dataOut_payload_128_331 = (_zz_dataOut_payload_128_330 ? _zz_dataOut_payload_128_267 : _zz_dataOut_payload_128_299);
  assign _zz_dataOut_payload_144_5 = (_zz_dataOut_payload_128_330 ? _zz_dataOut_payload_128_299 : _zz_dataOut_payload_128_267);
  assign _zz_dataOut_payload_128_332 = (_zz_dataOut_payload_128_269 < _zz_dataOut_payload_128_301);
  assign _zz_dataOut_payload_128_333 = (_zz_dataOut_payload_128_332 ? _zz_dataOut_payload_128_269 : _zz_dataOut_payload_128_301);
  assign _zz_dataOut_payload_144_6 = (_zz_dataOut_payload_128_332 ? _zz_dataOut_payload_128_301 : _zz_dataOut_payload_128_269);
  assign _zz_dataOut_payload_128_334 = (_zz_dataOut_payload_128_271 < _zz_dataOut_payload_128_303);
  assign _zz_dataOut_payload_128_335 = (_zz_dataOut_payload_128_334 ? _zz_dataOut_payload_128_271 : _zz_dataOut_payload_128_303);
  assign _zz_dataOut_payload_144_7 = (_zz_dataOut_payload_128_334 ? _zz_dataOut_payload_128_303 : _zz_dataOut_payload_128_271);
  assign _zz_dataOut_payload_128_336 = (_zz_dataOut_payload_128_273 < _zz_dataOut_payload_128_305);
  assign _zz_dataOut_payload_128_337 = (_zz_dataOut_payload_128_336 ? _zz_dataOut_payload_128_273 : _zz_dataOut_payload_128_305);
  assign _zz_dataOut_payload_144_8 = (_zz_dataOut_payload_128_336 ? _zz_dataOut_payload_128_305 : _zz_dataOut_payload_128_273);
  assign _zz_dataOut_payload_128_338 = (_zz_dataOut_payload_128_275 < _zz_dataOut_payload_128_307);
  assign _zz_dataOut_payload_128_339 = (_zz_dataOut_payload_128_338 ? _zz_dataOut_payload_128_275 : _zz_dataOut_payload_128_307);
  assign _zz_dataOut_payload_144_9 = (_zz_dataOut_payload_128_338 ? _zz_dataOut_payload_128_307 : _zz_dataOut_payload_128_275);
  assign _zz_dataOut_payload_128_340 = (_zz_dataOut_payload_128_277 < _zz_dataOut_payload_128_309);
  assign _zz_dataOut_payload_128_341 = (_zz_dataOut_payload_128_340 ? _zz_dataOut_payload_128_277 : _zz_dataOut_payload_128_309);
  assign _zz_dataOut_payload_144_10 = (_zz_dataOut_payload_128_340 ? _zz_dataOut_payload_128_309 : _zz_dataOut_payload_128_277);
  assign _zz_dataOut_payload_128_342 = (_zz_dataOut_payload_128_279 < _zz_dataOut_payload_128_311);
  assign _zz_dataOut_payload_128_343 = (_zz_dataOut_payload_128_342 ? _zz_dataOut_payload_128_279 : _zz_dataOut_payload_128_311);
  assign _zz_dataOut_payload_144_11 = (_zz_dataOut_payload_128_342 ? _zz_dataOut_payload_128_311 : _zz_dataOut_payload_128_279);
  assign _zz_dataOut_payload_128_344 = (_zz_dataOut_payload_128_281 < _zz_dataOut_payload_128_313);
  assign _zz_dataOut_payload_128_345 = (_zz_dataOut_payload_128_344 ? _zz_dataOut_payload_128_281 : _zz_dataOut_payload_128_313);
  assign _zz_dataOut_payload_144_12 = (_zz_dataOut_payload_128_344 ? _zz_dataOut_payload_128_313 : _zz_dataOut_payload_128_281);
  assign _zz_dataOut_payload_128_346 = (_zz_dataOut_payload_128_283 < _zz_dataOut_payload_128_315);
  assign _zz_dataOut_payload_128_347 = (_zz_dataOut_payload_128_346 ? _zz_dataOut_payload_128_283 : _zz_dataOut_payload_128_315);
  assign _zz_dataOut_payload_144_13 = (_zz_dataOut_payload_128_346 ? _zz_dataOut_payload_128_315 : _zz_dataOut_payload_128_283);
  assign _zz_dataOut_payload_128_348 = (_zz_dataOut_payload_128_285 < _zz_dataOut_payload_128_317);
  assign _zz_dataOut_payload_128_349 = (_zz_dataOut_payload_128_348 ? _zz_dataOut_payload_128_285 : _zz_dataOut_payload_128_317);
  assign _zz_dataOut_payload_144_14 = (_zz_dataOut_payload_128_348 ? _zz_dataOut_payload_128_317 : _zz_dataOut_payload_128_285);
  assign _zz_dataOut_payload_128_350 = (_zz_dataOut_payload_128_287 < _zz_dataOut_payload_128_319);
  assign _zz_dataOut_payload_128_351 = (_zz_dataOut_payload_128_350 ? _zz_dataOut_payload_128_287 : _zz_dataOut_payload_128_319);
  assign _zz_dataOut_payload_144_15 = (_zz_dataOut_payload_128_350 ? _zz_dataOut_payload_128_319 : _zz_dataOut_payload_128_287);
  assign _zz_dataOut_payload_128_352 = (_zz_dataOut_payload_128_321 < _zz_dataOut_payload_128_337);
  assign _zz_dataOut_payload_128_353 = (_zz_dataOut_payload_128_352 ? _zz_dataOut_payload_128_321 : _zz_dataOut_payload_128_337);
  assign _zz_dataOut_payload_136 = (_zz_dataOut_payload_128_352 ? _zz_dataOut_payload_128_337 : _zz_dataOut_payload_128_321);
  assign _zz_dataOut_payload_128_354 = (_zz_dataOut_payload_128_323 < _zz_dataOut_payload_128_339);
  assign _zz_dataOut_payload_128_355 = (_zz_dataOut_payload_128_354 ? _zz_dataOut_payload_128_323 : _zz_dataOut_payload_128_339);
  assign _zz_dataOut_payload_136_1 = (_zz_dataOut_payload_128_354 ? _zz_dataOut_payload_128_339 : _zz_dataOut_payload_128_323);
  assign _zz_dataOut_payload_128_356 = (_zz_dataOut_payload_128_325 < _zz_dataOut_payload_128_341);
  assign _zz_dataOut_payload_128_357 = (_zz_dataOut_payload_128_356 ? _zz_dataOut_payload_128_325 : _zz_dataOut_payload_128_341);
  assign _zz_dataOut_payload_136_2 = (_zz_dataOut_payload_128_356 ? _zz_dataOut_payload_128_341 : _zz_dataOut_payload_128_325);
  assign _zz_dataOut_payload_128_358 = (_zz_dataOut_payload_128_327 < _zz_dataOut_payload_128_343);
  assign _zz_dataOut_payload_128_359 = (_zz_dataOut_payload_128_358 ? _zz_dataOut_payload_128_327 : _zz_dataOut_payload_128_343);
  assign _zz_dataOut_payload_136_3 = (_zz_dataOut_payload_128_358 ? _zz_dataOut_payload_128_343 : _zz_dataOut_payload_128_327);
  assign _zz_dataOut_payload_128_360 = (_zz_dataOut_payload_128_329 < _zz_dataOut_payload_128_345);
  assign _zz_dataOut_payload_128_361 = (_zz_dataOut_payload_128_360 ? _zz_dataOut_payload_128_329 : _zz_dataOut_payload_128_345);
  assign _zz_dataOut_payload_136_4 = (_zz_dataOut_payload_128_360 ? _zz_dataOut_payload_128_345 : _zz_dataOut_payload_128_329);
  assign _zz_dataOut_payload_128_362 = (_zz_dataOut_payload_128_331 < _zz_dataOut_payload_128_347);
  assign _zz_dataOut_payload_128_363 = (_zz_dataOut_payload_128_362 ? _zz_dataOut_payload_128_331 : _zz_dataOut_payload_128_347);
  assign _zz_dataOut_payload_136_5 = (_zz_dataOut_payload_128_362 ? _zz_dataOut_payload_128_347 : _zz_dataOut_payload_128_331);
  assign _zz_dataOut_payload_128_364 = (_zz_dataOut_payload_128_333 < _zz_dataOut_payload_128_349);
  assign _zz_dataOut_payload_128_365 = (_zz_dataOut_payload_128_364 ? _zz_dataOut_payload_128_333 : _zz_dataOut_payload_128_349);
  assign _zz_dataOut_payload_136_6 = (_zz_dataOut_payload_128_364 ? _zz_dataOut_payload_128_349 : _zz_dataOut_payload_128_333);
  assign _zz_dataOut_payload_128_366 = (_zz_dataOut_payload_128_335 < _zz_dataOut_payload_128_351);
  assign _zz_dataOut_payload_128_367 = (_zz_dataOut_payload_128_366 ? _zz_dataOut_payload_128_335 : _zz_dataOut_payload_128_351);
  assign _zz_dataOut_payload_136_7 = (_zz_dataOut_payload_128_366 ? _zz_dataOut_payload_128_351 : _zz_dataOut_payload_128_335);
  assign _zz_dataOut_payload_128_368 = (_zz_dataOut_payload_128_353 < _zz_dataOut_payload_128_361);
  assign _zz_dataOut_payload_128_369 = (_zz_dataOut_payload_128_368 ? _zz_dataOut_payload_128_353 : _zz_dataOut_payload_128_361);
  assign _zz_dataOut_payload_132 = (_zz_dataOut_payload_128_368 ? _zz_dataOut_payload_128_361 : _zz_dataOut_payload_128_353);
  assign _zz_dataOut_payload_128_370 = (_zz_dataOut_payload_128_355 < _zz_dataOut_payload_128_363);
  assign _zz_dataOut_payload_128_371 = (_zz_dataOut_payload_128_370 ? _zz_dataOut_payload_128_355 : _zz_dataOut_payload_128_363);
  assign _zz_dataOut_payload_132_1 = (_zz_dataOut_payload_128_370 ? _zz_dataOut_payload_128_363 : _zz_dataOut_payload_128_355);
  assign _zz_dataOut_payload_128_372 = (_zz_dataOut_payload_128_357 < _zz_dataOut_payload_128_365);
  assign _zz_dataOut_payload_128_373 = (_zz_dataOut_payload_128_372 ? _zz_dataOut_payload_128_357 : _zz_dataOut_payload_128_365);
  assign _zz_dataOut_payload_132_2 = (_zz_dataOut_payload_128_372 ? _zz_dataOut_payload_128_365 : _zz_dataOut_payload_128_357);
  assign _zz_dataOut_payload_128_374 = (_zz_dataOut_payload_128_359 < _zz_dataOut_payload_128_367);
  assign _zz_dataOut_payload_128_375 = (_zz_dataOut_payload_128_374 ? _zz_dataOut_payload_128_359 : _zz_dataOut_payload_128_367);
  assign _zz_dataOut_payload_132_3 = (_zz_dataOut_payload_128_374 ? _zz_dataOut_payload_128_367 : _zz_dataOut_payload_128_359);
  assign _zz_dataOut_payload_128_376 = (_zz_dataOut_payload_128_369 < _zz_dataOut_payload_128_373);
  assign _zz_dataOut_payload_128_377 = (_zz_dataOut_payload_128_376 ? _zz_dataOut_payload_128_369 : _zz_dataOut_payload_128_373);
  assign _zz_dataOut_payload_130 = (_zz_dataOut_payload_128_376 ? _zz_dataOut_payload_128_373 : _zz_dataOut_payload_128_369);
  assign _zz_dataOut_payload_128_378 = (_zz_dataOut_payload_128_371 < _zz_dataOut_payload_128_375);
  assign _zz_dataOut_payload_128_379 = (_zz_dataOut_payload_128_378 ? _zz_dataOut_payload_128_371 : _zz_dataOut_payload_128_375);
  assign _zz_dataOut_payload_130_1 = (_zz_dataOut_payload_128_378 ? _zz_dataOut_payload_128_375 : _zz_dataOut_payload_128_371);
  assign _zz_dataOut_payload_128_380 = (_zz_dataOut_payload_128_377 < _zz_dataOut_payload_128_379);
  assign _zz_dataOut_payload_130_2 = (_zz_dataOut_payload_130 < _zz_dataOut_payload_130_1);
  assign _zz_dataOut_payload_132_4 = (_zz_dataOut_payload_132 < _zz_dataOut_payload_132_2);
  assign _zz_dataOut_payload_132_5 = (_zz_dataOut_payload_132_4 ? _zz_dataOut_payload_132 : _zz_dataOut_payload_132_2);
  assign _zz_dataOut_payload_134 = (_zz_dataOut_payload_132_4 ? _zz_dataOut_payload_132_2 : _zz_dataOut_payload_132);
  assign _zz_dataOut_payload_132_6 = (_zz_dataOut_payload_132_1 < _zz_dataOut_payload_132_3);
  assign _zz_dataOut_payload_132_7 = (_zz_dataOut_payload_132_6 ? _zz_dataOut_payload_132_1 : _zz_dataOut_payload_132_3);
  assign _zz_dataOut_payload_134_1 = (_zz_dataOut_payload_132_6 ? _zz_dataOut_payload_132_3 : _zz_dataOut_payload_132_1);
  assign _zz_dataOut_payload_132_8 = (_zz_dataOut_payload_132_5 < _zz_dataOut_payload_132_7);
  assign _zz_dataOut_payload_134_2 = (_zz_dataOut_payload_134 < _zz_dataOut_payload_134_1);
  assign _zz_dataOut_payload_136_8 = (_zz_dataOut_payload_136 < _zz_dataOut_payload_136_4);
  assign _zz_dataOut_payload_136_9 = (_zz_dataOut_payload_136_8 ? _zz_dataOut_payload_136 : _zz_dataOut_payload_136_4);
  assign _zz_dataOut_payload_140 = (_zz_dataOut_payload_136_8 ? _zz_dataOut_payload_136_4 : _zz_dataOut_payload_136);
  assign _zz_dataOut_payload_136_10 = (_zz_dataOut_payload_136_1 < _zz_dataOut_payload_136_5);
  assign _zz_dataOut_payload_136_11 = (_zz_dataOut_payload_136_10 ? _zz_dataOut_payload_136_1 : _zz_dataOut_payload_136_5);
  assign _zz_dataOut_payload_140_1 = (_zz_dataOut_payload_136_10 ? _zz_dataOut_payload_136_5 : _zz_dataOut_payload_136_1);
  assign _zz_dataOut_payload_136_12 = (_zz_dataOut_payload_136_2 < _zz_dataOut_payload_136_6);
  assign _zz_dataOut_payload_136_13 = (_zz_dataOut_payload_136_12 ? _zz_dataOut_payload_136_2 : _zz_dataOut_payload_136_6);
  assign _zz_dataOut_payload_140_2 = (_zz_dataOut_payload_136_12 ? _zz_dataOut_payload_136_6 : _zz_dataOut_payload_136_2);
  assign _zz_dataOut_payload_136_14 = (_zz_dataOut_payload_136_3 < _zz_dataOut_payload_136_7);
  assign _zz_dataOut_payload_136_15 = (_zz_dataOut_payload_136_14 ? _zz_dataOut_payload_136_3 : _zz_dataOut_payload_136_7);
  assign _zz_dataOut_payload_140_3 = (_zz_dataOut_payload_136_14 ? _zz_dataOut_payload_136_7 : _zz_dataOut_payload_136_3);
  assign _zz_dataOut_payload_136_16 = (_zz_dataOut_payload_136_9 < _zz_dataOut_payload_136_13);
  assign _zz_dataOut_payload_136_17 = (_zz_dataOut_payload_136_16 ? _zz_dataOut_payload_136_9 : _zz_dataOut_payload_136_13);
  assign _zz_dataOut_payload_138 = (_zz_dataOut_payload_136_16 ? _zz_dataOut_payload_136_13 : _zz_dataOut_payload_136_9);
  assign _zz_dataOut_payload_136_18 = (_zz_dataOut_payload_136_11 < _zz_dataOut_payload_136_15);
  assign _zz_dataOut_payload_136_19 = (_zz_dataOut_payload_136_18 ? _zz_dataOut_payload_136_11 : _zz_dataOut_payload_136_15);
  assign _zz_dataOut_payload_138_1 = (_zz_dataOut_payload_136_18 ? _zz_dataOut_payload_136_15 : _zz_dataOut_payload_136_11);
  assign _zz_dataOut_payload_136_20 = (_zz_dataOut_payload_136_17 < _zz_dataOut_payload_136_19);
  assign _zz_dataOut_payload_138_2 = (_zz_dataOut_payload_138 < _zz_dataOut_payload_138_1);
  assign _zz_dataOut_payload_140_4 = (_zz_dataOut_payload_140 < _zz_dataOut_payload_140_2);
  assign _zz_dataOut_payload_140_5 = (_zz_dataOut_payload_140_4 ? _zz_dataOut_payload_140 : _zz_dataOut_payload_140_2);
  assign _zz_dataOut_payload_142 = (_zz_dataOut_payload_140_4 ? _zz_dataOut_payload_140_2 : _zz_dataOut_payload_140);
  assign _zz_dataOut_payload_140_6 = (_zz_dataOut_payload_140_1 < _zz_dataOut_payload_140_3);
  assign _zz_dataOut_payload_140_7 = (_zz_dataOut_payload_140_6 ? _zz_dataOut_payload_140_1 : _zz_dataOut_payload_140_3);
  assign _zz_dataOut_payload_142_1 = (_zz_dataOut_payload_140_6 ? _zz_dataOut_payload_140_3 : _zz_dataOut_payload_140_1);
  assign _zz_dataOut_payload_140_8 = (_zz_dataOut_payload_140_5 < _zz_dataOut_payload_140_7);
  assign _zz_dataOut_payload_142_2 = (_zz_dataOut_payload_142 < _zz_dataOut_payload_142_1);
  assign _zz_dataOut_payload_144_16 = (_zz_dataOut_payload_144 < _zz_dataOut_payload_144_8);
  assign _zz_dataOut_payload_144_17 = (_zz_dataOut_payload_144_16 ? _zz_dataOut_payload_144 : _zz_dataOut_payload_144_8);
  assign _zz_dataOut_payload_152 = (_zz_dataOut_payload_144_16 ? _zz_dataOut_payload_144_8 : _zz_dataOut_payload_144);
  assign _zz_dataOut_payload_144_18 = (_zz_dataOut_payload_144_1 < _zz_dataOut_payload_144_9);
  assign _zz_dataOut_payload_144_19 = (_zz_dataOut_payload_144_18 ? _zz_dataOut_payload_144_1 : _zz_dataOut_payload_144_9);
  assign _zz_dataOut_payload_152_1 = (_zz_dataOut_payload_144_18 ? _zz_dataOut_payload_144_9 : _zz_dataOut_payload_144_1);
  assign _zz_dataOut_payload_144_20 = (_zz_dataOut_payload_144_2 < _zz_dataOut_payload_144_10);
  assign _zz_dataOut_payload_144_21 = (_zz_dataOut_payload_144_20 ? _zz_dataOut_payload_144_2 : _zz_dataOut_payload_144_10);
  assign _zz_dataOut_payload_152_2 = (_zz_dataOut_payload_144_20 ? _zz_dataOut_payload_144_10 : _zz_dataOut_payload_144_2);
  assign _zz_dataOut_payload_144_22 = (_zz_dataOut_payload_144_3 < _zz_dataOut_payload_144_11);
  assign _zz_dataOut_payload_144_23 = (_zz_dataOut_payload_144_22 ? _zz_dataOut_payload_144_3 : _zz_dataOut_payload_144_11);
  assign _zz_dataOut_payload_152_3 = (_zz_dataOut_payload_144_22 ? _zz_dataOut_payload_144_11 : _zz_dataOut_payload_144_3);
  assign _zz_dataOut_payload_144_24 = (_zz_dataOut_payload_144_4 < _zz_dataOut_payload_144_12);
  assign _zz_dataOut_payload_144_25 = (_zz_dataOut_payload_144_24 ? _zz_dataOut_payload_144_4 : _zz_dataOut_payload_144_12);
  assign _zz_dataOut_payload_152_4 = (_zz_dataOut_payload_144_24 ? _zz_dataOut_payload_144_12 : _zz_dataOut_payload_144_4);
  assign _zz_dataOut_payload_144_26 = (_zz_dataOut_payload_144_5 < _zz_dataOut_payload_144_13);
  assign _zz_dataOut_payload_144_27 = (_zz_dataOut_payload_144_26 ? _zz_dataOut_payload_144_5 : _zz_dataOut_payload_144_13);
  assign _zz_dataOut_payload_152_5 = (_zz_dataOut_payload_144_26 ? _zz_dataOut_payload_144_13 : _zz_dataOut_payload_144_5);
  assign _zz_dataOut_payload_144_28 = (_zz_dataOut_payload_144_6 < _zz_dataOut_payload_144_14);
  assign _zz_dataOut_payload_144_29 = (_zz_dataOut_payload_144_28 ? _zz_dataOut_payload_144_6 : _zz_dataOut_payload_144_14);
  assign _zz_dataOut_payload_152_6 = (_zz_dataOut_payload_144_28 ? _zz_dataOut_payload_144_14 : _zz_dataOut_payload_144_6);
  assign _zz_dataOut_payload_144_30 = (_zz_dataOut_payload_144_7 < _zz_dataOut_payload_144_15);
  assign _zz_dataOut_payload_144_31 = (_zz_dataOut_payload_144_30 ? _zz_dataOut_payload_144_7 : _zz_dataOut_payload_144_15);
  assign _zz_dataOut_payload_152_7 = (_zz_dataOut_payload_144_30 ? _zz_dataOut_payload_144_15 : _zz_dataOut_payload_144_7);
  assign _zz_dataOut_payload_144_32 = (_zz_dataOut_payload_144_17 < _zz_dataOut_payload_144_25);
  assign _zz_dataOut_payload_144_33 = (_zz_dataOut_payload_144_32 ? _zz_dataOut_payload_144_17 : _zz_dataOut_payload_144_25);
  assign _zz_dataOut_payload_148 = (_zz_dataOut_payload_144_32 ? _zz_dataOut_payload_144_25 : _zz_dataOut_payload_144_17);
  assign _zz_dataOut_payload_144_34 = (_zz_dataOut_payload_144_19 < _zz_dataOut_payload_144_27);
  assign _zz_dataOut_payload_144_35 = (_zz_dataOut_payload_144_34 ? _zz_dataOut_payload_144_19 : _zz_dataOut_payload_144_27);
  assign _zz_dataOut_payload_148_1 = (_zz_dataOut_payload_144_34 ? _zz_dataOut_payload_144_27 : _zz_dataOut_payload_144_19);
  assign _zz_dataOut_payload_144_36 = (_zz_dataOut_payload_144_21 < _zz_dataOut_payload_144_29);
  assign _zz_dataOut_payload_144_37 = (_zz_dataOut_payload_144_36 ? _zz_dataOut_payload_144_21 : _zz_dataOut_payload_144_29);
  assign _zz_dataOut_payload_148_2 = (_zz_dataOut_payload_144_36 ? _zz_dataOut_payload_144_29 : _zz_dataOut_payload_144_21);
  assign _zz_dataOut_payload_144_38 = (_zz_dataOut_payload_144_23 < _zz_dataOut_payload_144_31);
  assign _zz_dataOut_payload_144_39 = (_zz_dataOut_payload_144_38 ? _zz_dataOut_payload_144_23 : _zz_dataOut_payload_144_31);
  assign _zz_dataOut_payload_148_3 = (_zz_dataOut_payload_144_38 ? _zz_dataOut_payload_144_31 : _zz_dataOut_payload_144_23);
  assign _zz_dataOut_payload_144_40 = (_zz_dataOut_payload_144_33 < _zz_dataOut_payload_144_37);
  assign _zz_dataOut_payload_144_41 = (_zz_dataOut_payload_144_40 ? _zz_dataOut_payload_144_33 : _zz_dataOut_payload_144_37);
  assign _zz_dataOut_payload_146 = (_zz_dataOut_payload_144_40 ? _zz_dataOut_payload_144_37 : _zz_dataOut_payload_144_33);
  assign _zz_dataOut_payload_144_42 = (_zz_dataOut_payload_144_35 < _zz_dataOut_payload_144_39);
  assign _zz_dataOut_payload_144_43 = (_zz_dataOut_payload_144_42 ? _zz_dataOut_payload_144_35 : _zz_dataOut_payload_144_39);
  assign _zz_dataOut_payload_146_1 = (_zz_dataOut_payload_144_42 ? _zz_dataOut_payload_144_39 : _zz_dataOut_payload_144_35);
  assign _zz_dataOut_payload_144_44 = (_zz_dataOut_payload_144_41 < _zz_dataOut_payload_144_43);
  assign _zz_dataOut_payload_146_2 = (_zz_dataOut_payload_146 < _zz_dataOut_payload_146_1);
  assign _zz_dataOut_payload_148_4 = (_zz_dataOut_payload_148 < _zz_dataOut_payload_148_2);
  assign _zz_dataOut_payload_148_5 = (_zz_dataOut_payload_148_4 ? _zz_dataOut_payload_148 : _zz_dataOut_payload_148_2);
  assign _zz_dataOut_payload_150 = (_zz_dataOut_payload_148_4 ? _zz_dataOut_payload_148_2 : _zz_dataOut_payload_148);
  assign _zz_dataOut_payload_148_6 = (_zz_dataOut_payload_148_1 < _zz_dataOut_payload_148_3);
  assign _zz_dataOut_payload_148_7 = (_zz_dataOut_payload_148_6 ? _zz_dataOut_payload_148_1 : _zz_dataOut_payload_148_3);
  assign _zz_dataOut_payload_150_1 = (_zz_dataOut_payload_148_6 ? _zz_dataOut_payload_148_3 : _zz_dataOut_payload_148_1);
  assign _zz_dataOut_payload_148_8 = (_zz_dataOut_payload_148_5 < _zz_dataOut_payload_148_7);
  assign _zz_dataOut_payload_150_2 = (_zz_dataOut_payload_150 < _zz_dataOut_payload_150_1);
  assign _zz_dataOut_payload_152_8 = (_zz_dataOut_payload_152 < _zz_dataOut_payload_152_4);
  assign _zz_dataOut_payload_152_9 = (_zz_dataOut_payload_152_8 ? _zz_dataOut_payload_152 : _zz_dataOut_payload_152_4);
  assign _zz_dataOut_payload_156 = (_zz_dataOut_payload_152_8 ? _zz_dataOut_payload_152_4 : _zz_dataOut_payload_152);
  assign _zz_dataOut_payload_152_10 = (_zz_dataOut_payload_152_1 < _zz_dataOut_payload_152_5);
  assign _zz_dataOut_payload_152_11 = (_zz_dataOut_payload_152_10 ? _zz_dataOut_payload_152_1 : _zz_dataOut_payload_152_5);
  assign _zz_dataOut_payload_156_1 = (_zz_dataOut_payload_152_10 ? _zz_dataOut_payload_152_5 : _zz_dataOut_payload_152_1);
  assign _zz_dataOut_payload_152_12 = (_zz_dataOut_payload_152_2 < _zz_dataOut_payload_152_6);
  assign _zz_dataOut_payload_152_13 = (_zz_dataOut_payload_152_12 ? _zz_dataOut_payload_152_2 : _zz_dataOut_payload_152_6);
  assign _zz_dataOut_payload_156_2 = (_zz_dataOut_payload_152_12 ? _zz_dataOut_payload_152_6 : _zz_dataOut_payload_152_2);
  assign _zz_dataOut_payload_152_14 = (_zz_dataOut_payload_152_3 < _zz_dataOut_payload_152_7);
  assign _zz_dataOut_payload_152_15 = (_zz_dataOut_payload_152_14 ? _zz_dataOut_payload_152_3 : _zz_dataOut_payload_152_7);
  assign _zz_dataOut_payload_156_3 = (_zz_dataOut_payload_152_14 ? _zz_dataOut_payload_152_7 : _zz_dataOut_payload_152_3);
  assign _zz_dataOut_payload_152_16 = (_zz_dataOut_payload_152_9 < _zz_dataOut_payload_152_13);
  assign _zz_dataOut_payload_152_17 = (_zz_dataOut_payload_152_16 ? _zz_dataOut_payload_152_9 : _zz_dataOut_payload_152_13);
  assign _zz_dataOut_payload_154 = (_zz_dataOut_payload_152_16 ? _zz_dataOut_payload_152_13 : _zz_dataOut_payload_152_9);
  assign _zz_dataOut_payload_152_18 = (_zz_dataOut_payload_152_11 < _zz_dataOut_payload_152_15);
  assign _zz_dataOut_payload_152_19 = (_zz_dataOut_payload_152_18 ? _zz_dataOut_payload_152_11 : _zz_dataOut_payload_152_15);
  assign _zz_dataOut_payload_154_1 = (_zz_dataOut_payload_152_18 ? _zz_dataOut_payload_152_15 : _zz_dataOut_payload_152_11);
  assign _zz_dataOut_payload_152_20 = (_zz_dataOut_payload_152_17 < _zz_dataOut_payload_152_19);
  assign _zz_dataOut_payload_154_2 = (_zz_dataOut_payload_154 < _zz_dataOut_payload_154_1);
  assign _zz_dataOut_payload_156_4 = (_zz_dataOut_payload_156 < _zz_dataOut_payload_156_2);
  assign _zz_dataOut_payload_156_5 = (_zz_dataOut_payload_156_4 ? _zz_dataOut_payload_156 : _zz_dataOut_payload_156_2);
  assign _zz_dataOut_payload_158 = (_zz_dataOut_payload_156_4 ? _zz_dataOut_payload_156_2 : _zz_dataOut_payload_156);
  assign _zz_dataOut_payload_156_6 = (_zz_dataOut_payload_156_1 < _zz_dataOut_payload_156_3);
  assign _zz_dataOut_payload_156_7 = (_zz_dataOut_payload_156_6 ? _zz_dataOut_payload_156_1 : _zz_dataOut_payload_156_3);
  assign _zz_dataOut_payload_158_1 = (_zz_dataOut_payload_156_6 ? _zz_dataOut_payload_156_3 : _zz_dataOut_payload_156_1);
  assign _zz_dataOut_payload_156_8 = (_zz_dataOut_payload_156_5 < _zz_dataOut_payload_156_7);
  assign _zz_dataOut_payload_158_2 = (_zz_dataOut_payload_158 < _zz_dataOut_payload_158_1);
  assign _zz_dataOut_payload_160_32 = (_zz_dataOut_payload_160 < _zz_dataOut_payload_160_16);
  assign _zz_dataOut_payload_160_33 = (_zz_dataOut_payload_160_32 ? _zz_dataOut_payload_160 : _zz_dataOut_payload_160_16);
  assign _zz_dataOut_payload_176 = (_zz_dataOut_payload_160_32 ? _zz_dataOut_payload_160_16 : _zz_dataOut_payload_160);
  assign _zz_dataOut_payload_160_34 = (_zz_dataOut_payload_160_1 < _zz_dataOut_payload_160_17);
  assign _zz_dataOut_payload_160_35 = (_zz_dataOut_payload_160_34 ? _zz_dataOut_payload_160_1 : _zz_dataOut_payload_160_17);
  assign _zz_dataOut_payload_176_1 = (_zz_dataOut_payload_160_34 ? _zz_dataOut_payload_160_17 : _zz_dataOut_payload_160_1);
  assign _zz_dataOut_payload_160_36 = (_zz_dataOut_payload_160_2 < _zz_dataOut_payload_160_18);
  assign _zz_dataOut_payload_160_37 = (_zz_dataOut_payload_160_36 ? _zz_dataOut_payload_160_2 : _zz_dataOut_payload_160_18);
  assign _zz_dataOut_payload_176_2 = (_zz_dataOut_payload_160_36 ? _zz_dataOut_payload_160_18 : _zz_dataOut_payload_160_2);
  assign _zz_dataOut_payload_160_38 = (_zz_dataOut_payload_160_3 < _zz_dataOut_payload_160_19);
  assign _zz_dataOut_payload_160_39 = (_zz_dataOut_payload_160_38 ? _zz_dataOut_payload_160_3 : _zz_dataOut_payload_160_19);
  assign _zz_dataOut_payload_176_3 = (_zz_dataOut_payload_160_38 ? _zz_dataOut_payload_160_19 : _zz_dataOut_payload_160_3);
  assign _zz_dataOut_payload_160_40 = (_zz_dataOut_payload_160_4 < _zz_dataOut_payload_160_20);
  assign _zz_dataOut_payload_160_41 = (_zz_dataOut_payload_160_40 ? _zz_dataOut_payload_160_4 : _zz_dataOut_payload_160_20);
  assign _zz_dataOut_payload_176_4 = (_zz_dataOut_payload_160_40 ? _zz_dataOut_payload_160_20 : _zz_dataOut_payload_160_4);
  assign _zz_dataOut_payload_160_42 = (_zz_dataOut_payload_160_5 < _zz_dataOut_payload_160_21);
  assign _zz_dataOut_payload_160_43 = (_zz_dataOut_payload_160_42 ? _zz_dataOut_payload_160_5 : _zz_dataOut_payload_160_21);
  assign _zz_dataOut_payload_176_5 = (_zz_dataOut_payload_160_42 ? _zz_dataOut_payload_160_21 : _zz_dataOut_payload_160_5);
  assign _zz_dataOut_payload_160_44 = (_zz_dataOut_payload_160_6 < _zz_dataOut_payload_160_22);
  assign _zz_dataOut_payload_160_45 = (_zz_dataOut_payload_160_44 ? _zz_dataOut_payload_160_6 : _zz_dataOut_payload_160_22);
  assign _zz_dataOut_payload_176_6 = (_zz_dataOut_payload_160_44 ? _zz_dataOut_payload_160_22 : _zz_dataOut_payload_160_6);
  assign _zz_dataOut_payload_160_46 = (_zz_dataOut_payload_160_7 < _zz_dataOut_payload_160_23);
  assign _zz_dataOut_payload_160_47 = (_zz_dataOut_payload_160_46 ? _zz_dataOut_payload_160_7 : _zz_dataOut_payload_160_23);
  assign _zz_dataOut_payload_176_7 = (_zz_dataOut_payload_160_46 ? _zz_dataOut_payload_160_23 : _zz_dataOut_payload_160_7);
  assign _zz_dataOut_payload_160_48 = (_zz_dataOut_payload_160_8 < _zz_dataOut_payload_160_24);
  assign _zz_dataOut_payload_160_49 = (_zz_dataOut_payload_160_48 ? _zz_dataOut_payload_160_8 : _zz_dataOut_payload_160_24);
  assign _zz_dataOut_payload_176_8 = (_zz_dataOut_payload_160_48 ? _zz_dataOut_payload_160_24 : _zz_dataOut_payload_160_8);
  assign _zz_dataOut_payload_160_50 = (_zz_dataOut_payload_160_9 < _zz_dataOut_payload_160_25);
  assign _zz_dataOut_payload_160_51 = (_zz_dataOut_payload_160_50 ? _zz_dataOut_payload_160_9 : _zz_dataOut_payload_160_25);
  assign _zz_dataOut_payload_176_9 = (_zz_dataOut_payload_160_50 ? _zz_dataOut_payload_160_25 : _zz_dataOut_payload_160_9);
  assign _zz_dataOut_payload_160_52 = (_zz_dataOut_payload_160_10 < _zz_dataOut_payload_160_26);
  assign _zz_dataOut_payload_160_53 = (_zz_dataOut_payload_160_52 ? _zz_dataOut_payload_160_10 : _zz_dataOut_payload_160_26);
  assign _zz_dataOut_payload_176_10 = (_zz_dataOut_payload_160_52 ? _zz_dataOut_payload_160_26 : _zz_dataOut_payload_160_10);
  assign _zz_dataOut_payload_160_54 = (_zz_dataOut_payload_160_11 < _zz_dataOut_payload_160_27);
  assign _zz_dataOut_payload_160_55 = (_zz_dataOut_payload_160_54 ? _zz_dataOut_payload_160_11 : _zz_dataOut_payload_160_27);
  assign _zz_dataOut_payload_176_11 = (_zz_dataOut_payload_160_54 ? _zz_dataOut_payload_160_27 : _zz_dataOut_payload_160_11);
  assign _zz_dataOut_payload_160_56 = (_zz_dataOut_payload_160_12 < _zz_dataOut_payload_160_28);
  assign _zz_dataOut_payload_160_57 = (_zz_dataOut_payload_160_56 ? _zz_dataOut_payload_160_12 : _zz_dataOut_payload_160_28);
  assign _zz_dataOut_payload_176_12 = (_zz_dataOut_payload_160_56 ? _zz_dataOut_payload_160_28 : _zz_dataOut_payload_160_12);
  assign _zz_dataOut_payload_160_58 = (_zz_dataOut_payload_160_13 < _zz_dataOut_payload_160_29);
  assign _zz_dataOut_payload_160_59 = (_zz_dataOut_payload_160_58 ? _zz_dataOut_payload_160_13 : _zz_dataOut_payload_160_29);
  assign _zz_dataOut_payload_176_13 = (_zz_dataOut_payload_160_58 ? _zz_dataOut_payload_160_29 : _zz_dataOut_payload_160_13);
  assign _zz_dataOut_payload_160_60 = (_zz_dataOut_payload_160_14 < _zz_dataOut_payload_160_30);
  assign _zz_dataOut_payload_160_61 = (_zz_dataOut_payload_160_60 ? _zz_dataOut_payload_160_14 : _zz_dataOut_payload_160_30);
  assign _zz_dataOut_payload_176_14 = (_zz_dataOut_payload_160_60 ? _zz_dataOut_payload_160_30 : _zz_dataOut_payload_160_14);
  assign _zz_dataOut_payload_160_62 = (_zz_dataOut_payload_160_15 < _zz_dataOut_payload_160_31);
  assign _zz_dataOut_payload_160_63 = (_zz_dataOut_payload_160_62 ? _zz_dataOut_payload_160_15 : _zz_dataOut_payload_160_31);
  assign _zz_dataOut_payload_176_15 = (_zz_dataOut_payload_160_62 ? _zz_dataOut_payload_160_31 : _zz_dataOut_payload_160_15);
  assign _zz_dataOut_payload_160_64 = (_zz_dataOut_payload_160_33 < _zz_dataOut_payload_160_49);
  assign _zz_dataOut_payload_160_65 = (_zz_dataOut_payload_160_64 ? _zz_dataOut_payload_160_33 : _zz_dataOut_payload_160_49);
  assign _zz_dataOut_payload_168 = (_zz_dataOut_payload_160_64 ? _zz_dataOut_payload_160_49 : _zz_dataOut_payload_160_33);
  assign _zz_dataOut_payload_160_66 = (_zz_dataOut_payload_160_35 < _zz_dataOut_payload_160_51);
  assign _zz_dataOut_payload_160_67 = (_zz_dataOut_payload_160_66 ? _zz_dataOut_payload_160_35 : _zz_dataOut_payload_160_51);
  assign _zz_dataOut_payload_168_1 = (_zz_dataOut_payload_160_66 ? _zz_dataOut_payload_160_51 : _zz_dataOut_payload_160_35);
  assign _zz_dataOut_payload_160_68 = (_zz_dataOut_payload_160_37 < _zz_dataOut_payload_160_53);
  assign _zz_dataOut_payload_160_69 = (_zz_dataOut_payload_160_68 ? _zz_dataOut_payload_160_37 : _zz_dataOut_payload_160_53);
  assign _zz_dataOut_payload_168_2 = (_zz_dataOut_payload_160_68 ? _zz_dataOut_payload_160_53 : _zz_dataOut_payload_160_37);
  assign _zz_dataOut_payload_160_70 = (_zz_dataOut_payload_160_39 < _zz_dataOut_payload_160_55);
  assign _zz_dataOut_payload_160_71 = (_zz_dataOut_payload_160_70 ? _zz_dataOut_payload_160_39 : _zz_dataOut_payload_160_55);
  assign _zz_dataOut_payload_168_3 = (_zz_dataOut_payload_160_70 ? _zz_dataOut_payload_160_55 : _zz_dataOut_payload_160_39);
  assign _zz_dataOut_payload_160_72 = (_zz_dataOut_payload_160_41 < _zz_dataOut_payload_160_57);
  assign _zz_dataOut_payload_160_73 = (_zz_dataOut_payload_160_72 ? _zz_dataOut_payload_160_41 : _zz_dataOut_payload_160_57);
  assign _zz_dataOut_payload_168_4 = (_zz_dataOut_payload_160_72 ? _zz_dataOut_payload_160_57 : _zz_dataOut_payload_160_41);
  assign _zz_dataOut_payload_160_74 = (_zz_dataOut_payload_160_43 < _zz_dataOut_payload_160_59);
  assign _zz_dataOut_payload_160_75 = (_zz_dataOut_payload_160_74 ? _zz_dataOut_payload_160_43 : _zz_dataOut_payload_160_59);
  assign _zz_dataOut_payload_168_5 = (_zz_dataOut_payload_160_74 ? _zz_dataOut_payload_160_59 : _zz_dataOut_payload_160_43);
  assign _zz_dataOut_payload_160_76 = (_zz_dataOut_payload_160_45 < _zz_dataOut_payload_160_61);
  assign _zz_dataOut_payload_160_77 = (_zz_dataOut_payload_160_76 ? _zz_dataOut_payload_160_45 : _zz_dataOut_payload_160_61);
  assign _zz_dataOut_payload_168_6 = (_zz_dataOut_payload_160_76 ? _zz_dataOut_payload_160_61 : _zz_dataOut_payload_160_45);
  assign _zz_dataOut_payload_160_78 = (_zz_dataOut_payload_160_47 < _zz_dataOut_payload_160_63);
  assign _zz_dataOut_payload_160_79 = (_zz_dataOut_payload_160_78 ? _zz_dataOut_payload_160_47 : _zz_dataOut_payload_160_63);
  assign _zz_dataOut_payload_168_7 = (_zz_dataOut_payload_160_78 ? _zz_dataOut_payload_160_63 : _zz_dataOut_payload_160_47);
  assign _zz_dataOut_payload_160_80 = (_zz_dataOut_payload_160_65 < _zz_dataOut_payload_160_73);
  assign _zz_dataOut_payload_160_81 = (_zz_dataOut_payload_160_80 ? _zz_dataOut_payload_160_65 : _zz_dataOut_payload_160_73);
  assign _zz_dataOut_payload_164 = (_zz_dataOut_payload_160_80 ? _zz_dataOut_payload_160_73 : _zz_dataOut_payload_160_65);
  assign _zz_dataOut_payload_160_82 = (_zz_dataOut_payload_160_67 < _zz_dataOut_payload_160_75);
  assign _zz_dataOut_payload_160_83 = (_zz_dataOut_payload_160_82 ? _zz_dataOut_payload_160_67 : _zz_dataOut_payload_160_75);
  assign _zz_dataOut_payload_164_1 = (_zz_dataOut_payload_160_82 ? _zz_dataOut_payload_160_75 : _zz_dataOut_payload_160_67);
  assign _zz_dataOut_payload_160_84 = (_zz_dataOut_payload_160_69 < _zz_dataOut_payload_160_77);
  assign _zz_dataOut_payload_160_85 = (_zz_dataOut_payload_160_84 ? _zz_dataOut_payload_160_69 : _zz_dataOut_payload_160_77);
  assign _zz_dataOut_payload_164_2 = (_zz_dataOut_payload_160_84 ? _zz_dataOut_payload_160_77 : _zz_dataOut_payload_160_69);
  assign _zz_dataOut_payload_160_86 = (_zz_dataOut_payload_160_71 < _zz_dataOut_payload_160_79);
  assign _zz_dataOut_payload_160_87 = (_zz_dataOut_payload_160_86 ? _zz_dataOut_payload_160_71 : _zz_dataOut_payload_160_79);
  assign _zz_dataOut_payload_164_3 = (_zz_dataOut_payload_160_86 ? _zz_dataOut_payload_160_79 : _zz_dataOut_payload_160_71);
  assign _zz_dataOut_payload_160_88 = (_zz_dataOut_payload_160_81 < _zz_dataOut_payload_160_85);
  assign _zz_dataOut_payload_160_89 = (_zz_dataOut_payload_160_88 ? _zz_dataOut_payload_160_81 : _zz_dataOut_payload_160_85);
  assign _zz_dataOut_payload_162 = (_zz_dataOut_payload_160_88 ? _zz_dataOut_payload_160_85 : _zz_dataOut_payload_160_81);
  assign _zz_dataOut_payload_160_90 = (_zz_dataOut_payload_160_83 < _zz_dataOut_payload_160_87);
  assign _zz_dataOut_payload_160_91 = (_zz_dataOut_payload_160_90 ? _zz_dataOut_payload_160_83 : _zz_dataOut_payload_160_87);
  assign _zz_dataOut_payload_162_1 = (_zz_dataOut_payload_160_90 ? _zz_dataOut_payload_160_87 : _zz_dataOut_payload_160_83);
  assign _zz_dataOut_payload_160_92 = (_zz_dataOut_payload_160_89 < _zz_dataOut_payload_160_91);
  assign _zz_dataOut_payload_162_2 = (_zz_dataOut_payload_162 < _zz_dataOut_payload_162_1);
  assign _zz_dataOut_payload_164_4 = (_zz_dataOut_payload_164 < _zz_dataOut_payload_164_2);
  assign _zz_dataOut_payload_164_5 = (_zz_dataOut_payload_164_4 ? _zz_dataOut_payload_164 : _zz_dataOut_payload_164_2);
  assign _zz_dataOut_payload_166 = (_zz_dataOut_payload_164_4 ? _zz_dataOut_payload_164_2 : _zz_dataOut_payload_164);
  assign _zz_dataOut_payload_164_6 = (_zz_dataOut_payload_164_1 < _zz_dataOut_payload_164_3);
  assign _zz_dataOut_payload_164_7 = (_zz_dataOut_payload_164_6 ? _zz_dataOut_payload_164_1 : _zz_dataOut_payload_164_3);
  assign _zz_dataOut_payload_166_1 = (_zz_dataOut_payload_164_6 ? _zz_dataOut_payload_164_3 : _zz_dataOut_payload_164_1);
  assign _zz_dataOut_payload_164_8 = (_zz_dataOut_payload_164_5 < _zz_dataOut_payload_164_7);
  assign _zz_dataOut_payload_166_2 = (_zz_dataOut_payload_166 < _zz_dataOut_payload_166_1);
  assign _zz_dataOut_payload_168_8 = (_zz_dataOut_payload_168 < _zz_dataOut_payload_168_4);
  assign _zz_dataOut_payload_168_9 = (_zz_dataOut_payload_168_8 ? _zz_dataOut_payload_168 : _zz_dataOut_payload_168_4);
  assign _zz_dataOut_payload_172 = (_zz_dataOut_payload_168_8 ? _zz_dataOut_payload_168_4 : _zz_dataOut_payload_168);
  assign _zz_dataOut_payload_168_10 = (_zz_dataOut_payload_168_1 < _zz_dataOut_payload_168_5);
  assign _zz_dataOut_payload_168_11 = (_zz_dataOut_payload_168_10 ? _zz_dataOut_payload_168_1 : _zz_dataOut_payload_168_5);
  assign _zz_dataOut_payload_172_1 = (_zz_dataOut_payload_168_10 ? _zz_dataOut_payload_168_5 : _zz_dataOut_payload_168_1);
  assign _zz_dataOut_payload_168_12 = (_zz_dataOut_payload_168_2 < _zz_dataOut_payload_168_6);
  assign _zz_dataOut_payload_168_13 = (_zz_dataOut_payload_168_12 ? _zz_dataOut_payload_168_2 : _zz_dataOut_payload_168_6);
  assign _zz_dataOut_payload_172_2 = (_zz_dataOut_payload_168_12 ? _zz_dataOut_payload_168_6 : _zz_dataOut_payload_168_2);
  assign _zz_dataOut_payload_168_14 = (_zz_dataOut_payload_168_3 < _zz_dataOut_payload_168_7);
  assign _zz_dataOut_payload_168_15 = (_zz_dataOut_payload_168_14 ? _zz_dataOut_payload_168_3 : _zz_dataOut_payload_168_7);
  assign _zz_dataOut_payload_172_3 = (_zz_dataOut_payload_168_14 ? _zz_dataOut_payload_168_7 : _zz_dataOut_payload_168_3);
  assign _zz_dataOut_payload_168_16 = (_zz_dataOut_payload_168_9 < _zz_dataOut_payload_168_13);
  assign _zz_dataOut_payload_168_17 = (_zz_dataOut_payload_168_16 ? _zz_dataOut_payload_168_9 : _zz_dataOut_payload_168_13);
  assign _zz_dataOut_payload_170 = (_zz_dataOut_payload_168_16 ? _zz_dataOut_payload_168_13 : _zz_dataOut_payload_168_9);
  assign _zz_dataOut_payload_168_18 = (_zz_dataOut_payload_168_11 < _zz_dataOut_payload_168_15);
  assign _zz_dataOut_payload_168_19 = (_zz_dataOut_payload_168_18 ? _zz_dataOut_payload_168_11 : _zz_dataOut_payload_168_15);
  assign _zz_dataOut_payload_170_1 = (_zz_dataOut_payload_168_18 ? _zz_dataOut_payload_168_15 : _zz_dataOut_payload_168_11);
  assign _zz_dataOut_payload_168_20 = (_zz_dataOut_payload_168_17 < _zz_dataOut_payload_168_19);
  assign _zz_dataOut_payload_170_2 = (_zz_dataOut_payload_170 < _zz_dataOut_payload_170_1);
  assign _zz_dataOut_payload_172_4 = (_zz_dataOut_payload_172 < _zz_dataOut_payload_172_2);
  assign _zz_dataOut_payload_172_5 = (_zz_dataOut_payload_172_4 ? _zz_dataOut_payload_172 : _zz_dataOut_payload_172_2);
  assign _zz_dataOut_payload_174 = (_zz_dataOut_payload_172_4 ? _zz_dataOut_payload_172_2 : _zz_dataOut_payload_172);
  assign _zz_dataOut_payload_172_6 = (_zz_dataOut_payload_172_1 < _zz_dataOut_payload_172_3);
  assign _zz_dataOut_payload_172_7 = (_zz_dataOut_payload_172_6 ? _zz_dataOut_payload_172_1 : _zz_dataOut_payload_172_3);
  assign _zz_dataOut_payload_174_1 = (_zz_dataOut_payload_172_6 ? _zz_dataOut_payload_172_3 : _zz_dataOut_payload_172_1);
  assign _zz_dataOut_payload_172_8 = (_zz_dataOut_payload_172_5 < _zz_dataOut_payload_172_7);
  assign _zz_dataOut_payload_174_2 = (_zz_dataOut_payload_174 < _zz_dataOut_payload_174_1);
  assign _zz_dataOut_payload_176_16 = (_zz_dataOut_payload_176 < _zz_dataOut_payload_176_8);
  assign _zz_dataOut_payload_176_17 = (_zz_dataOut_payload_176_16 ? _zz_dataOut_payload_176 : _zz_dataOut_payload_176_8);
  assign _zz_dataOut_payload_184 = (_zz_dataOut_payload_176_16 ? _zz_dataOut_payload_176_8 : _zz_dataOut_payload_176);
  assign _zz_dataOut_payload_176_18 = (_zz_dataOut_payload_176_1 < _zz_dataOut_payload_176_9);
  assign _zz_dataOut_payload_176_19 = (_zz_dataOut_payload_176_18 ? _zz_dataOut_payload_176_1 : _zz_dataOut_payload_176_9);
  assign _zz_dataOut_payload_184_1 = (_zz_dataOut_payload_176_18 ? _zz_dataOut_payload_176_9 : _zz_dataOut_payload_176_1);
  assign _zz_dataOut_payload_176_20 = (_zz_dataOut_payload_176_2 < _zz_dataOut_payload_176_10);
  assign _zz_dataOut_payload_176_21 = (_zz_dataOut_payload_176_20 ? _zz_dataOut_payload_176_2 : _zz_dataOut_payload_176_10);
  assign _zz_dataOut_payload_184_2 = (_zz_dataOut_payload_176_20 ? _zz_dataOut_payload_176_10 : _zz_dataOut_payload_176_2);
  assign _zz_dataOut_payload_176_22 = (_zz_dataOut_payload_176_3 < _zz_dataOut_payload_176_11);
  assign _zz_dataOut_payload_176_23 = (_zz_dataOut_payload_176_22 ? _zz_dataOut_payload_176_3 : _zz_dataOut_payload_176_11);
  assign _zz_dataOut_payload_184_3 = (_zz_dataOut_payload_176_22 ? _zz_dataOut_payload_176_11 : _zz_dataOut_payload_176_3);
  assign _zz_dataOut_payload_176_24 = (_zz_dataOut_payload_176_4 < _zz_dataOut_payload_176_12);
  assign _zz_dataOut_payload_176_25 = (_zz_dataOut_payload_176_24 ? _zz_dataOut_payload_176_4 : _zz_dataOut_payload_176_12);
  assign _zz_dataOut_payload_184_4 = (_zz_dataOut_payload_176_24 ? _zz_dataOut_payload_176_12 : _zz_dataOut_payload_176_4);
  assign _zz_dataOut_payload_176_26 = (_zz_dataOut_payload_176_5 < _zz_dataOut_payload_176_13);
  assign _zz_dataOut_payload_176_27 = (_zz_dataOut_payload_176_26 ? _zz_dataOut_payload_176_5 : _zz_dataOut_payload_176_13);
  assign _zz_dataOut_payload_184_5 = (_zz_dataOut_payload_176_26 ? _zz_dataOut_payload_176_13 : _zz_dataOut_payload_176_5);
  assign _zz_dataOut_payload_176_28 = (_zz_dataOut_payload_176_6 < _zz_dataOut_payload_176_14);
  assign _zz_dataOut_payload_176_29 = (_zz_dataOut_payload_176_28 ? _zz_dataOut_payload_176_6 : _zz_dataOut_payload_176_14);
  assign _zz_dataOut_payload_184_6 = (_zz_dataOut_payload_176_28 ? _zz_dataOut_payload_176_14 : _zz_dataOut_payload_176_6);
  assign _zz_dataOut_payload_176_30 = (_zz_dataOut_payload_176_7 < _zz_dataOut_payload_176_15);
  assign _zz_dataOut_payload_176_31 = (_zz_dataOut_payload_176_30 ? _zz_dataOut_payload_176_7 : _zz_dataOut_payload_176_15);
  assign _zz_dataOut_payload_184_7 = (_zz_dataOut_payload_176_30 ? _zz_dataOut_payload_176_15 : _zz_dataOut_payload_176_7);
  assign _zz_dataOut_payload_176_32 = (_zz_dataOut_payload_176_17 < _zz_dataOut_payload_176_25);
  assign _zz_dataOut_payload_176_33 = (_zz_dataOut_payload_176_32 ? _zz_dataOut_payload_176_17 : _zz_dataOut_payload_176_25);
  assign _zz_dataOut_payload_180 = (_zz_dataOut_payload_176_32 ? _zz_dataOut_payload_176_25 : _zz_dataOut_payload_176_17);
  assign _zz_dataOut_payload_176_34 = (_zz_dataOut_payload_176_19 < _zz_dataOut_payload_176_27);
  assign _zz_dataOut_payload_176_35 = (_zz_dataOut_payload_176_34 ? _zz_dataOut_payload_176_19 : _zz_dataOut_payload_176_27);
  assign _zz_dataOut_payload_180_1 = (_zz_dataOut_payload_176_34 ? _zz_dataOut_payload_176_27 : _zz_dataOut_payload_176_19);
  assign _zz_dataOut_payload_176_36 = (_zz_dataOut_payload_176_21 < _zz_dataOut_payload_176_29);
  assign _zz_dataOut_payload_176_37 = (_zz_dataOut_payload_176_36 ? _zz_dataOut_payload_176_21 : _zz_dataOut_payload_176_29);
  assign _zz_dataOut_payload_180_2 = (_zz_dataOut_payload_176_36 ? _zz_dataOut_payload_176_29 : _zz_dataOut_payload_176_21);
  assign _zz_dataOut_payload_176_38 = (_zz_dataOut_payload_176_23 < _zz_dataOut_payload_176_31);
  assign _zz_dataOut_payload_176_39 = (_zz_dataOut_payload_176_38 ? _zz_dataOut_payload_176_23 : _zz_dataOut_payload_176_31);
  assign _zz_dataOut_payload_180_3 = (_zz_dataOut_payload_176_38 ? _zz_dataOut_payload_176_31 : _zz_dataOut_payload_176_23);
  assign _zz_dataOut_payload_176_40 = (_zz_dataOut_payload_176_33 < _zz_dataOut_payload_176_37);
  assign _zz_dataOut_payload_176_41 = (_zz_dataOut_payload_176_40 ? _zz_dataOut_payload_176_33 : _zz_dataOut_payload_176_37);
  assign _zz_dataOut_payload_178 = (_zz_dataOut_payload_176_40 ? _zz_dataOut_payload_176_37 : _zz_dataOut_payload_176_33);
  assign _zz_dataOut_payload_176_42 = (_zz_dataOut_payload_176_35 < _zz_dataOut_payload_176_39);
  assign _zz_dataOut_payload_176_43 = (_zz_dataOut_payload_176_42 ? _zz_dataOut_payload_176_35 : _zz_dataOut_payload_176_39);
  assign _zz_dataOut_payload_178_1 = (_zz_dataOut_payload_176_42 ? _zz_dataOut_payload_176_39 : _zz_dataOut_payload_176_35);
  assign _zz_dataOut_payload_176_44 = (_zz_dataOut_payload_176_41 < _zz_dataOut_payload_176_43);
  assign _zz_dataOut_payload_178_2 = (_zz_dataOut_payload_178 < _zz_dataOut_payload_178_1);
  assign _zz_dataOut_payload_180_4 = (_zz_dataOut_payload_180 < _zz_dataOut_payload_180_2);
  assign _zz_dataOut_payload_180_5 = (_zz_dataOut_payload_180_4 ? _zz_dataOut_payload_180 : _zz_dataOut_payload_180_2);
  assign _zz_dataOut_payload_182 = (_zz_dataOut_payload_180_4 ? _zz_dataOut_payload_180_2 : _zz_dataOut_payload_180);
  assign _zz_dataOut_payload_180_6 = (_zz_dataOut_payload_180_1 < _zz_dataOut_payload_180_3);
  assign _zz_dataOut_payload_180_7 = (_zz_dataOut_payload_180_6 ? _zz_dataOut_payload_180_1 : _zz_dataOut_payload_180_3);
  assign _zz_dataOut_payload_182_1 = (_zz_dataOut_payload_180_6 ? _zz_dataOut_payload_180_3 : _zz_dataOut_payload_180_1);
  assign _zz_dataOut_payload_180_8 = (_zz_dataOut_payload_180_5 < _zz_dataOut_payload_180_7);
  assign _zz_dataOut_payload_182_2 = (_zz_dataOut_payload_182 < _zz_dataOut_payload_182_1);
  assign _zz_dataOut_payload_184_8 = (_zz_dataOut_payload_184 < _zz_dataOut_payload_184_4);
  assign _zz_dataOut_payload_184_9 = (_zz_dataOut_payload_184_8 ? _zz_dataOut_payload_184 : _zz_dataOut_payload_184_4);
  assign _zz_dataOut_payload_188 = (_zz_dataOut_payload_184_8 ? _zz_dataOut_payload_184_4 : _zz_dataOut_payload_184);
  assign _zz_dataOut_payload_184_10 = (_zz_dataOut_payload_184_1 < _zz_dataOut_payload_184_5);
  assign _zz_dataOut_payload_184_11 = (_zz_dataOut_payload_184_10 ? _zz_dataOut_payload_184_1 : _zz_dataOut_payload_184_5);
  assign _zz_dataOut_payload_188_1 = (_zz_dataOut_payload_184_10 ? _zz_dataOut_payload_184_5 : _zz_dataOut_payload_184_1);
  assign _zz_dataOut_payload_184_12 = (_zz_dataOut_payload_184_2 < _zz_dataOut_payload_184_6);
  assign _zz_dataOut_payload_184_13 = (_zz_dataOut_payload_184_12 ? _zz_dataOut_payload_184_2 : _zz_dataOut_payload_184_6);
  assign _zz_dataOut_payload_188_2 = (_zz_dataOut_payload_184_12 ? _zz_dataOut_payload_184_6 : _zz_dataOut_payload_184_2);
  assign _zz_dataOut_payload_184_14 = (_zz_dataOut_payload_184_3 < _zz_dataOut_payload_184_7);
  assign _zz_dataOut_payload_184_15 = (_zz_dataOut_payload_184_14 ? _zz_dataOut_payload_184_3 : _zz_dataOut_payload_184_7);
  assign _zz_dataOut_payload_188_3 = (_zz_dataOut_payload_184_14 ? _zz_dataOut_payload_184_7 : _zz_dataOut_payload_184_3);
  assign _zz_dataOut_payload_184_16 = (_zz_dataOut_payload_184_9 < _zz_dataOut_payload_184_13);
  assign _zz_dataOut_payload_184_17 = (_zz_dataOut_payload_184_16 ? _zz_dataOut_payload_184_9 : _zz_dataOut_payload_184_13);
  assign _zz_dataOut_payload_186 = (_zz_dataOut_payload_184_16 ? _zz_dataOut_payload_184_13 : _zz_dataOut_payload_184_9);
  assign _zz_dataOut_payload_184_18 = (_zz_dataOut_payload_184_11 < _zz_dataOut_payload_184_15);
  assign _zz_dataOut_payload_184_19 = (_zz_dataOut_payload_184_18 ? _zz_dataOut_payload_184_11 : _zz_dataOut_payload_184_15);
  assign _zz_dataOut_payload_186_1 = (_zz_dataOut_payload_184_18 ? _zz_dataOut_payload_184_15 : _zz_dataOut_payload_184_11);
  assign _zz_dataOut_payload_184_20 = (_zz_dataOut_payload_184_17 < _zz_dataOut_payload_184_19);
  assign _zz_dataOut_payload_186_2 = (_zz_dataOut_payload_186 < _zz_dataOut_payload_186_1);
  assign _zz_dataOut_payload_188_4 = (_zz_dataOut_payload_188 < _zz_dataOut_payload_188_2);
  assign _zz_dataOut_payload_188_5 = (_zz_dataOut_payload_188_4 ? _zz_dataOut_payload_188 : _zz_dataOut_payload_188_2);
  assign _zz_dataOut_payload_190 = (_zz_dataOut_payload_188_4 ? _zz_dataOut_payload_188_2 : _zz_dataOut_payload_188);
  assign _zz_dataOut_payload_188_6 = (_zz_dataOut_payload_188_1 < _zz_dataOut_payload_188_3);
  assign _zz_dataOut_payload_188_7 = (_zz_dataOut_payload_188_6 ? _zz_dataOut_payload_188_1 : _zz_dataOut_payload_188_3);
  assign _zz_dataOut_payload_190_1 = (_zz_dataOut_payload_188_6 ? _zz_dataOut_payload_188_3 : _zz_dataOut_payload_188_1);
  assign _zz_dataOut_payload_188_8 = (_zz_dataOut_payload_188_5 < _zz_dataOut_payload_188_7);
  assign _zz_dataOut_payload_190_2 = (_zz_dataOut_payload_190 < _zz_dataOut_payload_190_1);
  assign _zz_dataOut_payload_192_64 = (_zz_dataOut_payload_192 < _zz_dataOut_payload_192_32);
  assign _zz_dataOut_payload_192_65 = (_zz_dataOut_payload_192_64 ? _zz_dataOut_payload_192 : _zz_dataOut_payload_192_32);
  assign _zz_dataOut_payload_224 = (_zz_dataOut_payload_192_64 ? _zz_dataOut_payload_192_32 : _zz_dataOut_payload_192);
  assign _zz_dataOut_payload_192_66 = (_zz_dataOut_payload_192_1 < _zz_dataOut_payload_192_33);
  assign _zz_dataOut_payload_192_67 = (_zz_dataOut_payload_192_66 ? _zz_dataOut_payload_192_1 : _zz_dataOut_payload_192_33);
  assign _zz_dataOut_payload_224_1 = (_zz_dataOut_payload_192_66 ? _zz_dataOut_payload_192_33 : _zz_dataOut_payload_192_1);
  assign _zz_dataOut_payload_192_68 = (_zz_dataOut_payload_192_2 < _zz_dataOut_payload_192_34);
  assign _zz_dataOut_payload_192_69 = (_zz_dataOut_payload_192_68 ? _zz_dataOut_payload_192_2 : _zz_dataOut_payload_192_34);
  assign _zz_dataOut_payload_224_2 = (_zz_dataOut_payload_192_68 ? _zz_dataOut_payload_192_34 : _zz_dataOut_payload_192_2);
  assign _zz_dataOut_payload_192_70 = (_zz_dataOut_payload_192_3 < _zz_dataOut_payload_192_35);
  assign _zz_dataOut_payload_192_71 = (_zz_dataOut_payload_192_70 ? _zz_dataOut_payload_192_3 : _zz_dataOut_payload_192_35);
  assign _zz_dataOut_payload_224_3 = (_zz_dataOut_payload_192_70 ? _zz_dataOut_payload_192_35 : _zz_dataOut_payload_192_3);
  assign _zz_dataOut_payload_192_72 = (_zz_dataOut_payload_192_4 < _zz_dataOut_payload_192_36);
  assign _zz_dataOut_payload_192_73 = (_zz_dataOut_payload_192_72 ? _zz_dataOut_payload_192_4 : _zz_dataOut_payload_192_36);
  assign _zz_dataOut_payload_224_4 = (_zz_dataOut_payload_192_72 ? _zz_dataOut_payload_192_36 : _zz_dataOut_payload_192_4);
  assign _zz_dataOut_payload_192_74 = (_zz_dataOut_payload_192_5 < _zz_dataOut_payload_192_37);
  assign _zz_dataOut_payload_192_75 = (_zz_dataOut_payload_192_74 ? _zz_dataOut_payload_192_5 : _zz_dataOut_payload_192_37);
  assign _zz_dataOut_payload_224_5 = (_zz_dataOut_payload_192_74 ? _zz_dataOut_payload_192_37 : _zz_dataOut_payload_192_5);
  assign _zz_dataOut_payload_192_76 = (_zz_dataOut_payload_192_6 < _zz_dataOut_payload_192_38);
  assign _zz_dataOut_payload_192_77 = (_zz_dataOut_payload_192_76 ? _zz_dataOut_payload_192_6 : _zz_dataOut_payload_192_38);
  assign _zz_dataOut_payload_224_6 = (_zz_dataOut_payload_192_76 ? _zz_dataOut_payload_192_38 : _zz_dataOut_payload_192_6);
  assign _zz_dataOut_payload_192_78 = (_zz_dataOut_payload_192_7 < _zz_dataOut_payload_192_39);
  assign _zz_dataOut_payload_192_79 = (_zz_dataOut_payload_192_78 ? _zz_dataOut_payload_192_7 : _zz_dataOut_payload_192_39);
  assign _zz_dataOut_payload_224_7 = (_zz_dataOut_payload_192_78 ? _zz_dataOut_payload_192_39 : _zz_dataOut_payload_192_7);
  assign _zz_dataOut_payload_192_80 = (_zz_dataOut_payload_192_8 < _zz_dataOut_payload_192_40);
  assign _zz_dataOut_payload_192_81 = (_zz_dataOut_payload_192_80 ? _zz_dataOut_payload_192_8 : _zz_dataOut_payload_192_40);
  assign _zz_dataOut_payload_224_8 = (_zz_dataOut_payload_192_80 ? _zz_dataOut_payload_192_40 : _zz_dataOut_payload_192_8);
  assign _zz_dataOut_payload_192_82 = (_zz_dataOut_payload_192_9 < _zz_dataOut_payload_192_41);
  assign _zz_dataOut_payload_192_83 = (_zz_dataOut_payload_192_82 ? _zz_dataOut_payload_192_9 : _zz_dataOut_payload_192_41);
  assign _zz_dataOut_payload_224_9 = (_zz_dataOut_payload_192_82 ? _zz_dataOut_payload_192_41 : _zz_dataOut_payload_192_9);
  assign _zz_dataOut_payload_192_84 = (_zz_dataOut_payload_192_10 < _zz_dataOut_payload_192_42);
  assign _zz_dataOut_payload_192_85 = (_zz_dataOut_payload_192_84 ? _zz_dataOut_payload_192_10 : _zz_dataOut_payload_192_42);
  assign _zz_dataOut_payload_224_10 = (_zz_dataOut_payload_192_84 ? _zz_dataOut_payload_192_42 : _zz_dataOut_payload_192_10);
  assign _zz_dataOut_payload_192_86 = (_zz_dataOut_payload_192_11 < _zz_dataOut_payload_192_43);
  assign _zz_dataOut_payload_192_87 = (_zz_dataOut_payload_192_86 ? _zz_dataOut_payload_192_11 : _zz_dataOut_payload_192_43);
  assign _zz_dataOut_payload_224_11 = (_zz_dataOut_payload_192_86 ? _zz_dataOut_payload_192_43 : _zz_dataOut_payload_192_11);
  assign _zz_dataOut_payload_192_88 = (_zz_dataOut_payload_192_12 < _zz_dataOut_payload_192_44);
  assign _zz_dataOut_payload_192_89 = (_zz_dataOut_payload_192_88 ? _zz_dataOut_payload_192_12 : _zz_dataOut_payload_192_44);
  assign _zz_dataOut_payload_224_12 = (_zz_dataOut_payload_192_88 ? _zz_dataOut_payload_192_44 : _zz_dataOut_payload_192_12);
  assign _zz_dataOut_payload_192_90 = (_zz_dataOut_payload_192_13 < _zz_dataOut_payload_192_45);
  assign _zz_dataOut_payload_192_91 = (_zz_dataOut_payload_192_90 ? _zz_dataOut_payload_192_13 : _zz_dataOut_payload_192_45);
  assign _zz_dataOut_payload_224_13 = (_zz_dataOut_payload_192_90 ? _zz_dataOut_payload_192_45 : _zz_dataOut_payload_192_13);
  assign _zz_dataOut_payload_192_92 = (_zz_dataOut_payload_192_14 < _zz_dataOut_payload_192_46);
  assign _zz_dataOut_payload_192_93 = (_zz_dataOut_payload_192_92 ? _zz_dataOut_payload_192_14 : _zz_dataOut_payload_192_46);
  assign _zz_dataOut_payload_224_14 = (_zz_dataOut_payload_192_92 ? _zz_dataOut_payload_192_46 : _zz_dataOut_payload_192_14);
  assign _zz_dataOut_payload_192_94 = (_zz_dataOut_payload_192_15 < _zz_dataOut_payload_192_47);
  assign _zz_dataOut_payload_192_95 = (_zz_dataOut_payload_192_94 ? _zz_dataOut_payload_192_15 : _zz_dataOut_payload_192_47);
  assign _zz_dataOut_payload_224_15 = (_zz_dataOut_payload_192_94 ? _zz_dataOut_payload_192_47 : _zz_dataOut_payload_192_15);
  assign _zz_dataOut_payload_192_96 = (_zz_dataOut_payload_192_16 < _zz_dataOut_payload_192_48);
  assign _zz_dataOut_payload_192_97 = (_zz_dataOut_payload_192_96 ? _zz_dataOut_payload_192_16 : _zz_dataOut_payload_192_48);
  assign _zz_dataOut_payload_224_16 = (_zz_dataOut_payload_192_96 ? _zz_dataOut_payload_192_48 : _zz_dataOut_payload_192_16);
  assign _zz_dataOut_payload_192_98 = (_zz_dataOut_payload_192_17 < _zz_dataOut_payload_192_49);
  assign _zz_dataOut_payload_192_99 = (_zz_dataOut_payload_192_98 ? _zz_dataOut_payload_192_17 : _zz_dataOut_payload_192_49);
  assign _zz_dataOut_payload_224_17 = (_zz_dataOut_payload_192_98 ? _zz_dataOut_payload_192_49 : _zz_dataOut_payload_192_17);
  assign _zz_dataOut_payload_192_100 = (_zz_dataOut_payload_192_18 < _zz_dataOut_payload_192_50);
  assign _zz_dataOut_payload_192_101 = (_zz_dataOut_payload_192_100 ? _zz_dataOut_payload_192_18 : _zz_dataOut_payload_192_50);
  assign _zz_dataOut_payload_224_18 = (_zz_dataOut_payload_192_100 ? _zz_dataOut_payload_192_50 : _zz_dataOut_payload_192_18);
  assign _zz_dataOut_payload_192_102 = (_zz_dataOut_payload_192_19 < _zz_dataOut_payload_192_51);
  assign _zz_dataOut_payload_192_103 = (_zz_dataOut_payload_192_102 ? _zz_dataOut_payload_192_19 : _zz_dataOut_payload_192_51);
  assign _zz_dataOut_payload_224_19 = (_zz_dataOut_payload_192_102 ? _zz_dataOut_payload_192_51 : _zz_dataOut_payload_192_19);
  assign _zz_dataOut_payload_192_104 = (_zz_dataOut_payload_192_20 < _zz_dataOut_payload_192_52);
  assign _zz_dataOut_payload_192_105 = (_zz_dataOut_payload_192_104 ? _zz_dataOut_payload_192_20 : _zz_dataOut_payload_192_52);
  assign _zz_dataOut_payload_224_20 = (_zz_dataOut_payload_192_104 ? _zz_dataOut_payload_192_52 : _zz_dataOut_payload_192_20);
  assign _zz_dataOut_payload_192_106 = (_zz_dataOut_payload_192_21 < _zz_dataOut_payload_192_53);
  assign _zz_dataOut_payload_192_107 = (_zz_dataOut_payload_192_106 ? _zz_dataOut_payload_192_21 : _zz_dataOut_payload_192_53);
  assign _zz_dataOut_payload_224_21 = (_zz_dataOut_payload_192_106 ? _zz_dataOut_payload_192_53 : _zz_dataOut_payload_192_21);
  assign _zz_dataOut_payload_192_108 = (_zz_dataOut_payload_192_22 < _zz_dataOut_payload_192_54);
  assign _zz_dataOut_payload_192_109 = (_zz_dataOut_payload_192_108 ? _zz_dataOut_payload_192_22 : _zz_dataOut_payload_192_54);
  assign _zz_dataOut_payload_224_22 = (_zz_dataOut_payload_192_108 ? _zz_dataOut_payload_192_54 : _zz_dataOut_payload_192_22);
  assign _zz_dataOut_payload_192_110 = (_zz_dataOut_payload_192_23 < _zz_dataOut_payload_192_55);
  assign _zz_dataOut_payload_192_111 = (_zz_dataOut_payload_192_110 ? _zz_dataOut_payload_192_23 : _zz_dataOut_payload_192_55);
  assign _zz_dataOut_payload_224_23 = (_zz_dataOut_payload_192_110 ? _zz_dataOut_payload_192_55 : _zz_dataOut_payload_192_23);
  assign _zz_dataOut_payload_192_112 = (_zz_dataOut_payload_192_24 < _zz_dataOut_payload_192_56);
  assign _zz_dataOut_payload_192_113 = (_zz_dataOut_payload_192_112 ? _zz_dataOut_payload_192_24 : _zz_dataOut_payload_192_56);
  assign _zz_dataOut_payload_224_24 = (_zz_dataOut_payload_192_112 ? _zz_dataOut_payload_192_56 : _zz_dataOut_payload_192_24);
  assign _zz_dataOut_payload_192_114 = (_zz_dataOut_payload_192_25 < _zz_dataOut_payload_192_57);
  assign _zz_dataOut_payload_192_115 = (_zz_dataOut_payload_192_114 ? _zz_dataOut_payload_192_25 : _zz_dataOut_payload_192_57);
  assign _zz_dataOut_payload_224_25 = (_zz_dataOut_payload_192_114 ? _zz_dataOut_payload_192_57 : _zz_dataOut_payload_192_25);
  assign _zz_dataOut_payload_192_116 = (_zz_dataOut_payload_192_26 < _zz_dataOut_payload_192_58);
  assign _zz_dataOut_payload_192_117 = (_zz_dataOut_payload_192_116 ? _zz_dataOut_payload_192_26 : _zz_dataOut_payload_192_58);
  assign _zz_dataOut_payload_224_26 = (_zz_dataOut_payload_192_116 ? _zz_dataOut_payload_192_58 : _zz_dataOut_payload_192_26);
  assign _zz_dataOut_payload_192_118 = (_zz_dataOut_payload_192_27 < _zz_dataOut_payload_192_59);
  assign _zz_dataOut_payload_192_119 = (_zz_dataOut_payload_192_118 ? _zz_dataOut_payload_192_27 : _zz_dataOut_payload_192_59);
  assign _zz_dataOut_payload_224_27 = (_zz_dataOut_payload_192_118 ? _zz_dataOut_payload_192_59 : _zz_dataOut_payload_192_27);
  assign _zz_dataOut_payload_192_120 = (_zz_dataOut_payload_192_28 < _zz_dataOut_payload_192_60);
  assign _zz_dataOut_payload_192_121 = (_zz_dataOut_payload_192_120 ? _zz_dataOut_payload_192_28 : _zz_dataOut_payload_192_60);
  assign _zz_dataOut_payload_224_28 = (_zz_dataOut_payload_192_120 ? _zz_dataOut_payload_192_60 : _zz_dataOut_payload_192_28);
  assign _zz_dataOut_payload_192_122 = (_zz_dataOut_payload_192_29 < _zz_dataOut_payload_192_61);
  assign _zz_dataOut_payload_192_123 = (_zz_dataOut_payload_192_122 ? _zz_dataOut_payload_192_29 : _zz_dataOut_payload_192_61);
  assign _zz_dataOut_payload_224_29 = (_zz_dataOut_payload_192_122 ? _zz_dataOut_payload_192_61 : _zz_dataOut_payload_192_29);
  assign _zz_dataOut_payload_192_124 = (_zz_dataOut_payload_192_30 < _zz_dataOut_payload_192_62);
  assign _zz_dataOut_payload_192_125 = (_zz_dataOut_payload_192_124 ? _zz_dataOut_payload_192_30 : _zz_dataOut_payload_192_62);
  assign _zz_dataOut_payload_224_30 = (_zz_dataOut_payload_192_124 ? _zz_dataOut_payload_192_62 : _zz_dataOut_payload_192_30);
  assign _zz_dataOut_payload_192_126 = (_zz_dataOut_payload_192_31 < _zz_dataOut_payload_192_63);
  assign _zz_dataOut_payload_192_127 = (_zz_dataOut_payload_192_126 ? _zz_dataOut_payload_192_31 : _zz_dataOut_payload_192_63);
  assign _zz_dataOut_payload_224_31 = (_zz_dataOut_payload_192_126 ? _zz_dataOut_payload_192_63 : _zz_dataOut_payload_192_31);
  assign _zz_dataOut_payload_192_128 = (_zz_dataOut_payload_192_65 < _zz_dataOut_payload_192_97);
  assign _zz_dataOut_payload_192_129 = (_zz_dataOut_payload_192_128 ? _zz_dataOut_payload_192_65 : _zz_dataOut_payload_192_97);
  assign _zz_dataOut_payload_208 = (_zz_dataOut_payload_192_128 ? _zz_dataOut_payload_192_97 : _zz_dataOut_payload_192_65);
  assign _zz_dataOut_payload_192_130 = (_zz_dataOut_payload_192_67 < _zz_dataOut_payload_192_99);
  assign _zz_dataOut_payload_192_131 = (_zz_dataOut_payload_192_130 ? _zz_dataOut_payload_192_67 : _zz_dataOut_payload_192_99);
  assign _zz_dataOut_payload_208_1 = (_zz_dataOut_payload_192_130 ? _zz_dataOut_payload_192_99 : _zz_dataOut_payload_192_67);
  assign _zz_dataOut_payload_192_132 = (_zz_dataOut_payload_192_69 < _zz_dataOut_payload_192_101);
  assign _zz_dataOut_payload_192_133 = (_zz_dataOut_payload_192_132 ? _zz_dataOut_payload_192_69 : _zz_dataOut_payload_192_101);
  assign _zz_dataOut_payload_208_2 = (_zz_dataOut_payload_192_132 ? _zz_dataOut_payload_192_101 : _zz_dataOut_payload_192_69);
  assign _zz_dataOut_payload_192_134 = (_zz_dataOut_payload_192_71 < _zz_dataOut_payload_192_103);
  assign _zz_dataOut_payload_192_135 = (_zz_dataOut_payload_192_134 ? _zz_dataOut_payload_192_71 : _zz_dataOut_payload_192_103);
  assign _zz_dataOut_payload_208_3 = (_zz_dataOut_payload_192_134 ? _zz_dataOut_payload_192_103 : _zz_dataOut_payload_192_71);
  assign _zz_dataOut_payload_192_136 = (_zz_dataOut_payload_192_73 < _zz_dataOut_payload_192_105);
  assign _zz_dataOut_payload_192_137 = (_zz_dataOut_payload_192_136 ? _zz_dataOut_payload_192_73 : _zz_dataOut_payload_192_105);
  assign _zz_dataOut_payload_208_4 = (_zz_dataOut_payload_192_136 ? _zz_dataOut_payload_192_105 : _zz_dataOut_payload_192_73);
  assign _zz_dataOut_payload_192_138 = (_zz_dataOut_payload_192_75 < _zz_dataOut_payload_192_107);
  assign _zz_dataOut_payload_192_139 = (_zz_dataOut_payload_192_138 ? _zz_dataOut_payload_192_75 : _zz_dataOut_payload_192_107);
  assign _zz_dataOut_payload_208_5 = (_zz_dataOut_payload_192_138 ? _zz_dataOut_payload_192_107 : _zz_dataOut_payload_192_75);
  assign _zz_dataOut_payload_192_140 = (_zz_dataOut_payload_192_77 < _zz_dataOut_payload_192_109);
  assign _zz_dataOut_payload_192_141 = (_zz_dataOut_payload_192_140 ? _zz_dataOut_payload_192_77 : _zz_dataOut_payload_192_109);
  assign _zz_dataOut_payload_208_6 = (_zz_dataOut_payload_192_140 ? _zz_dataOut_payload_192_109 : _zz_dataOut_payload_192_77);
  assign _zz_dataOut_payload_192_142 = (_zz_dataOut_payload_192_79 < _zz_dataOut_payload_192_111);
  assign _zz_dataOut_payload_192_143 = (_zz_dataOut_payload_192_142 ? _zz_dataOut_payload_192_79 : _zz_dataOut_payload_192_111);
  assign _zz_dataOut_payload_208_7 = (_zz_dataOut_payload_192_142 ? _zz_dataOut_payload_192_111 : _zz_dataOut_payload_192_79);
  assign _zz_dataOut_payload_192_144 = (_zz_dataOut_payload_192_81 < _zz_dataOut_payload_192_113);
  assign _zz_dataOut_payload_192_145 = (_zz_dataOut_payload_192_144 ? _zz_dataOut_payload_192_81 : _zz_dataOut_payload_192_113);
  assign _zz_dataOut_payload_208_8 = (_zz_dataOut_payload_192_144 ? _zz_dataOut_payload_192_113 : _zz_dataOut_payload_192_81);
  assign _zz_dataOut_payload_192_146 = (_zz_dataOut_payload_192_83 < _zz_dataOut_payload_192_115);
  assign _zz_dataOut_payload_192_147 = (_zz_dataOut_payload_192_146 ? _zz_dataOut_payload_192_83 : _zz_dataOut_payload_192_115);
  assign _zz_dataOut_payload_208_9 = (_zz_dataOut_payload_192_146 ? _zz_dataOut_payload_192_115 : _zz_dataOut_payload_192_83);
  assign _zz_dataOut_payload_192_148 = (_zz_dataOut_payload_192_85 < _zz_dataOut_payload_192_117);
  assign _zz_dataOut_payload_192_149 = (_zz_dataOut_payload_192_148 ? _zz_dataOut_payload_192_85 : _zz_dataOut_payload_192_117);
  assign _zz_dataOut_payload_208_10 = (_zz_dataOut_payload_192_148 ? _zz_dataOut_payload_192_117 : _zz_dataOut_payload_192_85);
  assign _zz_dataOut_payload_192_150 = (_zz_dataOut_payload_192_87 < _zz_dataOut_payload_192_119);
  assign _zz_dataOut_payload_192_151 = (_zz_dataOut_payload_192_150 ? _zz_dataOut_payload_192_87 : _zz_dataOut_payload_192_119);
  assign _zz_dataOut_payload_208_11 = (_zz_dataOut_payload_192_150 ? _zz_dataOut_payload_192_119 : _zz_dataOut_payload_192_87);
  assign _zz_dataOut_payload_192_152 = (_zz_dataOut_payload_192_89 < _zz_dataOut_payload_192_121);
  assign _zz_dataOut_payload_192_153 = (_zz_dataOut_payload_192_152 ? _zz_dataOut_payload_192_89 : _zz_dataOut_payload_192_121);
  assign _zz_dataOut_payload_208_12 = (_zz_dataOut_payload_192_152 ? _zz_dataOut_payload_192_121 : _zz_dataOut_payload_192_89);
  assign _zz_dataOut_payload_192_154 = (_zz_dataOut_payload_192_91 < _zz_dataOut_payload_192_123);
  assign _zz_dataOut_payload_192_155 = (_zz_dataOut_payload_192_154 ? _zz_dataOut_payload_192_91 : _zz_dataOut_payload_192_123);
  assign _zz_dataOut_payload_208_13 = (_zz_dataOut_payload_192_154 ? _zz_dataOut_payload_192_123 : _zz_dataOut_payload_192_91);
  assign _zz_dataOut_payload_192_156 = (_zz_dataOut_payload_192_93 < _zz_dataOut_payload_192_125);
  assign _zz_dataOut_payload_192_157 = (_zz_dataOut_payload_192_156 ? _zz_dataOut_payload_192_93 : _zz_dataOut_payload_192_125);
  assign _zz_dataOut_payload_208_14 = (_zz_dataOut_payload_192_156 ? _zz_dataOut_payload_192_125 : _zz_dataOut_payload_192_93);
  assign _zz_dataOut_payload_192_158 = (_zz_dataOut_payload_192_95 < _zz_dataOut_payload_192_127);
  assign _zz_dataOut_payload_192_159 = (_zz_dataOut_payload_192_158 ? _zz_dataOut_payload_192_95 : _zz_dataOut_payload_192_127);
  assign _zz_dataOut_payload_208_15 = (_zz_dataOut_payload_192_158 ? _zz_dataOut_payload_192_127 : _zz_dataOut_payload_192_95);
  assign _zz_dataOut_payload_192_160 = (_zz_dataOut_payload_192_129 < _zz_dataOut_payload_192_145);
  assign _zz_dataOut_payload_192_161 = (_zz_dataOut_payload_192_160 ? _zz_dataOut_payload_192_129 : _zz_dataOut_payload_192_145);
  assign _zz_dataOut_payload_200 = (_zz_dataOut_payload_192_160 ? _zz_dataOut_payload_192_145 : _zz_dataOut_payload_192_129);
  assign _zz_dataOut_payload_192_162 = (_zz_dataOut_payload_192_131 < _zz_dataOut_payload_192_147);
  assign _zz_dataOut_payload_192_163 = (_zz_dataOut_payload_192_162 ? _zz_dataOut_payload_192_131 : _zz_dataOut_payload_192_147);
  assign _zz_dataOut_payload_200_1 = (_zz_dataOut_payload_192_162 ? _zz_dataOut_payload_192_147 : _zz_dataOut_payload_192_131);
  assign _zz_dataOut_payload_192_164 = (_zz_dataOut_payload_192_133 < _zz_dataOut_payload_192_149);
  assign _zz_dataOut_payload_192_165 = (_zz_dataOut_payload_192_164 ? _zz_dataOut_payload_192_133 : _zz_dataOut_payload_192_149);
  assign _zz_dataOut_payload_200_2 = (_zz_dataOut_payload_192_164 ? _zz_dataOut_payload_192_149 : _zz_dataOut_payload_192_133);
  assign _zz_dataOut_payload_192_166 = (_zz_dataOut_payload_192_135 < _zz_dataOut_payload_192_151);
  assign _zz_dataOut_payload_192_167 = (_zz_dataOut_payload_192_166 ? _zz_dataOut_payload_192_135 : _zz_dataOut_payload_192_151);
  assign _zz_dataOut_payload_200_3 = (_zz_dataOut_payload_192_166 ? _zz_dataOut_payload_192_151 : _zz_dataOut_payload_192_135);
  assign _zz_dataOut_payload_192_168 = (_zz_dataOut_payload_192_137 < _zz_dataOut_payload_192_153);
  assign _zz_dataOut_payload_192_169 = (_zz_dataOut_payload_192_168 ? _zz_dataOut_payload_192_137 : _zz_dataOut_payload_192_153);
  assign _zz_dataOut_payload_200_4 = (_zz_dataOut_payload_192_168 ? _zz_dataOut_payload_192_153 : _zz_dataOut_payload_192_137);
  assign _zz_dataOut_payload_192_170 = (_zz_dataOut_payload_192_139 < _zz_dataOut_payload_192_155);
  assign _zz_dataOut_payload_192_171 = (_zz_dataOut_payload_192_170 ? _zz_dataOut_payload_192_139 : _zz_dataOut_payload_192_155);
  assign _zz_dataOut_payload_200_5 = (_zz_dataOut_payload_192_170 ? _zz_dataOut_payload_192_155 : _zz_dataOut_payload_192_139);
  assign _zz_dataOut_payload_192_172 = (_zz_dataOut_payload_192_141 < _zz_dataOut_payload_192_157);
  assign _zz_dataOut_payload_192_173 = (_zz_dataOut_payload_192_172 ? _zz_dataOut_payload_192_141 : _zz_dataOut_payload_192_157);
  assign _zz_dataOut_payload_200_6 = (_zz_dataOut_payload_192_172 ? _zz_dataOut_payload_192_157 : _zz_dataOut_payload_192_141);
  assign _zz_dataOut_payload_192_174 = (_zz_dataOut_payload_192_143 < _zz_dataOut_payload_192_159);
  assign _zz_dataOut_payload_192_175 = (_zz_dataOut_payload_192_174 ? _zz_dataOut_payload_192_143 : _zz_dataOut_payload_192_159);
  assign _zz_dataOut_payload_200_7 = (_zz_dataOut_payload_192_174 ? _zz_dataOut_payload_192_159 : _zz_dataOut_payload_192_143);
  assign _zz_dataOut_payload_192_176 = (_zz_dataOut_payload_192_161 < _zz_dataOut_payload_192_169);
  assign _zz_dataOut_payload_192_177 = (_zz_dataOut_payload_192_176 ? _zz_dataOut_payload_192_161 : _zz_dataOut_payload_192_169);
  assign _zz_dataOut_payload_196 = (_zz_dataOut_payload_192_176 ? _zz_dataOut_payload_192_169 : _zz_dataOut_payload_192_161);
  assign _zz_dataOut_payload_192_178 = (_zz_dataOut_payload_192_163 < _zz_dataOut_payload_192_171);
  assign _zz_dataOut_payload_192_179 = (_zz_dataOut_payload_192_178 ? _zz_dataOut_payload_192_163 : _zz_dataOut_payload_192_171);
  assign _zz_dataOut_payload_196_1 = (_zz_dataOut_payload_192_178 ? _zz_dataOut_payload_192_171 : _zz_dataOut_payload_192_163);
  assign _zz_dataOut_payload_192_180 = (_zz_dataOut_payload_192_165 < _zz_dataOut_payload_192_173);
  assign _zz_dataOut_payload_192_181 = (_zz_dataOut_payload_192_180 ? _zz_dataOut_payload_192_165 : _zz_dataOut_payload_192_173);
  assign _zz_dataOut_payload_196_2 = (_zz_dataOut_payload_192_180 ? _zz_dataOut_payload_192_173 : _zz_dataOut_payload_192_165);
  assign _zz_dataOut_payload_192_182 = (_zz_dataOut_payload_192_167 < _zz_dataOut_payload_192_175);
  assign _zz_dataOut_payload_192_183 = (_zz_dataOut_payload_192_182 ? _zz_dataOut_payload_192_167 : _zz_dataOut_payload_192_175);
  assign _zz_dataOut_payload_196_3 = (_zz_dataOut_payload_192_182 ? _zz_dataOut_payload_192_175 : _zz_dataOut_payload_192_167);
  assign _zz_dataOut_payload_192_184 = (_zz_dataOut_payload_192_177 < _zz_dataOut_payload_192_181);
  assign _zz_dataOut_payload_192_185 = (_zz_dataOut_payload_192_184 ? _zz_dataOut_payload_192_177 : _zz_dataOut_payload_192_181);
  assign _zz_dataOut_payload_194 = (_zz_dataOut_payload_192_184 ? _zz_dataOut_payload_192_181 : _zz_dataOut_payload_192_177);
  assign _zz_dataOut_payload_192_186 = (_zz_dataOut_payload_192_179 < _zz_dataOut_payload_192_183);
  assign _zz_dataOut_payload_192_187 = (_zz_dataOut_payload_192_186 ? _zz_dataOut_payload_192_179 : _zz_dataOut_payload_192_183);
  assign _zz_dataOut_payload_194_1 = (_zz_dataOut_payload_192_186 ? _zz_dataOut_payload_192_183 : _zz_dataOut_payload_192_179);
  assign _zz_dataOut_payload_192_188 = (_zz_dataOut_payload_192_185 < _zz_dataOut_payload_192_187);
  assign _zz_dataOut_payload_194_2 = (_zz_dataOut_payload_194 < _zz_dataOut_payload_194_1);
  assign _zz_dataOut_payload_196_4 = (_zz_dataOut_payload_196 < _zz_dataOut_payload_196_2);
  assign _zz_dataOut_payload_196_5 = (_zz_dataOut_payload_196_4 ? _zz_dataOut_payload_196 : _zz_dataOut_payload_196_2);
  assign _zz_dataOut_payload_198 = (_zz_dataOut_payload_196_4 ? _zz_dataOut_payload_196_2 : _zz_dataOut_payload_196);
  assign _zz_dataOut_payload_196_6 = (_zz_dataOut_payload_196_1 < _zz_dataOut_payload_196_3);
  assign _zz_dataOut_payload_196_7 = (_zz_dataOut_payload_196_6 ? _zz_dataOut_payload_196_1 : _zz_dataOut_payload_196_3);
  assign _zz_dataOut_payload_198_1 = (_zz_dataOut_payload_196_6 ? _zz_dataOut_payload_196_3 : _zz_dataOut_payload_196_1);
  assign _zz_dataOut_payload_196_8 = (_zz_dataOut_payload_196_5 < _zz_dataOut_payload_196_7);
  assign _zz_dataOut_payload_198_2 = (_zz_dataOut_payload_198 < _zz_dataOut_payload_198_1);
  assign _zz_dataOut_payload_200_8 = (_zz_dataOut_payload_200 < _zz_dataOut_payload_200_4);
  assign _zz_dataOut_payload_200_9 = (_zz_dataOut_payload_200_8 ? _zz_dataOut_payload_200 : _zz_dataOut_payload_200_4);
  assign _zz_dataOut_payload_204 = (_zz_dataOut_payload_200_8 ? _zz_dataOut_payload_200_4 : _zz_dataOut_payload_200);
  assign _zz_dataOut_payload_200_10 = (_zz_dataOut_payload_200_1 < _zz_dataOut_payload_200_5);
  assign _zz_dataOut_payload_200_11 = (_zz_dataOut_payload_200_10 ? _zz_dataOut_payload_200_1 : _zz_dataOut_payload_200_5);
  assign _zz_dataOut_payload_204_1 = (_zz_dataOut_payload_200_10 ? _zz_dataOut_payload_200_5 : _zz_dataOut_payload_200_1);
  assign _zz_dataOut_payload_200_12 = (_zz_dataOut_payload_200_2 < _zz_dataOut_payload_200_6);
  assign _zz_dataOut_payload_200_13 = (_zz_dataOut_payload_200_12 ? _zz_dataOut_payload_200_2 : _zz_dataOut_payload_200_6);
  assign _zz_dataOut_payload_204_2 = (_zz_dataOut_payload_200_12 ? _zz_dataOut_payload_200_6 : _zz_dataOut_payload_200_2);
  assign _zz_dataOut_payload_200_14 = (_zz_dataOut_payload_200_3 < _zz_dataOut_payload_200_7);
  assign _zz_dataOut_payload_200_15 = (_zz_dataOut_payload_200_14 ? _zz_dataOut_payload_200_3 : _zz_dataOut_payload_200_7);
  assign _zz_dataOut_payload_204_3 = (_zz_dataOut_payload_200_14 ? _zz_dataOut_payload_200_7 : _zz_dataOut_payload_200_3);
  assign _zz_dataOut_payload_200_16 = (_zz_dataOut_payload_200_9 < _zz_dataOut_payload_200_13);
  assign _zz_dataOut_payload_200_17 = (_zz_dataOut_payload_200_16 ? _zz_dataOut_payload_200_9 : _zz_dataOut_payload_200_13);
  assign _zz_dataOut_payload_202 = (_zz_dataOut_payload_200_16 ? _zz_dataOut_payload_200_13 : _zz_dataOut_payload_200_9);
  assign _zz_dataOut_payload_200_18 = (_zz_dataOut_payload_200_11 < _zz_dataOut_payload_200_15);
  assign _zz_dataOut_payload_200_19 = (_zz_dataOut_payload_200_18 ? _zz_dataOut_payload_200_11 : _zz_dataOut_payload_200_15);
  assign _zz_dataOut_payload_202_1 = (_zz_dataOut_payload_200_18 ? _zz_dataOut_payload_200_15 : _zz_dataOut_payload_200_11);
  assign _zz_dataOut_payload_200_20 = (_zz_dataOut_payload_200_17 < _zz_dataOut_payload_200_19);
  assign _zz_dataOut_payload_202_2 = (_zz_dataOut_payload_202 < _zz_dataOut_payload_202_1);
  assign _zz_dataOut_payload_204_4 = (_zz_dataOut_payload_204 < _zz_dataOut_payload_204_2);
  assign _zz_dataOut_payload_204_5 = (_zz_dataOut_payload_204_4 ? _zz_dataOut_payload_204 : _zz_dataOut_payload_204_2);
  assign _zz_dataOut_payload_206 = (_zz_dataOut_payload_204_4 ? _zz_dataOut_payload_204_2 : _zz_dataOut_payload_204);
  assign _zz_dataOut_payload_204_6 = (_zz_dataOut_payload_204_1 < _zz_dataOut_payload_204_3);
  assign _zz_dataOut_payload_204_7 = (_zz_dataOut_payload_204_6 ? _zz_dataOut_payload_204_1 : _zz_dataOut_payload_204_3);
  assign _zz_dataOut_payload_206_1 = (_zz_dataOut_payload_204_6 ? _zz_dataOut_payload_204_3 : _zz_dataOut_payload_204_1);
  assign _zz_dataOut_payload_204_8 = (_zz_dataOut_payload_204_5 < _zz_dataOut_payload_204_7);
  assign _zz_dataOut_payload_206_2 = (_zz_dataOut_payload_206 < _zz_dataOut_payload_206_1);
  assign _zz_dataOut_payload_208_16 = (_zz_dataOut_payload_208 < _zz_dataOut_payload_208_8);
  assign _zz_dataOut_payload_208_17 = (_zz_dataOut_payload_208_16 ? _zz_dataOut_payload_208 : _zz_dataOut_payload_208_8);
  assign _zz_dataOut_payload_216 = (_zz_dataOut_payload_208_16 ? _zz_dataOut_payload_208_8 : _zz_dataOut_payload_208);
  assign _zz_dataOut_payload_208_18 = (_zz_dataOut_payload_208_1 < _zz_dataOut_payload_208_9);
  assign _zz_dataOut_payload_208_19 = (_zz_dataOut_payload_208_18 ? _zz_dataOut_payload_208_1 : _zz_dataOut_payload_208_9);
  assign _zz_dataOut_payload_216_1 = (_zz_dataOut_payload_208_18 ? _zz_dataOut_payload_208_9 : _zz_dataOut_payload_208_1);
  assign _zz_dataOut_payload_208_20 = (_zz_dataOut_payload_208_2 < _zz_dataOut_payload_208_10);
  assign _zz_dataOut_payload_208_21 = (_zz_dataOut_payload_208_20 ? _zz_dataOut_payload_208_2 : _zz_dataOut_payload_208_10);
  assign _zz_dataOut_payload_216_2 = (_zz_dataOut_payload_208_20 ? _zz_dataOut_payload_208_10 : _zz_dataOut_payload_208_2);
  assign _zz_dataOut_payload_208_22 = (_zz_dataOut_payload_208_3 < _zz_dataOut_payload_208_11);
  assign _zz_dataOut_payload_208_23 = (_zz_dataOut_payload_208_22 ? _zz_dataOut_payload_208_3 : _zz_dataOut_payload_208_11);
  assign _zz_dataOut_payload_216_3 = (_zz_dataOut_payload_208_22 ? _zz_dataOut_payload_208_11 : _zz_dataOut_payload_208_3);
  assign _zz_dataOut_payload_208_24 = (_zz_dataOut_payload_208_4 < _zz_dataOut_payload_208_12);
  assign _zz_dataOut_payload_208_25 = (_zz_dataOut_payload_208_24 ? _zz_dataOut_payload_208_4 : _zz_dataOut_payload_208_12);
  assign _zz_dataOut_payload_216_4 = (_zz_dataOut_payload_208_24 ? _zz_dataOut_payload_208_12 : _zz_dataOut_payload_208_4);
  assign _zz_dataOut_payload_208_26 = (_zz_dataOut_payload_208_5 < _zz_dataOut_payload_208_13);
  assign _zz_dataOut_payload_208_27 = (_zz_dataOut_payload_208_26 ? _zz_dataOut_payload_208_5 : _zz_dataOut_payload_208_13);
  assign _zz_dataOut_payload_216_5 = (_zz_dataOut_payload_208_26 ? _zz_dataOut_payload_208_13 : _zz_dataOut_payload_208_5);
  assign _zz_dataOut_payload_208_28 = (_zz_dataOut_payload_208_6 < _zz_dataOut_payload_208_14);
  assign _zz_dataOut_payload_208_29 = (_zz_dataOut_payload_208_28 ? _zz_dataOut_payload_208_6 : _zz_dataOut_payload_208_14);
  assign _zz_dataOut_payload_216_6 = (_zz_dataOut_payload_208_28 ? _zz_dataOut_payload_208_14 : _zz_dataOut_payload_208_6);
  assign _zz_dataOut_payload_208_30 = (_zz_dataOut_payload_208_7 < _zz_dataOut_payload_208_15);
  assign _zz_dataOut_payload_208_31 = (_zz_dataOut_payload_208_30 ? _zz_dataOut_payload_208_7 : _zz_dataOut_payload_208_15);
  assign _zz_dataOut_payload_216_7 = (_zz_dataOut_payload_208_30 ? _zz_dataOut_payload_208_15 : _zz_dataOut_payload_208_7);
  assign _zz_dataOut_payload_208_32 = (_zz_dataOut_payload_208_17 < _zz_dataOut_payload_208_25);
  assign _zz_dataOut_payload_208_33 = (_zz_dataOut_payload_208_32 ? _zz_dataOut_payload_208_17 : _zz_dataOut_payload_208_25);
  assign _zz_dataOut_payload_212 = (_zz_dataOut_payload_208_32 ? _zz_dataOut_payload_208_25 : _zz_dataOut_payload_208_17);
  assign _zz_dataOut_payload_208_34 = (_zz_dataOut_payload_208_19 < _zz_dataOut_payload_208_27);
  assign _zz_dataOut_payload_208_35 = (_zz_dataOut_payload_208_34 ? _zz_dataOut_payload_208_19 : _zz_dataOut_payload_208_27);
  assign _zz_dataOut_payload_212_1 = (_zz_dataOut_payload_208_34 ? _zz_dataOut_payload_208_27 : _zz_dataOut_payload_208_19);
  assign _zz_dataOut_payload_208_36 = (_zz_dataOut_payload_208_21 < _zz_dataOut_payload_208_29);
  assign _zz_dataOut_payload_208_37 = (_zz_dataOut_payload_208_36 ? _zz_dataOut_payload_208_21 : _zz_dataOut_payload_208_29);
  assign _zz_dataOut_payload_212_2 = (_zz_dataOut_payload_208_36 ? _zz_dataOut_payload_208_29 : _zz_dataOut_payload_208_21);
  assign _zz_dataOut_payload_208_38 = (_zz_dataOut_payload_208_23 < _zz_dataOut_payload_208_31);
  assign _zz_dataOut_payload_208_39 = (_zz_dataOut_payload_208_38 ? _zz_dataOut_payload_208_23 : _zz_dataOut_payload_208_31);
  assign _zz_dataOut_payload_212_3 = (_zz_dataOut_payload_208_38 ? _zz_dataOut_payload_208_31 : _zz_dataOut_payload_208_23);
  assign _zz_dataOut_payload_208_40 = (_zz_dataOut_payload_208_33 < _zz_dataOut_payload_208_37);
  assign _zz_dataOut_payload_208_41 = (_zz_dataOut_payload_208_40 ? _zz_dataOut_payload_208_33 : _zz_dataOut_payload_208_37);
  assign _zz_dataOut_payload_210 = (_zz_dataOut_payload_208_40 ? _zz_dataOut_payload_208_37 : _zz_dataOut_payload_208_33);
  assign _zz_dataOut_payload_208_42 = (_zz_dataOut_payload_208_35 < _zz_dataOut_payload_208_39);
  assign _zz_dataOut_payload_208_43 = (_zz_dataOut_payload_208_42 ? _zz_dataOut_payload_208_35 : _zz_dataOut_payload_208_39);
  assign _zz_dataOut_payload_210_1 = (_zz_dataOut_payload_208_42 ? _zz_dataOut_payload_208_39 : _zz_dataOut_payload_208_35);
  assign _zz_dataOut_payload_208_44 = (_zz_dataOut_payload_208_41 < _zz_dataOut_payload_208_43);
  assign _zz_dataOut_payload_210_2 = (_zz_dataOut_payload_210 < _zz_dataOut_payload_210_1);
  assign _zz_dataOut_payload_212_4 = (_zz_dataOut_payload_212 < _zz_dataOut_payload_212_2);
  assign _zz_dataOut_payload_212_5 = (_zz_dataOut_payload_212_4 ? _zz_dataOut_payload_212 : _zz_dataOut_payload_212_2);
  assign _zz_dataOut_payload_214 = (_zz_dataOut_payload_212_4 ? _zz_dataOut_payload_212_2 : _zz_dataOut_payload_212);
  assign _zz_dataOut_payload_212_6 = (_zz_dataOut_payload_212_1 < _zz_dataOut_payload_212_3);
  assign _zz_dataOut_payload_212_7 = (_zz_dataOut_payload_212_6 ? _zz_dataOut_payload_212_1 : _zz_dataOut_payload_212_3);
  assign _zz_dataOut_payload_214_1 = (_zz_dataOut_payload_212_6 ? _zz_dataOut_payload_212_3 : _zz_dataOut_payload_212_1);
  assign _zz_dataOut_payload_212_8 = (_zz_dataOut_payload_212_5 < _zz_dataOut_payload_212_7);
  assign _zz_dataOut_payload_214_2 = (_zz_dataOut_payload_214 < _zz_dataOut_payload_214_1);
  assign _zz_dataOut_payload_216_8 = (_zz_dataOut_payload_216 < _zz_dataOut_payload_216_4);
  assign _zz_dataOut_payload_216_9 = (_zz_dataOut_payload_216_8 ? _zz_dataOut_payload_216 : _zz_dataOut_payload_216_4);
  assign _zz_dataOut_payload_220 = (_zz_dataOut_payload_216_8 ? _zz_dataOut_payload_216_4 : _zz_dataOut_payload_216);
  assign _zz_dataOut_payload_216_10 = (_zz_dataOut_payload_216_1 < _zz_dataOut_payload_216_5);
  assign _zz_dataOut_payload_216_11 = (_zz_dataOut_payload_216_10 ? _zz_dataOut_payload_216_1 : _zz_dataOut_payload_216_5);
  assign _zz_dataOut_payload_220_1 = (_zz_dataOut_payload_216_10 ? _zz_dataOut_payload_216_5 : _zz_dataOut_payload_216_1);
  assign _zz_dataOut_payload_216_12 = (_zz_dataOut_payload_216_2 < _zz_dataOut_payload_216_6);
  assign _zz_dataOut_payload_216_13 = (_zz_dataOut_payload_216_12 ? _zz_dataOut_payload_216_2 : _zz_dataOut_payload_216_6);
  assign _zz_dataOut_payload_220_2 = (_zz_dataOut_payload_216_12 ? _zz_dataOut_payload_216_6 : _zz_dataOut_payload_216_2);
  assign _zz_dataOut_payload_216_14 = (_zz_dataOut_payload_216_3 < _zz_dataOut_payload_216_7);
  assign _zz_dataOut_payload_216_15 = (_zz_dataOut_payload_216_14 ? _zz_dataOut_payload_216_3 : _zz_dataOut_payload_216_7);
  assign _zz_dataOut_payload_220_3 = (_zz_dataOut_payload_216_14 ? _zz_dataOut_payload_216_7 : _zz_dataOut_payload_216_3);
  assign _zz_dataOut_payload_216_16 = (_zz_dataOut_payload_216_9 < _zz_dataOut_payload_216_13);
  assign _zz_dataOut_payload_216_17 = (_zz_dataOut_payload_216_16 ? _zz_dataOut_payload_216_9 : _zz_dataOut_payload_216_13);
  assign _zz_dataOut_payload_218 = (_zz_dataOut_payload_216_16 ? _zz_dataOut_payload_216_13 : _zz_dataOut_payload_216_9);
  assign _zz_dataOut_payload_216_18 = (_zz_dataOut_payload_216_11 < _zz_dataOut_payload_216_15);
  assign _zz_dataOut_payload_216_19 = (_zz_dataOut_payload_216_18 ? _zz_dataOut_payload_216_11 : _zz_dataOut_payload_216_15);
  assign _zz_dataOut_payload_218_1 = (_zz_dataOut_payload_216_18 ? _zz_dataOut_payload_216_15 : _zz_dataOut_payload_216_11);
  assign _zz_dataOut_payload_216_20 = (_zz_dataOut_payload_216_17 < _zz_dataOut_payload_216_19);
  assign _zz_dataOut_payload_218_2 = (_zz_dataOut_payload_218 < _zz_dataOut_payload_218_1);
  assign _zz_dataOut_payload_220_4 = (_zz_dataOut_payload_220 < _zz_dataOut_payload_220_2);
  assign _zz_dataOut_payload_220_5 = (_zz_dataOut_payload_220_4 ? _zz_dataOut_payload_220 : _zz_dataOut_payload_220_2);
  assign _zz_dataOut_payload_222 = (_zz_dataOut_payload_220_4 ? _zz_dataOut_payload_220_2 : _zz_dataOut_payload_220);
  assign _zz_dataOut_payload_220_6 = (_zz_dataOut_payload_220_1 < _zz_dataOut_payload_220_3);
  assign _zz_dataOut_payload_220_7 = (_zz_dataOut_payload_220_6 ? _zz_dataOut_payload_220_1 : _zz_dataOut_payload_220_3);
  assign _zz_dataOut_payload_222_1 = (_zz_dataOut_payload_220_6 ? _zz_dataOut_payload_220_3 : _zz_dataOut_payload_220_1);
  assign _zz_dataOut_payload_220_8 = (_zz_dataOut_payload_220_5 < _zz_dataOut_payload_220_7);
  assign _zz_dataOut_payload_222_2 = (_zz_dataOut_payload_222 < _zz_dataOut_payload_222_1);
  assign _zz_dataOut_payload_224_32 = (_zz_dataOut_payload_224 < _zz_dataOut_payload_224_16);
  assign _zz_dataOut_payload_224_33 = (_zz_dataOut_payload_224_32 ? _zz_dataOut_payload_224 : _zz_dataOut_payload_224_16);
  assign _zz_dataOut_payload_240 = (_zz_dataOut_payload_224_32 ? _zz_dataOut_payload_224_16 : _zz_dataOut_payload_224);
  assign _zz_dataOut_payload_224_34 = (_zz_dataOut_payload_224_1 < _zz_dataOut_payload_224_17);
  assign _zz_dataOut_payload_224_35 = (_zz_dataOut_payload_224_34 ? _zz_dataOut_payload_224_1 : _zz_dataOut_payload_224_17);
  assign _zz_dataOut_payload_240_1 = (_zz_dataOut_payload_224_34 ? _zz_dataOut_payload_224_17 : _zz_dataOut_payload_224_1);
  assign _zz_dataOut_payload_224_36 = (_zz_dataOut_payload_224_2 < _zz_dataOut_payload_224_18);
  assign _zz_dataOut_payload_224_37 = (_zz_dataOut_payload_224_36 ? _zz_dataOut_payload_224_2 : _zz_dataOut_payload_224_18);
  assign _zz_dataOut_payload_240_2 = (_zz_dataOut_payload_224_36 ? _zz_dataOut_payload_224_18 : _zz_dataOut_payload_224_2);
  assign _zz_dataOut_payload_224_38 = (_zz_dataOut_payload_224_3 < _zz_dataOut_payload_224_19);
  assign _zz_dataOut_payload_224_39 = (_zz_dataOut_payload_224_38 ? _zz_dataOut_payload_224_3 : _zz_dataOut_payload_224_19);
  assign _zz_dataOut_payload_240_3 = (_zz_dataOut_payload_224_38 ? _zz_dataOut_payload_224_19 : _zz_dataOut_payload_224_3);
  assign _zz_dataOut_payload_224_40 = (_zz_dataOut_payload_224_4 < _zz_dataOut_payload_224_20);
  assign _zz_dataOut_payload_224_41 = (_zz_dataOut_payload_224_40 ? _zz_dataOut_payload_224_4 : _zz_dataOut_payload_224_20);
  assign _zz_dataOut_payload_240_4 = (_zz_dataOut_payload_224_40 ? _zz_dataOut_payload_224_20 : _zz_dataOut_payload_224_4);
  assign _zz_dataOut_payload_224_42 = (_zz_dataOut_payload_224_5 < _zz_dataOut_payload_224_21);
  assign _zz_dataOut_payload_224_43 = (_zz_dataOut_payload_224_42 ? _zz_dataOut_payload_224_5 : _zz_dataOut_payload_224_21);
  assign _zz_dataOut_payload_240_5 = (_zz_dataOut_payload_224_42 ? _zz_dataOut_payload_224_21 : _zz_dataOut_payload_224_5);
  assign _zz_dataOut_payload_224_44 = (_zz_dataOut_payload_224_6 < _zz_dataOut_payload_224_22);
  assign _zz_dataOut_payload_224_45 = (_zz_dataOut_payload_224_44 ? _zz_dataOut_payload_224_6 : _zz_dataOut_payload_224_22);
  assign _zz_dataOut_payload_240_6 = (_zz_dataOut_payload_224_44 ? _zz_dataOut_payload_224_22 : _zz_dataOut_payload_224_6);
  assign _zz_dataOut_payload_224_46 = (_zz_dataOut_payload_224_7 < _zz_dataOut_payload_224_23);
  assign _zz_dataOut_payload_224_47 = (_zz_dataOut_payload_224_46 ? _zz_dataOut_payload_224_7 : _zz_dataOut_payload_224_23);
  assign _zz_dataOut_payload_240_7 = (_zz_dataOut_payload_224_46 ? _zz_dataOut_payload_224_23 : _zz_dataOut_payload_224_7);
  assign _zz_dataOut_payload_224_48 = (_zz_dataOut_payload_224_8 < _zz_dataOut_payload_224_24);
  assign _zz_dataOut_payload_224_49 = (_zz_dataOut_payload_224_48 ? _zz_dataOut_payload_224_8 : _zz_dataOut_payload_224_24);
  assign _zz_dataOut_payload_240_8 = (_zz_dataOut_payload_224_48 ? _zz_dataOut_payload_224_24 : _zz_dataOut_payload_224_8);
  assign _zz_dataOut_payload_224_50 = (_zz_dataOut_payload_224_9 < _zz_dataOut_payload_224_25);
  assign _zz_dataOut_payload_224_51 = (_zz_dataOut_payload_224_50 ? _zz_dataOut_payload_224_9 : _zz_dataOut_payload_224_25);
  assign _zz_dataOut_payload_240_9 = (_zz_dataOut_payload_224_50 ? _zz_dataOut_payload_224_25 : _zz_dataOut_payload_224_9);
  assign _zz_dataOut_payload_224_52 = (_zz_dataOut_payload_224_10 < _zz_dataOut_payload_224_26);
  assign _zz_dataOut_payload_224_53 = (_zz_dataOut_payload_224_52 ? _zz_dataOut_payload_224_10 : _zz_dataOut_payload_224_26);
  assign _zz_dataOut_payload_240_10 = (_zz_dataOut_payload_224_52 ? _zz_dataOut_payload_224_26 : _zz_dataOut_payload_224_10);
  assign _zz_dataOut_payload_224_54 = (_zz_dataOut_payload_224_11 < _zz_dataOut_payload_224_27);
  assign _zz_dataOut_payload_224_55 = (_zz_dataOut_payload_224_54 ? _zz_dataOut_payload_224_11 : _zz_dataOut_payload_224_27);
  assign _zz_dataOut_payload_240_11 = (_zz_dataOut_payload_224_54 ? _zz_dataOut_payload_224_27 : _zz_dataOut_payload_224_11);
  assign _zz_dataOut_payload_224_56 = (_zz_dataOut_payload_224_12 < _zz_dataOut_payload_224_28);
  assign _zz_dataOut_payload_224_57 = (_zz_dataOut_payload_224_56 ? _zz_dataOut_payload_224_12 : _zz_dataOut_payload_224_28);
  assign _zz_dataOut_payload_240_12 = (_zz_dataOut_payload_224_56 ? _zz_dataOut_payload_224_28 : _zz_dataOut_payload_224_12);
  assign _zz_dataOut_payload_224_58 = (_zz_dataOut_payload_224_13 < _zz_dataOut_payload_224_29);
  assign _zz_dataOut_payload_224_59 = (_zz_dataOut_payload_224_58 ? _zz_dataOut_payload_224_13 : _zz_dataOut_payload_224_29);
  assign _zz_dataOut_payload_240_13 = (_zz_dataOut_payload_224_58 ? _zz_dataOut_payload_224_29 : _zz_dataOut_payload_224_13);
  assign _zz_dataOut_payload_224_60 = (_zz_dataOut_payload_224_14 < _zz_dataOut_payload_224_30);
  assign _zz_dataOut_payload_224_61 = (_zz_dataOut_payload_224_60 ? _zz_dataOut_payload_224_14 : _zz_dataOut_payload_224_30);
  assign _zz_dataOut_payload_240_14 = (_zz_dataOut_payload_224_60 ? _zz_dataOut_payload_224_30 : _zz_dataOut_payload_224_14);
  assign _zz_dataOut_payload_224_62 = (_zz_dataOut_payload_224_15 < _zz_dataOut_payload_224_31);
  assign _zz_dataOut_payload_224_63 = (_zz_dataOut_payload_224_62 ? _zz_dataOut_payload_224_15 : _zz_dataOut_payload_224_31);
  assign _zz_dataOut_payload_240_15 = (_zz_dataOut_payload_224_62 ? _zz_dataOut_payload_224_31 : _zz_dataOut_payload_224_15);
  assign _zz_dataOut_payload_224_64 = (_zz_dataOut_payload_224_33 < _zz_dataOut_payload_224_49);
  assign _zz_dataOut_payload_224_65 = (_zz_dataOut_payload_224_64 ? _zz_dataOut_payload_224_33 : _zz_dataOut_payload_224_49);
  assign _zz_dataOut_payload_232 = (_zz_dataOut_payload_224_64 ? _zz_dataOut_payload_224_49 : _zz_dataOut_payload_224_33);
  assign _zz_dataOut_payload_224_66 = (_zz_dataOut_payload_224_35 < _zz_dataOut_payload_224_51);
  assign _zz_dataOut_payload_224_67 = (_zz_dataOut_payload_224_66 ? _zz_dataOut_payload_224_35 : _zz_dataOut_payload_224_51);
  assign _zz_dataOut_payload_232_1 = (_zz_dataOut_payload_224_66 ? _zz_dataOut_payload_224_51 : _zz_dataOut_payload_224_35);
  assign _zz_dataOut_payload_224_68 = (_zz_dataOut_payload_224_37 < _zz_dataOut_payload_224_53);
  assign _zz_dataOut_payload_224_69 = (_zz_dataOut_payload_224_68 ? _zz_dataOut_payload_224_37 : _zz_dataOut_payload_224_53);
  assign _zz_dataOut_payload_232_2 = (_zz_dataOut_payload_224_68 ? _zz_dataOut_payload_224_53 : _zz_dataOut_payload_224_37);
  assign _zz_dataOut_payload_224_70 = (_zz_dataOut_payload_224_39 < _zz_dataOut_payload_224_55);
  assign _zz_dataOut_payload_224_71 = (_zz_dataOut_payload_224_70 ? _zz_dataOut_payload_224_39 : _zz_dataOut_payload_224_55);
  assign _zz_dataOut_payload_232_3 = (_zz_dataOut_payload_224_70 ? _zz_dataOut_payload_224_55 : _zz_dataOut_payload_224_39);
  assign _zz_dataOut_payload_224_72 = (_zz_dataOut_payload_224_41 < _zz_dataOut_payload_224_57);
  assign _zz_dataOut_payload_224_73 = (_zz_dataOut_payload_224_72 ? _zz_dataOut_payload_224_41 : _zz_dataOut_payload_224_57);
  assign _zz_dataOut_payload_232_4 = (_zz_dataOut_payload_224_72 ? _zz_dataOut_payload_224_57 : _zz_dataOut_payload_224_41);
  assign _zz_dataOut_payload_224_74 = (_zz_dataOut_payload_224_43 < _zz_dataOut_payload_224_59);
  assign _zz_dataOut_payload_224_75 = (_zz_dataOut_payload_224_74 ? _zz_dataOut_payload_224_43 : _zz_dataOut_payload_224_59);
  assign _zz_dataOut_payload_232_5 = (_zz_dataOut_payload_224_74 ? _zz_dataOut_payload_224_59 : _zz_dataOut_payload_224_43);
  assign _zz_dataOut_payload_224_76 = (_zz_dataOut_payload_224_45 < _zz_dataOut_payload_224_61);
  assign _zz_dataOut_payload_224_77 = (_zz_dataOut_payload_224_76 ? _zz_dataOut_payload_224_45 : _zz_dataOut_payload_224_61);
  assign _zz_dataOut_payload_232_6 = (_zz_dataOut_payload_224_76 ? _zz_dataOut_payload_224_61 : _zz_dataOut_payload_224_45);
  assign _zz_dataOut_payload_224_78 = (_zz_dataOut_payload_224_47 < _zz_dataOut_payload_224_63);
  assign _zz_dataOut_payload_224_79 = (_zz_dataOut_payload_224_78 ? _zz_dataOut_payload_224_47 : _zz_dataOut_payload_224_63);
  assign _zz_dataOut_payload_232_7 = (_zz_dataOut_payload_224_78 ? _zz_dataOut_payload_224_63 : _zz_dataOut_payload_224_47);
  assign _zz_dataOut_payload_224_80 = (_zz_dataOut_payload_224_65 < _zz_dataOut_payload_224_73);
  assign _zz_dataOut_payload_224_81 = (_zz_dataOut_payload_224_80 ? _zz_dataOut_payload_224_65 : _zz_dataOut_payload_224_73);
  assign _zz_dataOut_payload_228 = (_zz_dataOut_payload_224_80 ? _zz_dataOut_payload_224_73 : _zz_dataOut_payload_224_65);
  assign _zz_dataOut_payload_224_82 = (_zz_dataOut_payload_224_67 < _zz_dataOut_payload_224_75);
  assign _zz_dataOut_payload_224_83 = (_zz_dataOut_payload_224_82 ? _zz_dataOut_payload_224_67 : _zz_dataOut_payload_224_75);
  assign _zz_dataOut_payload_228_1 = (_zz_dataOut_payload_224_82 ? _zz_dataOut_payload_224_75 : _zz_dataOut_payload_224_67);
  assign _zz_dataOut_payload_224_84 = (_zz_dataOut_payload_224_69 < _zz_dataOut_payload_224_77);
  assign _zz_dataOut_payload_224_85 = (_zz_dataOut_payload_224_84 ? _zz_dataOut_payload_224_69 : _zz_dataOut_payload_224_77);
  assign _zz_dataOut_payload_228_2 = (_zz_dataOut_payload_224_84 ? _zz_dataOut_payload_224_77 : _zz_dataOut_payload_224_69);
  assign _zz_dataOut_payload_224_86 = (_zz_dataOut_payload_224_71 < _zz_dataOut_payload_224_79);
  assign _zz_dataOut_payload_224_87 = (_zz_dataOut_payload_224_86 ? _zz_dataOut_payload_224_71 : _zz_dataOut_payload_224_79);
  assign _zz_dataOut_payload_228_3 = (_zz_dataOut_payload_224_86 ? _zz_dataOut_payload_224_79 : _zz_dataOut_payload_224_71);
  assign _zz_dataOut_payload_224_88 = (_zz_dataOut_payload_224_81 < _zz_dataOut_payload_224_85);
  assign _zz_dataOut_payload_224_89 = (_zz_dataOut_payload_224_88 ? _zz_dataOut_payload_224_81 : _zz_dataOut_payload_224_85);
  assign _zz_dataOut_payload_226 = (_zz_dataOut_payload_224_88 ? _zz_dataOut_payload_224_85 : _zz_dataOut_payload_224_81);
  assign _zz_dataOut_payload_224_90 = (_zz_dataOut_payload_224_83 < _zz_dataOut_payload_224_87);
  assign _zz_dataOut_payload_224_91 = (_zz_dataOut_payload_224_90 ? _zz_dataOut_payload_224_83 : _zz_dataOut_payload_224_87);
  assign _zz_dataOut_payload_226_1 = (_zz_dataOut_payload_224_90 ? _zz_dataOut_payload_224_87 : _zz_dataOut_payload_224_83);
  assign _zz_dataOut_payload_224_92 = (_zz_dataOut_payload_224_89 < _zz_dataOut_payload_224_91);
  assign _zz_dataOut_payload_226_2 = (_zz_dataOut_payload_226 < _zz_dataOut_payload_226_1);
  assign _zz_dataOut_payload_228_4 = (_zz_dataOut_payload_228 < _zz_dataOut_payload_228_2);
  assign _zz_dataOut_payload_228_5 = (_zz_dataOut_payload_228_4 ? _zz_dataOut_payload_228 : _zz_dataOut_payload_228_2);
  assign _zz_dataOut_payload_230 = (_zz_dataOut_payload_228_4 ? _zz_dataOut_payload_228_2 : _zz_dataOut_payload_228);
  assign _zz_dataOut_payload_228_6 = (_zz_dataOut_payload_228_1 < _zz_dataOut_payload_228_3);
  assign _zz_dataOut_payload_228_7 = (_zz_dataOut_payload_228_6 ? _zz_dataOut_payload_228_1 : _zz_dataOut_payload_228_3);
  assign _zz_dataOut_payload_230_1 = (_zz_dataOut_payload_228_6 ? _zz_dataOut_payload_228_3 : _zz_dataOut_payload_228_1);
  assign _zz_dataOut_payload_228_8 = (_zz_dataOut_payload_228_5 < _zz_dataOut_payload_228_7);
  assign _zz_dataOut_payload_230_2 = (_zz_dataOut_payload_230 < _zz_dataOut_payload_230_1);
  assign _zz_dataOut_payload_232_8 = (_zz_dataOut_payload_232 < _zz_dataOut_payload_232_4);
  assign _zz_dataOut_payload_232_9 = (_zz_dataOut_payload_232_8 ? _zz_dataOut_payload_232 : _zz_dataOut_payload_232_4);
  assign _zz_dataOut_payload_236 = (_zz_dataOut_payload_232_8 ? _zz_dataOut_payload_232_4 : _zz_dataOut_payload_232);
  assign _zz_dataOut_payload_232_10 = (_zz_dataOut_payload_232_1 < _zz_dataOut_payload_232_5);
  assign _zz_dataOut_payload_232_11 = (_zz_dataOut_payload_232_10 ? _zz_dataOut_payload_232_1 : _zz_dataOut_payload_232_5);
  assign _zz_dataOut_payload_236_1 = (_zz_dataOut_payload_232_10 ? _zz_dataOut_payload_232_5 : _zz_dataOut_payload_232_1);
  assign _zz_dataOut_payload_232_12 = (_zz_dataOut_payload_232_2 < _zz_dataOut_payload_232_6);
  assign _zz_dataOut_payload_232_13 = (_zz_dataOut_payload_232_12 ? _zz_dataOut_payload_232_2 : _zz_dataOut_payload_232_6);
  assign _zz_dataOut_payload_236_2 = (_zz_dataOut_payload_232_12 ? _zz_dataOut_payload_232_6 : _zz_dataOut_payload_232_2);
  assign _zz_dataOut_payload_232_14 = (_zz_dataOut_payload_232_3 < _zz_dataOut_payload_232_7);
  assign _zz_dataOut_payload_232_15 = (_zz_dataOut_payload_232_14 ? _zz_dataOut_payload_232_3 : _zz_dataOut_payload_232_7);
  assign _zz_dataOut_payload_236_3 = (_zz_dataOut_payload_232_14 ? _zz_dataOut_payload_232_7 : _zz_dataOut_payload_232_3);
  assign _zz_dataOut_payload_232_16 = (_zz_dataOut_payload_232_9 < _zz_dataOut_payload_232_13);
  assign _zz_dataOut_payload_232_17 = (_zz_dataOut_payload_232_16 ? _zz_dataOut_payload_232_9 : _zz_dataOut_payload_232_13);
  assign _zz_dataOut_payload_234 = (_zz_dataOut_payload_232_16 ? _zz_dataOut_payload_232_13 : _zz_dataOut_payload_232_9);
  assign _zz_dataOut_payload_232_18 = (_zz_dataOut_payload_232_11 < _zz_dataOut_payload_232_15);
  assign _zz_dataOut_payload_232_19 = (_zz_dataOut_payload_232_18 ? _zz_dataOut_payload_232_11 : _zz_dataOut_payload_232_15);
  assign _zz_dataOut_payload_234_1 = (_zz_dataOut_payload_232_18 ? _zz_dataOut_payload_232_15 : _zz_dataOut_payload_232_11);
  assign _zz_dataOut_payload_232_20 = (_zz_dataOut_payload_232_17 < _zz_dataOut_payload_232_19);
  assign _zz_dataOut_payload_234_2 = (_zz_dataOut_payload_234 < _zz_dataOut_payload_234_1);
  assign _zz_dataOut_payload_236_4 = (_zz_dataOut_payload_236 < _zz_dataOut_payload_236_2);
  assign _zz_dataOut_payload_236_5 = (_zz_dataOut_payload_236_4 ? _zz_dataOut_payload_236 : _zz_dataOut_payload_236_2);
  assign _zz_dataOut_payload_238 = (_zz_dataOut_payload_236_4 ? _zz_dataOut_payload_236_2 : _zz_dataOut_payload_236);
  assign _zz_dataOut_payload_236_6 = (_zz_dataOut_payload_236_1 < _zz_dataOut_payload_236_3);
  assign _zz_dataOut_payload_236_7 = (_zz_dataOut_payload_236_6 ? _zz_dataOut_payload_236_1 : _zz_dataOut_payload_236_3);
  assign _zz_dataOut_payload_238_1 = (_zz_dataOut_payload_236_6 ? _zz_dataOut_payload_236_3 : _zz_dataOut_payload_236_1);
  assign _zz_dataOut_payload_236_8 = (_zz_dataOut_payload_236_5 < _zz_dataOut_payload_236_7);
  assign _zz_dataOut_payload_238_2 = (_zz_dataOut_payload_238 < _zz_dataOut_payload_238_1);
  assign _zz_dataOut_payload_240_16 = (_zz_dataOut_payload_240 < _zz_dataOut_payload_240_8);
  assign _zz_dataOut_payload_240_17 = (_zz_dataOut_payload_240_16 ? _zz_dataOut_payload_240 : _zz_dataOut_payload_240_8);
  assign _zz_dataOut_payload_248 = (_zz_dataOut_payload_240_16 ? _zz_dataOut_payload_240_8 : _zz_dataOut_payload_240);
  assign _zz_dataOut_payload_240_18 = (_zz_dataOut_payload_240_1 < _zz_dataOut_payload_240_9);
  assign _zz_dataOut_payload_240_19 = (_zz_dataOut_payload_240_18 ? _zz_dataOut_payload_240_1 : _zz_dataOut_payload_240_9);
  assign _zz_dataOut_payload_248_1 = (_zz_dataOut_payload_240_18 ? _zz_dataOut_payload_240_9 : _zz_dataOut_payload_240_1);
  assign _zz_dataOut_payload_240_20 = (_zz_dataOut_payload_240_2 < _zz_dataOut_payload_240_10);
  assign _zz_dataOut_payload_240_21 = (_zz_dataOut_payload_240_20 ? _zz_dataOut_payload_240_2 : _zz_dataOut_payload_240_10);
  assign _zz_dataOut_payload_248_2 = (_zz_dataOut_payload_240_20 ? _zz_dataOut_payload_240_10 : _zz_dataOut_payload_240_2);
  assign _zz_dataOut_payload_240_22 = (_zz_dataOut_payload_240_3 < _zz_dataOut_payload_240_11);
  assign _zz_dataOut_payload_240_23 = (_zz_dataOut_payload_240_22 ? _zz_dataOut_payload_240_3 : _zz_dataOut_payload_240_11);
  assign _zz_dataOut_payload_248_3 = (_zz_dataOut_payload_240_22 ? _zz_dataOut_payload_240_11 : _zz_dataOut_payload_240_3);
  assign _zz_dataOut_payload_240_24 = (_zz_dataOut_payload_240_4 < _zz_dataOut_payload_240_12);
  assign _zz_dataOut_payload_240_25 = (_zz_dataOut_payload_240_24 ? _zz_dataOut_payload_240_4 : _zz_dataOut_payload_240_12);
  assign _zz_dataOut_payload_248_4 = (_zz_dataOut_payload_240_24 ? _zz_dataOut_payload_240_12 : _zz_dataOut_payload_240_4);
  assign _zz_dataOut_payload_240_26 = (_zz_dataOut_payload_240_5 < _zz_dataOut_payload_240_13);
  assign _zz_dataOut_payload_240_27 = (_zz_dataOut_payload_240_26 ? _zz_dataOut_payload_240_5 : _zz_dataOut_payload_240_13);
  assign _zz_dataOut_payload_248_5 = (_zz_dataOut_payload_240_26 ? _zz_dataOut_payload_240_13 : _zz_dataOut_payload_240_5);
  assign _zz_dataOut_payload_240_28 = (_zz_dataOut_payload_240_6 < _zz_dataOut_payload_240_14);
  assign _zz_dataOut_payload_240_29 = (_zz_dataOut_payload_240_28 ? _zz_dataOut_payload_240_6 : _zz_dataOut_payload_240_14);
  assign _zz_dataOut_payload_248_6 = (_zz_dataOut_payload_240_28 ? _zz_dataOut_payload_240_14 : _zz_dataOut_payload_240_6);
  assign _zz_dataOut_payload_240_30 = (_zz_dataOut_payload_240_7 < _zz_dataOut_payload_240_15);
  assign _zz_dataOut_payload_240_31 = (_zz_dataOut_payload_240_30 ? _zz_dataOut_payload_240_7 : _zz_dataOut_payload_240_15);
  assign _zz_dataOut_payload_248_7 = (_zz_dataOut_payload_240_30 ? _zz_dataOut_payload_240_15 : _zz_dataOut_payload_240_7);
  assign _zz_dataOut_payload_240_32 = (_zz_dataOut_payload_240_17 < _zz_dataOut_payload_240_25);
  assign _zz_dataOut_payload_240_33 = (_zz_dataOut_payload_240_32 ? _zz_dataOut_payload_240_17 : _zz_dataOut_payload_240_25);
  assign _zz_dataOut_payload_244 = (_zz_dataOut_payload_240_32 ? _zz_dataOut_payload_240_25 : _zz_dataOut_payload_240_17);
  assign _zz_dataOut_payload_240_34 = (_zz_dataOut_payload_240_19 < _zz_dataOut_payload_240_27);
  assign _zz_dataOut_payload_240_35 = (_zz_dataOut_payload_240_34 ? _zz_dataOut_payload_240_19 : _zz_dataOut_payload_240_27);
  assign _zz_dataOut_payload_244_1 = (_zz_dataOut_payload_240_34 ? _zz_dataOut_payload_240_27 : _zz_dataOut_payload_240_19);
  assign _zz_dataOut_payload_240_36 = (_zz_dataOut_payload_240_21 < _zz_dataOut_payload_240_29);
  assign _zz_dataOut_payload_240_37 = (_zz_dataOut_payload_240_36 ? _zz_dataOut_payload_240_21 : _zz_dataOut_payload_240_29);
  assign _zz_dataOut_payload_244_2 = (_zz_dataOut_payload_240_36 ? _zz_dataOut_payload_240_29 : _zz_dataOut_payload_240_21);
  assign _zz_dataOut_payload_240_38 = (_zz_dataOut_payload_240_23 < _zz_dataOut_payload_240_31);
  assign _zz_dataOut_payload_240_39 = (_zz_dataOut_payload_240_38 ? _zz_dataOut_payload_240_23 : _zz_dataOut_payload_240_31);
  assign _zz_dataOut_payload_244_3 = (_zz_dataOut_payload_240_38 ? _zz_dataOut_payload_240_31 : _zz_dataOut_payload_240_23);
  assign _zz_dataOut_payload_240_40 = (_zz_dataOut_payload_240_33 < _zz_dataOut_payload_240_37);
  assign _zz_dataOut_payload_240_41 = (_zz_dataOut_payload_240_40 ? _zz_dataOut_payload_240_33 : _zz_dataOut_payload_240_37);
  assign _zz_dataOut_payload_242 = (_zz_dataOut_payload_240_40 ? _zz_dataOut_payload_240_37 : _zz_dataOut_payload_240_33);
  assign _zz_dataOut_payload_240_42 = (_zz_dataOut_payload_240_35 < _zz_dataOut_payload_240_39);
  assign _zz_dataOut_payload_240_43 = (_zz_dataOut_payload_240_42 ? _zz_dataOut_payload_240_35 : _zz_dataOut_payload_240_39);
  assign _zz_dataOut_payload_242_1 = (_zz_dataOut_payload_240_42 ? _zz_dataOut_payload_240_39 : _zz_dataOut_payload_240_35);
  assign _zz_dataOut_payload_240_44 = (_zz_dataOut_payload_240_41 < _zz_dataOut_payload_240_43);
  assign _zz_dataOut_payload_242_2 = (_zz_dataOut_payload_242 < _zz_dataOut_payload_242_1);
  assign _zz_dataOut_payload_244_4 = (_zz_dataOut_payload_244 < _zz_dataOut_payload_244_2);
  assign _zz_dataOut_payload_244_5 = (_zz_dataOut_payload_244_4 ? _zz_dataOut_payload_244 : _zz_dataOut_payload_244_2);
  assign _zz_dataOut_payload_246 = (_zz_dataOut_payload_244_4 ? _zz_dataOut_payload_244_2 : _zz_dataOut_payload_244);
  assign _zz_dataOut_payload_244_6 = (_zz_dataOut_payload_244_1 < _zz_dataOut_payload_244_3);
  assign _zz_dataOut_payload_244_7 = (_zz_dataOut_payload_244_6 ? _zz_dataOut_payload_244_1 : _zz_dataOut_payload_244_3);
  assign _zz_dataOut_payload_246_1 = (_zz_dataOut_payload_244_6 ? _zz_dataOut_payload_244_3 : _zz_dataOut_payload_244_1);
  assign _zz_dataOut_payload_244_8 = (_zz_dataOut_payload_244_5 < _zz_dataOut_payload_244_7);
  assign _zz_dataOut_payload_246_2 = (_zz_dataOut_payload_246 < _zz_dataOut_payload_246_1);
  assign _zz_dataOut_payload_248_8 = (_zz_dataOut_payload_248 < _zz_dataOut_payload_248_4);
  assign _zz_dataOut_payload_248_9 = (_zz_dataOut_payload_248_8 ? _zz_dataOut_payload_248 : _zz_dataOut_payload_248_4);
  assign _zz_dataOut_payload_252 = (_zz_dataOut_payload_248_8 ? _zz_dataOut_payload_248_4 : _zz_dataOut_payload_248);
  assign _zz_dataOut_payload_248_10 = (_zz_dataOut_payload_248_1 < _zz_dataOut_payload_248_5);
  assign _zz_dataOut_payload_248_11 = (_zz_dataOut_payload_248_10 ? _zz_dataOut_payload_248_1 : _zz_dataOut_payload_248_5);
  assign _zz_dataOut_payload_252_1 = (_zz_dataOut_payload_248_10 ? _zz_dataOut_payload_248_5 : _zz_dataOut_payload_248_1);
  assign _zz_dataOut_payload_248_12 = (_zz_dataOut_payload_248_2 < _zz_dataOut_payload_248_6);
  assign _zz_dataOut_payload_248_13 = (_zz_dataOut_payload_248_12 ? _zz_dataOut_payload_248_2 : _zz_dataOut_payload_248_6);
  assign _zz_dataOut_payload_252_2 = (_zz_dataOut_payload_248_12 ? _zz_dataOut_payload_248_6 : _zz_dataOut_payload_248_2);
  assign _zz_dataOut_payload_248_14 = (_zz_dataOut_payload_248_3 < _zz_dataOut_payload_248_7);
  assign _zz_dataOut_payload_248_15 = (_zz_dataOut_payload_248_14 ? _zz_dataOut_payload_248_3 : _zz_dataOut_payload_248_7);
  assign _zz_dataOut_payload_252_3 = (_zz_dataOut_payload_248_14 ? _zz_dataOut_payload_248_7 : _zz_dataOut_payload_248_3);
  assign _zz_dataOut_payload_248_16 = (_zz_dataOut_payload_248_9 < _zz_dataOut_payload_248_13);
  assign _zz_dataOut_payload_248_17 = (_zz_dataOut_payload_248_16 ? _zz_dataOut_payload_248_9 : _zz_dataOut_payload_248_13);
  assign _zz_dataOut_payload_250 = (_zz_dataOut_payload_248_16 ? _zz_dataOut_payload_248_13 : _zz_dataOut_payload_248_9);
  assign _zz_dataOut_payload_248_18 = (_zz_dataOut_payload_248_11 < _zz_dataOut_payload_248_15);
  assign _zz_dataOut_payload_248_19 = (_zz_dataOut_payload_248_18 ? _zz_dataOut_payload_248_11 : _zz_dataOut_payload_248_15);
  assign _zz_dataOut_payload_250_1 = (_zz_dataOut_payload_248_18 ? _zz_dataOut_payload_248_15 : _zz_dataOut_payload_248_11);
  assign _zz_dataOut_payload_248_20 = (_zz_dataOut_payload_248_17 < _zz_dataOut_payload_248_19);
  assign _zz_dataOut_payload_250_2 = (_zz_dataOut_payload_250 < _zz_dataOut_payload_250_1);
  assign _zz_dataOut_payload_252_4 = (_zz_dataOut_payload_252 < _zz_dataOut_payload_252_2);
  assign _zz_dataOut_payload_252_5 = (_zz_dataOut_payload_252_4 ? _zz_dataOut_payload_252 : _zz_dataOut_payload_252_2);
  assign _zz_dataOut_payload_254 = (_zz_dataOut_payload_252_4 ? _zz_dataOut_payload_252_2 : _zz_dataOut_payload_252);
  assign _zz_dataOut_payload_252_6 = (_zz_dataOut_payload_252_1 < _zz_dataOut_payload_252_3);
  assign _zz_dataOut_payload_252_7 = (_zz_dataOut_payload_252_6 ? _zz_dataOut_payload_252_1 : _zz_dataOut_payload_252_3);
  assign _zz_dataOut_payload_254_1 = (_zz_dataOut_payload_252_6 ? _zz_dataOut_payload_252_3 : _zz_dataOut_payload_252_1);
  assign _zz_dataOut_payload_252_8 = (_zz_dataOut_payload_252_5 < _zz_dataOut_payload_252_7);
  assign _zz_dataOut_payload_254_2 = (_zz_dataOut_payload_254 < _zz_dataOut_payload_254_1);
  assign dataOut_payload_0 = _zz_dataOut_payload_0_16644;
  assign dataOut_payload_1 = _zz_dataOut_payload_1_7;
  assign dataOut_payload_2 = _zz_dataOut_payload_2_10;
  assign dataOut_payload_3 = _zz_dataOut_payload_3_7;
  assign dataOut_payload_4 = _zz_dataOut_payload_4_16;
  assign dataOut_payload_5 = _zz_dataOut_payload_5_7;
  assign dataOut_payload_6 = _zz_dataOut_payload_6_10;
  assign dataOut_payload_7 = _zz_dataOut_payload_7_7;
  assign dataOut_payload_8 = _zz_dataOut_payload_8_28;
  assign dataOut_payload_9 = _zz_dataOut_payload_9_7;
  assign dataOut_payload_10 = _zz_dataOut_payload_10_10;
  assign dataOut_payload_11 = _zz_dataOut_payload_11_7;
  assign dataOut_payload_12 = _zz_dataOut_payload_12_16;
  assign dataOut_payload_13 = _zz_dataOut_payload_13_7;
  assign dataOut_payload_14 = _zz_dataOut_payload_14_10;
  assign dataOut_payload_15 = _zz_dataOut_payload_15_7;
  assign dataOut_payload_16 = _zz_dataOut_payload_16_52;
  assign dataOut_payload_17 = _zz_dataOut_payload_17_7;
  assign dataOut_payload_18 = _zz_dataOut_payload_18_10;
  assign dataOut_payload_19 = _zz_dataOut_payload_19_7;
  assign dataOut_payload_20 = _zz_dataOut_payload_20_16;
  assign dataOut_payload_21 = _zz_dataOut_payload_21_7;
  assign dataOut_payload_22 = _zz_dataOut_payload_22_10;
  assign dataOut_payload_23 = _zz_dataOut_payload_23_7;
  assign dataOut_payload_24 = _zz_dataOut_payload_24_28;
  assign dataOut_payload_25 = _zz_dataOut_payload_25_7;
  assign dataOut_payload_26 = _zz_dataOut_payload_26_10;
  assign dataOut_payload_27 = _zz_dataOut_payload_27_7;
  assign dataOut_payload_28 = _zz_dataOut_payload_28_16;
  assign dataOut_payload_29 = _zz_dataOut_payload_29_7;
  assign dataOut_payload_30 = _zz_dataOut_payload_30_10;
  assign dataOut_payload_31 = _zz_dataOut_payload_31_7;
  assign dataOut_payload_32 = _zz_dataOut_payload_32_100;
  assign dataOut_payload_33 = _zz_dataOut_payload_33_7;
  assign dataOut_payload_34 = _zz_dataOut_payload_34_10;
  assign dataOut_payload_35 = _zz_dataOut_payload_35_7;
  assign dataOut_payload_36 = _zz_dataOut_payload_36_16;
  assign dataOut_payload_37 = _zz_dataOut_payload_37_7;
  assign dataOut_payload_38 = _zz_dataOut_payload_38_10;
  assign dataOut_payload_39 = _zz_dataOut_payload_39_7;
  assign dataOut_payload_40 = _zz_dataOut_payload_40_28;
  assign dataOut_payload_41 = _zz_dataOut_payload_41_7;
  assign dataOut_payload_42 = _zz_dataOut_payload_42_10;
  assign dataOut_payload_43 = _zz_dataOut_payload_43_7;
  assign dataOut_payload_44 = _zz_dataOut_payload_44_16;
  assign dataOut_payload_45 = _zz_dataOut_payload_45_7;
  assign dataOut_payload_46 = _zz_dataOut_payload_46_10;
  assign dataOut_payload_47 = _zz_dataOut_payload_47_7;
  assign dataOut_payload_48 = _zz_dataOut_payload_48_52;
  assign dataOut_payload_49 = _zz_dataOut_payload_49_7;
  assign dataOut_payload_50 = _zz_dataOut_payload_50_10;
  assign dataOut_payload_51 = _zz_dataOut_payload_51_7;
  assign dataOut_payload_52 = _zz_dataOut_payload_52_16;
  assign dataOut_payload_53 = _zz_dataOut_payload_53_7;
  assign dataOut_payload_54 = _zz_dataOut_payload_54_10;
  assign dataOut_payload_55 = _zz_dataOut_payload_55_7;
  assign dataOut_payload_56 = _zz_dataOut_payload_56_28;
  assign dataOut_payload_57 = _zz_dataOut_payload_57_7;
  assign dataOut_payload_58 = _zz_dataOut_payload_58_10;
  assign dataOut_payload_59 = _zz_dataOut_payload_59_7;
  assign dataOut_payload_60 = _zz_dataOut_payload_60_16;
  assign dataOut_payload_61 = _zz_dataOut_payload_61_7;
  assign dataOut_payload_62 = _zz_dataOut_payload_62_10;
  assign dataOut_payload_63 = _zz_dataOut_payload_63_7;
  assign dataOut_payload_64 = _zz_dataOut_payload_64_196;
  assign dataOut_payload_65 = _zz_dataOut_payload_65_7;
  assign dataOut_payload_66 = _zz_dataOut_payload_66_10;
  assign dataOut_payload_67 = _zz_dataOut_payload_67_7;
  assign dataOut_payload_68 = _zz_dataOut_payload_68_16;
  assign dataOut_payload_69 = _zz_dataOut_payload_69_7;
  assign dataOut_payload_70 = _zz_dataOut_payload_70_10;
  assign dataOut_payload_71 = _zz_dataOut_payload_71_7;
  assign dataOut_payload_72 = _zz_dataOut_payload_72_28;
  assign dataOut_payload_73 = _zz_dataOut_payload_73_7;
  assign dataOut_payload_74 = _zz_dataOut_payload_74_10;
  assign dataOut_payload_75 = _zz_dataOut_payload_75_7;
  assign dataOut_payload_76 = _zz_dataOut_payload_76_16;
  assign dataOut_payload_77 = _zz_dataOut_payload_77_7;
  assign dataOut_payload_78 = _zz_dataOut_payload_78_10;
  assign dataOut_payload_79 = _zz_dataOut_payload_79_7;
  assign dataOut_payload_80 = _zz_dataOut_payload_80_52;
  assign dataOut_payload_81 = _zz_dataOut_payload_81_7;
  assign dataOut_payload_82 = _zz_dataOut_payload_82_10;
  assign dataOut_payload_83 = _zz_dataOut_payload_83_7;
  assign dataOut_payload_84 = _zz_dataOut_payload_84_16;
  assign dataOut_payload_85 = _zz_dataOut_payload_85_7;
  assign dataOut_payload_86 = _zz_dataOut_payload_86_10;
  assign dataOut_payload_87 = _zz_dataOut_payload_87_7;
  assign dataOut_payload_88 = _zz_dataOut_payload_88_28;
  assign dataOut_payload_89 = _zz_dataOut_payload_89_7;
  assign dataOut_payload_90 = _zz_dataOut_payload_90_10;
  assign dataOut_payload_91 = _zz_dataOut_payload_91_7;
  assign dataOut_payload_92 = _zz_dataOut_payload_92_16;
  assign dataOut_payload_93 = _zz_dataOut_payload_93_7;
  assign dataOut_payload_94 = _zz_dataOut_payload_94_10;
  assign dataOut_payload_95 = _zz_dataOut_payload_95_7;
  assign dataOut_payload_96 = _zz_dataOut_payload_96_100;
  assign dataOut_payload_97 = _zz_dataOut_payload_97_7;
  assign dataOut_payload_98 = _zz_dataOut_payload_98_10;
  assign dataOut_payload_99 = _zz_dataOut_payload_99_7;
  assign dataOut_payload_100 = _zz_dataOut_payload_100_16;
  assign dataOut_payload_101 = _zz_dataOut_payload_101_7;
  assign dataOut_payload_102 = _zz_dataOut_payload_102_10;
  assign dataOut_payload_103 = _zz_dataOut_payload_103_7;
  assign dataOut_payload_104 = _zz_dataOut_payload_104_28;
  assign dataOut_payload_105 = _zz_dataOut_payload_105_7;
  assign dataOut_payload_106 = _zz_dataOut_payload_106_10;
  assign dataOut_payload_107 = _zz_dataOut_payload_107_7;
  assign dataOut_payload_108 = _zz_dataOut_payload_108_16;
  assign dataOut_payload_109 = _zz_dataOut_payload_109_7;
  assign dataOut_payload_110 = _zz_dataOut_payload_110_10;
  assign dataOut_payload_111 = _zz_dataOut_payload_111_7;
  assign dataOut_payload_112 = _zz_dataOut_payload_112_52;
  assign dataOut_payload_113 = _zz_dataOut_payload_113_7;
  assign dataOut_payload_114 = _zz_dataOut_payload_114_10;
  assign dataOut_payload_115 = _zz_dataOut_payload_115_7;
  assign dataOut_payload_116 = _zz_dataOut_payload_116_16;
  assign dataOut_payload_117 = _zz_dataOut_payload_117_7;
  assign dataOut_payload_118 = _zz_dataOut_payload_118_10;
  assign dataOut_payload_119 = _zz_dataOut_payload_119_7;
  assign dataOut_payload_120 = _zz_dataOut_payload_120_28;
  assign dataOut_payload_121 = _zz_dataOut_payload_121_7;
  assign dataOut_payload_122 = _zz_dataOut_payload_122_10;
  assign dataOut_payload_123 = _zz_dataOut_payload_123_7;
  assign dataOut_payload_124 = _zz_dataOut_payload_124_16;
  assign dataOut_payload_125 = _zz_dataOut_payload_125_7;
  assign dataOut_payload_126 = _zz_dataOut_payload_126_10;
  assign dataOut_payload_127 = _zz_dataOut_payload_127_7;
  assign dataOut_payload_128 = _zz_dataOut_payload_128_388;
  assign dataOut_payload_129 = _zz_dataOut_payload_129_7;
  assign dataOut_payload_130 = _zz_dataOut_payload_130_10;
  assign dataOut_payload_131 = _zz_dataOut_payload_131_7;
  assign dataOut_payload_132 = _zz_dataOut_payload_132_16;
  assign dataOut_payload_133 = _zz_dataOut_payload_133_7;
  assign dataOut_payload_134 = _zz_dataOut_payload_134_10;
  assign dataOut_payload_135 = _zz_dataOut_payload_135_7;
  assign dataOut_payload_136 = _zz_dataOut_payload_136_28;
  assign dataOut_payload_137 = _zz_dataOut_payload_137_7;
  assign dataOut_payload_138 = _zz_dataOut_payload_138_10;
  assign dataOut_payload_139 = _zz_dataOut_payload_139_7;
  assign dataOut_payload_140 = _zz_dataOut_payload_140_16;
  assign dataOut_payload_141 = _zz_dataOut_payload_141_7;
  assign dataOut_payload_142 = _zz_dataOut_payload_142_10;
  assign dataOut_payload_143 = _zz_dataOut_payload_143_7;
  assign dataOut_payload_144 = _zz_dataOut_payload_144_52;
  assign dataOut_payload_145 = _zz_dataOut_payload_145_7;
  assign dataOut_payload_146 = _zz_dataOut_payload_146_10;
  assign dataOut_payload_147 = _zz_dataOut_payload_147_7;
  assign dataOut_payload_148 = _zz_dataOut_payload_148_16;
  assign dataOut_payload_149 = _zz_dataOut_payload_149_7;
  assign dataOut_payload_150 = _zz_dataOut_payload_150_10;
  assign dataOut_payload_151 = _zz_dataOut_payload_151_7;
  assign dataOut_payload_152 = _zz_dataOut_payload_152_28;
  assign dataOut_payload_153 = _zz_dataOut_payload_153_7;
  assign dataOut_payload_154 = _zz_dataOut_payload_154_10;
  assign dataOut_payload_155 = _zz_dataOut_payload_155_7;
  assign dataOut_payload_156 = _zz_dataOut_payload_156_16;
  assign dataOut_payload_157 = _zz_dataOut_payload_157_7;
  assign dataOut_payload_158 = _zz_dataOut_payload_158_10;
  assign dataOut_payload_159 = _zz_dataOut_payload_159_7;
  assign dataOut_payload_160 = _zz_dataOut_payload_160_100;
  assign dataOut_payload_161 = _zz_dataOut_payload_161_7;
  assign dataOut_payload_162 = _zz_dataOut_payload_162_10;
  assign dataOut_payload_163 = _zz_dataOut_payload_163_7;
  assign dataOut_payload_164 = _zz_dataOut_payload_164_16;
  assign dataOut_payload_165 = _zz_dataOut_payload_165_7;
  assign dataOut_payload_166 = _zz_dataOut_payload_166_10;
  assign dataOut_payload_167 = _zz_dataOut_payload_167_7;
  assign dataOut_payload_168 = _zz_dataOut_payload_168_28;
  assign dataOut_payload_169 = _zz_dataOut_payload_169_7;
  assign dataOut_payload_170 = _zz_dataOut_payload_170_10;
  assign dataOut_payload_171 = _zz_dataOut_payload_171_7;
  assign dataOut_payload_172 = _zz_dataOut_payload_172_16;
  assign dataOut_payload_173 = _zz_dataOut_payload_173_7;
  assign dataOut_payload_174 = _zz_dataOut_payload_174_10;
  assign dataOut_payload_175 = _zz_dataOut_payload_175_7;
  assign dataOut_payload_176 = _zz_dataOut_payload_176_52;
  assign dataOut_payload_177 = _zz_dataOut_payload_177_7;
  assign dataOut_payload_178 = _zz_dataOut_payload_178_10;
  assign dataOut_payload_179 = _zz_dataOut_payload_179_7;
  assign dataOut_payload_180 = _zz_dataOut_payload_180_16;
  assign dataOut_payload_181 = _zz_dataOut_payload_181_7;
  assign dataOut_payload_182 = _zz_dataOut_payload_182_10;
  assign dataOut_payload_183 = _zz_dataOut_payload_183_7;
  assign dataOut_payload_184 = _zz_dataOut_payload_184_28;
  assign dataOut_payload_185 = _zz_dataOut_payload_185_7;
  assign dataOut_payload_186 = _zz_dataOut_payload_186_10;
  assign dataOut_payload_187 = _zz_dataOut_payload_187_7;
  assign dataOut_payload_188 = _zz_dataOut_payload_188_16;
  assign dataOut_payload_189 = _zz_dataOut_payload_189_7;
  assign dataOut_payload_190 = _zz_dataOut_payload_190_10;
  assign dataOut_payload_191 = _zz_dataOut_payload_191_7;
  assign dataOut_payload_192 = _zz_dataOut_payload_192_196;
  assign dataOut_payload_193 = _zz_dataOut_payload_193_7;
  assign dataOut_payload_194 = _zz_dataOut_payload_194_10;
  assign dataOut_payload_195 = _zz_dataOut_payload_195_7;
  assign dataOut_payload_196 = _zz_dataOut_payload_196_16;
  assign dataOut_payload_197 = _zz_dataOut_payload_197_7;
  assign dataOut_payload_198 = _zz_dataOut_payload_198_10;
  assign dataOut_payload_199 = _zz_dataOut_payload_199_7;
  assign dataOut_payload_200 = _zz_dataOut_payload_200_28;
  assign dataOut_payload_201 = _zz_dataOut_payload_201_7;
  assign dataOut_payload_202 = _zz_dataOut_payload_202_10;
  assign dataOut_payload_203 = _zz_dataOut_payload_203_7;
  assign dataOut_payload_204 = _zz_dataOut_payload_204_16;
  assign dataOut_payload_205 = _zz_dataOut_payload_205_7;
  assign dataOut_payload_206 = _zz_dataOut_payload_206_10;
  assign dataOut_payload_207 = _zz_dataOut_payload_207_7;
  assign dataOut_payload_208 = _zz_dataOut_payload_208_52;
  assign dataOut_payload_209 = _zz_dataOut_payload_209_7;
  assign dataOut_payload_210 = _zz_dataOut_payload_210_10;
  assign dataOut_payload_211 = _zz_dataOut_payload_211_7;
  assign dataOut_payload_212 = _zz_dataOut_payload_212_16;
  assign dataOut_payload_213 = _zz_dataOut_payload_213_7;
  assign dataOut_payload_214 = _zz_dataOut_payload_214_10;
  assign dataOut_payload_215 = _zz_dataOut_payload_215_7;
  assign dataOut_payload_216 = _zz_dataOut_payload_216_28;
  assign dataOut_payload_217 = _zz_dataOut_payload_217_7;
  assign dataOut_payload_218 = _zz_dataOut_payload_218_10;
  assign dataOut_payload_219 = _zz_dataOut_payload_219_7;
  assign dataOut_payload_220 = _zz_dataOut_payload_220_16;
  assign dataOut_payload_221 = _zz_dataOut_payload_221_7;
  assign dataOut_payload_222 = _zz_dataOut_payload_222_10;
  assign dataOut_payload_223 = _zz_dataOut_payload_223_7;
  assign dataOut_payload_224 = _zz_dataOut_payload_224_100;
  assign dataOut_payload_225 = _zz_dataOut_payload_225_7;
  assign dataOut_payload_226 = _zz_dataOut_payload_226_10;
  assign dataOut_payload_227 = _zz_dataOut_payload_227_7;
  assign dataOut_payload_228 = _zz_dataOut_payload_228_16;
  assign dataOut_payload_229 = _zz_dataOut_payload_229_7;
  assign dataOut_payload_230 = _zz_dataOut_payload_230_10;
  assign dataOut_payload_231 = _zz_dataOut_payload_231_7;
  assign dataOut_payload_232 = _zz_dataOut_payload_232_28;
  assign dataOut_payload_233 = _zz_dataOut_payload_233_7;
  assign dataOut_payload_234 = _zz_dataOut_payload_234_10;
  assign dataOut_payload_235 = _zz_dataOut_payload_235_7;
  assign dataOut_payload_236 = _zz_dataOut_payload_236_16;
  assign dataOut_payload_237 = _zz_dataOut_payload_237_7;
  assign dataOut_payload_238 = _zz_dataOut_payload_238_10;
  assign dataOut_payload_239 = _zz_dataOut_payload_239_7;
  assign dataOut_payload_240 = _zz_dataOut_payload_240_52;
  assign dataOut_payload_241 = _zz_dataOut_payload_241_7;
  assign dataOut_payload_242 = _zz_dataOut_payload_242_10;
  assign dataOut_payload_243 = _zz_dataOut_payload_243_7;
  assign dataOut_payload_244 = _zz_dataOut_payload_244_16;
  assign dataOut_payload_245 = _zz_dataOut_payload_245_7;
  assign dataOut_payload_246 = _zz_dataOut_payload_246_10;
  assign dataOut_payload_247 = _zz_dataOut_payload_247_7;
  assign dataOut_payload_248 = _zz_dataOut_payload_248_28;
  assign dataOut_payload_249 = _zz_dataOut_payload_249_7;
  assign dataOut_payload_250 = _zz_dataOut_payload_250_10;
  assign dataOut_payload_251 = _zz_dataOut_payload_251_7;
  assign dataOut_payload_252 = _zz_dataOut_payload_252_16;
  assign dataOut_payload_253 = _zz_dataOut_payload_253_7;
  assign dataOut_payload_254 = _zz_dataOut_payload_254_10;
  assign dataOut_payload_255 = _zz_dataOut_payload_255_7;
  assign dataOut_valid = dataIn_valid_delay_36;
  always @(posedge clk) begin
    _zz_dataOut_payload_0_128 <= (_zz_dataOut_payload_0 ? dataIn_payload_0 : dataIn_payload_1);
    _zz_dataOut_payload_0_129 <= (_zz_dataOut_payload_0 ? dataIn_payload_1 : dataIn_payload_0);
    _zz_dataOut_payload_0_130 <= (_zz_dataOut_payload_0_1 ? dataIn_payload_2 : dataIn_payload_3);
    _zz_dataOut_payload_0_131 <= (_zz_dataOut_payload_0_1 ? dataIn_payload_3 : dataIn_payload_2);
    _zz_dataOut_payload_0_132 <= (_zz_dataOut_payload_0_2 ? dataIn_payload_4 : dataIn_payload_5);
    _zz_dataOut_payload_0_133 <= (_zz_dataOut_payload_0_2 ? dataIn_payload_5 : dataIn_payload_4);
    _zz_dataOut_payload_0_134 <= (_zz_dataOut_payload_0_3 ? dataIn_payload_6 : dataIn_payload_7);
    _zz_dataOut_payload_0_135 <= (_zz_dataOut_payload_0_3 ? dataIn_payload_7 : dataIn_payload_6);
    _zz_dataOut_payload_0_136 <= (_zz_dataOut_payload_0_4 ? dataIn_payload_8 : dataIn_payload_9);
    _zz_dataOut_payload_0_137 <= (_zz_dataOut_payload_0_4 ? dataIn_payload_9 : dataIn_payload_8);
    _zz_dataOut_payload_0_138 <= (_zz_dataOut_payload_0_5 ? dataIn_payload_10 : dataIn_payload_11);
    _zz_dataOut_payload_0_139 <= (_zz_dataOut_payload_0_5 ? dataIn_payload_11 : dataIn_payload_10);
    _zz_dataOut_payload_0_140 <= (_zz_dataOut_payload_0_6 ? dataIn_payload_12 : dataIn_payload_13);
    _zz_dataOut_payload_0_141 <= (_zz_dataOut_payload_0_6 ? dataIn_payload_13 : dataIn_payload_12);
    _zz_dataOut_payload_0_142 <= (_zz_dataOut_payload_0_7 ? dataIn_payload_14 : dataIn_payload_15);
    _zz_dataOut_payload_0_143 <= (_zz_dataOut_payload_0_7 ? dataIn_payload_15 : dataIn_payload_14);
    _zz_dataOut_payload_0_144 <= (_zz_dataOut_payload_0_8 ? dataIn_payload_16 : dataIn_payload_17);
    _zz_dataOut_payload_0_145 <= (_zz_dataOut_payload_0_8 ? dataIn_payload_17 : dataIn_payload_16);
    _zz_dataOut_payload_0_146 <= (_zz_dataOut_payload_0_9 ? dataIn_payload_18 : dataIn_payload_19);
    _zz_dataOut_payload_0_147 <= (_zz_dataOut_payload_0_9 ? dataIn_payload_19 : dataIn_payload_18);
    _zz_dataOut_payload_0_148 <= (_zz_dataOut_payload_0_10 ? dataIn_payload_20 : dataIn_payload_21);
    _zz_dataOut_payload_0_149 <= (_zz_dataOut_payload_0_10 ? dataIn_payload_21 : dataIn_payload_20);
    _zz_dataOut_payload_0_150 <= (_zz_dataOut_payload_0_11 ? dataIn_payload_22 : dataIn_payload_23);
    _zz_dataOut_payload_0_151 <= (_zz_dataOut_payload_0_11 ? dataIn_payload_23 : dataIn_payload_22);
    _zz_dataOut_payload_0_152 <= (_zz_dataOut_payload_0_12 ? dataIn_payload_24 : dataIn_payload_25);
    _zz_dataOut_payload_0_153 <= (_zz_dataOut_payload_0_12 ? dataIn_payload_25 : dataIn_payload_24);
    _zz_dataOut_payload_0_154 <= (_zz_dataOut_payload_0_13 ? dataIn_payload_26 : dataIn_payload_27);
    _zz_dataOut_payload_0_155 <= (_zz_dataOut_payload_0_13 ? dataIn_payload_27 : dataIn_payload_26);
    _zz_dataOut_payload_0_156 <= (_zz_dataOut_payload_0_14 ? dataIn_payload_28 : dataIn_payload_29);
    _zz_dataOut_payload_0_157 <= (_zz_dataOut_payload_0_14 ? dataIn_payload_29 : dataIn_payload_28);
    _zz_dataOut_payload_0_158 <= (_zz_dataOut_payload_0_15 ? dataIn_payload_30 : dataIn_payload_31);
    _zz_dataOut_payload_0_159 <= (_zz_dataOut_payload_0_15 ? dataIn_payload_31 : dataIn_payload_30);
    _zz_dataOut_payload_0_160 <= (_zz_dataOut_payload_0_16 ? dataIn_payload_32 : dataIn_payload_33);
    _zz_dataOut_payload_0_161 <= (_zz_dataOut_payload_0_16 ? dataIn_payload_33 : dataIn_payload_32);
    _zz_dataOut_payload_0_162 <= (_zz_dataOut_payload_0_17 ? dataIn_payload_34 : dataIn_payload_35);
    _zz_dataOut_payload_0_163 <= (_zz_dataOut_payload_0_17 ? dataIn_payload_35 : dataIn_payload_34);
    _zz_dataOut_payload_0_164 <= (_zz_dataOut_payload_0_18 ? dataIn_payload_36 : dataIn_payload_37);
    _zz_dataOut_payload_0_165 <= (_zz_dataOut_payload_0_18 ? dataIn_payload_37 : dataIn_payload_36);
    _zz_dataOut_payload_0_166 <= (_zz_dataOut_payload_0_19 ? dataIn_payload_38 : dataIn_payload_39);
    _zz_dataOut_payload_0_167 <= (_zz_dataOut_payload_0_19 ? dataIn_payload_39 : dataIn_payload_38);
    _zz_dataOut_payload_0_168 <= (_zz_dataOut_payload_0_20 ? dataIn_payload_40 : dataIn_payload_41);
    _zz_dataOut_payload_0_169 <= (_zz_dataOut_payload_0_20 ? dataIn_payload_41 : dataIn_payload_40);
    _zz_dataOut_payload_0_170 <= (_zz_dataOut_payload_0_21 ? dataIn_payload_42 : dataIn_payload_43);
    _zz_dataOut_payload_0_171 <= (_zz_dataOut_payload_0_21 ? dataIn_payload_43 : dataIn_payload_42);
    _zz_dataOut_payload_0_172 <= (_zz_dataOut_payload_0_22 ? dataIn_payload_44 : dataIn_payload_45);
    _zz_dataOut_payload_0_173 <= (_zz_dataOut_payload_0_22 ? dataIn_payload_45 : dataIn_payload_44);
    _zz_dataOut_payload_0_174 <= (_zz_dataOut_payload_0_23 ? dataIn_payload_46 : dataIn_payload_47);
    _zz_dataOut_payload_0_175 <= (_zz_dataOut_payload_0_23 ? dataIn_payload_47 : dataIn_payload_46);
    _zz_dataOut_payload_0_176 <= (_zz_dataOut_payload_0_24 ? dataIn_payload_48 : dataIn_payload_49);
    _zz_dataOut_payload_0_177 <= (_zz_dataOut_payload_0_24 ? dataIn_payload_49 : dataIn_payload_48);
    _zz_dataOut_payload_0_178 <= (_zz_dataOut_payload_0_25 ? dataIn_payload_50 : dataIn_payload_51);
    _zz_dataOut_payload_0_179 <= (_zz_dataOut_payload_0_25 ? dataIn_payload_51 : dataIn_payload_50);
    _zz_dataOut_payload_0_180 <= (_zz_dataOut_payload_0_26 ? dataIn_payload_52 : dataIn_payload_53);
    _zz_dataOut_payload_0_181 <= (_zz_dataOut_payload_0_26 ? dataIn_payload_53 : dataIn_payload_52);
    _zz_dataOut_payload_0_182 <= (_zz_dataOut_payload_0_27 ? dataIn_payload_54 : dataIn_payload_55);
    _zz_dataOut_payload_0_183 <= (_zz_dataOut_payload_0_27 ? dataIn_payload_55 : dataIn_payload_54);
    _zz_dataOut_payload_0_184 <= (_zz_dataOut_payload_0_28 ? dataIn_payload_56 : dataIn_payload_57);
    _zz_dataOut_payload_0_185 <= (_zz_dataOut_payload_0_28 ? dataIn_payload_57 : dataIn_payload_56);
    _zz_dataOut_payload_0_186 <= (_zz_dataOut_payload_0_29 ? dataIn_payload_58 : dataIn_payload_59);
    _zz_dataOut_payload_0_187 <= (_zz_dataOut_payload_0_29 ? dataIn_payload_59 : dataIn_payload_58);
    _zz_dataOut_payload_0_188 <= (_zz_dataOut_payload_0_30 ? dataIn_payload_60 : dataIn_payload_61);
    _zz_dataOut_payload_0_189 <= (_zz_dataOut_payload_0_30 ? dataIn_payload_61 : dataIn_payload_60);
    _zz_dataOut_payload_0_190 <= (_zz_dataOut_payload_0_31 ? dataIn_payload_62 : dataIn_payload_63);
    _zz_dataOut_payload_0_191 <= (_zz_dataOut_payload_0_31 ? dataIn_payload_63 : dataIn_payload_62);
    _zz_dataOut_payload_0_192 <= (_zz_dataOut_payload_0_32 ? dataIn_payload_64 : dataIn_payload_65);
    _zz_dataOut_payload_0_193 <= (_zz_dataOut_payload_0_32 ? dataIn_payload_65 : dataIn_payload_64);
    _zz_dataOut_payload_0_194 <= (_zz_dataOut_payload_0_33 ? dataIn_payload_66 : dataIn_payload_67);
    _zz_dataOut_payload_0_195 <= (_zz_dataOut_payload_0_33 ? dataIn_payload_67 : dataIn_payload_66);
    _zz_dataOut_payload_0_196 <= (_zz_dataOut_payload_0_34 ? dataIn_payload_68 : dataIn_payload_69);
    _zz_dataOut_payload_0_197 <= (_zz_dataOut_payload_0_34 ? dataIn_payload_69 : dataIn_payload_68);
    _zz_dataOut_payload_0_198 <= (_zz_dataOut_payload_0_35 ? dataIn_payload_70 : dataIn_payload_71);
    _zz_dataOut_payload_0_199 <= (_zz_dataOut_payload_0_35 ? dataIn_payload_71 : dataIn_payload_70);
    _zz_dataOut_payload_0_200 <= (_zz_dataOut_payload_0_36 ? dataIn_payload_72 : dataIn_payload_73);
    _zz_dataOut_payload_0_201 <= (_zz_dataOut_payload_0_36 ? dataIn_payload_73 : dataIn_payload_72);
    _zz_dataOut_payload_0_202 <= (_zz_dataOut_payload_0_37 ? dataIn_payload_74 : dataIn_payload_75);
    _zz_dataOut_payload_0_203 <= (_zz_dataOut_payload_0_37 ? dataIn_payload_75 : dataIn_payload_74);
    _zz_dataOut_payload_0_204 <= (_zz_dataOut_payload_0_38 ? dataIn_payload_76 : dataIn_payload_77);
    _zz_dataOut_payload_0_205 <= (_zz_dataOut_payload_0_38 ? dataIn_payload_77 : dataIn_payload_76);
    _zz_dataOut_payload_0_206 <= (_zz_dataOut_payload_0_39 ? dataIn_payload_78 : dataIn_payload_79);
    _zz_dataOut_payload_0_207 <= (_zz_dataOut_payload_0_39 ? dataIn_payload_79 : dataIn_payload_78);
    _zz_dataOut_payload_0_208 <= (_zz_dataOut_payload_0_40 ? dataIn_payload_80 : dataIn_payload_81);
    _zz_dataOut_payload_0_209 <= (_zz_dataOut_payload_0_40 ? dataIn_payload_81 : dataIn_payload_80);
    _zz_dataOut_payload_0_210 <= (_zz_dataOut_payload_0_41 ? dataIn_payload_82 : dataIn_payload_83);
    _zz_dataOut_payload_0_211 <= (_zz_dataOut_payload_0_41 ? dataIn_payload_83 : dataIn_payload_82);
    _zz_dataOut_payload_0_212 <= (_zz_dataOut_payload_0_42 ? dataIn_payload_84 : dataIn_payload_85);
    _zz_dataOut_payload_0_213 <= (_zz_dataOut_payload_0_42 ? dataIn_payload_85 : dataIn_payload_84);
    _zz_dataOut_payload_0_214 <= (_zz_dataOut_payload_0_43 ? dataIn_payload_86 : dataIn_payload_87);
    _zz_dataOut_payload_0_215 <= (_zz_dataOut_payload_0_43 ? dataIn_payload_87 : dataIn_payload_86);
    _zz_dataOut_payload_0_216 <= (_zz_dataOut_payload_0_44 ? dataIn_payload_88 : dataIn_payload_89);
    _zz_dataOut_payload_0_217 <= (_zz_dataOut_payload_0_44 ? dataIn_payload_89 : dataIn_payload_88);
    _zz_dataOut_payload_0_218 <= (_zz_dataOut_payload_0_45 ? dataIn_payload_90 : dataIn_payload_91);
    _zz_dataOut_payload_0_219 <= (_zz_dataOut_payload_0_45 ? dataIn_payload_91 : dataIn_payload_90);
    _zz_dataOut_payload_0_220 <= (_zz_dataOut_payload_0_46 ? dataIn_payload_92 : dataIn_payload_93);
    _zz_dataOut_payload_0_221 <= (_zz_dataOut_payload_0_46 ? dataIn_payload_93 : dataIn_payload_92);
    _zz_dataOut_payload_0_222 <= (_zz_dataOut_payload_0_47 ? dataIn_payload_94 : dataIn_payload_95);
    _zz_dataOut_payload_0_223 <= (_zz_dataOut_payload_0_47 ? dataIn_payload_95 : dataIn_payload_94);
    _zz_dataOut_payload_0_224 <= (_zz_dataOut_payload_0_48 ? dataIn_payload_96 : dataIn_payload_97);
    _zz_dataOut_payload_0_225 <= (_zz_dataOut_payload_0_48 ? dataIn_payload_97 : dataIn_payload_96);
    _zz_dataOut_payload_0_226 <= (_zz_dataOut_payload_0_49 ? dataIn_payload_98 : dataIn_payload_99);
    _zz_dataOut_payload_0_227 <= (_zz_dataOut_payload_0_49 ? dataIn_payload_99 : dataIn_payload_98);
    _zz_dataOut_payload_0_228 <= (_zz_dataOut_payload_0_50 ? dataIn_payload_100 : dataIn_payload_101);
    _zz_dataOut_payload_0_229 <= (_zz_dataOut_payload_0_50 ? dataIn_payload_101 : dataIn_payload_100);
    _zz_dataOut_payload_0_230 <= (_zz_dataOut_payload_0_51 ? dataIn_payload_102 : dataIn_payload_103);
    _zz_dataOut_payload_0_231 <= (_zz_dataOut_payload_0_51 ? dataIn_payload_103 : dataIn_payload_102);
    _zz_dataOut_payload_0_232 <= (_zz_dataOut_payload_0_52 ? dataIn_payload_104 : dataIn_payload_105);
    _zz_dataOut_payload_0_233 <= (_zz_dataOut_payload_0_52 ? dataIn_payload_105 : dataIn_payload_104);
    _zz_dataOut_payload_0_234 <= (_zz_dataOut_payload_0_53 ? dataIn_payload_106 : dataIn_payload_107);
    _zz_dataOut_payload_0_235 <= (_zz_dataOut_payload_0_53 ? dataIn_payload_107 : dataIn_payload_106);
    _zz_dataOut_payload_0_236 <= (_zz_dataOut_payload_0_54 ? dataIn_payload_108 : dataIn_payload_109);
    _zz_dataOut_payload_0_237 <= (_zz_dataOut_payload_0_54 ? dataIn_payload_109 : dataIn_payload_108);
    _zz_dataOut_payload_0_238 <= (_zz_dataOut_payload_0_55 ? dataIn_payload_110 : dataIn_payload_111);
    _zz_dataOut_payload_0_239 <= (_zz_dataOut_payload_0_55 ? dataIn_payload_111 : dataIn_payload_110);
    _zz_dataOut_payload_0_240 <= (_zz_dataOut_payload_0_56 ? dataIn_payload_112 : dataIn_payload_113);
    _zz_dataOut_payload_0_241 <= (_zz_dataOut_payload_0_56 ? dataIn_payload_113 : dataIn_payload_112);
    _zz_dataOut_payload_0_242 <= (_zz_dataOut_payload_0_57 ? dataIn_payload_114 : dataIn_payload_115);
    _zz_dataOut_payload_0_243 <= (_zz_dataOut_payload_0_57 ? dataIn_payload_115 : dataIn_payload_114);
    _zz_dataOut_payload_0_244 <= (_zz_dataOut_payload_0_58 ? dataIn_payload_116 : dataIn_payload_117);
    _zz_dataOut_payload_0_245 <= (_zz_dataOut_payload_0_58 ? dataIn_payload_117 : dataIn_payload_116);
    _zz_dataOut_payload_0_246 <= (_zz_dataOut_payload_0_59 ? dataIn_payload_118 : dataIn_payload_119);
    _zz_dataOut_payload_0_247 <= (_zz_dataOut_payload_0_59 ? dataIn_payload_119 : dataIn_payload_118);
    _zz_dataOut_payload_0_248 <= (_zz_dataOut_payload_0_60 ? dataIn_payload_120 : dataIn_payload_121);
    _zz_dataOut_payload_0_249 <= (_zz_dataOut_payload_0_60 ? dataIn_payload_121 : dataIn_payload_120);
    _zz_dataOut_payload_0_250 <= (_zz_dataOut_payload_0_61 ? dataIn_payload_122 : dataIn_payload_123);
    _zz_dataOut_payload_0_251 <= (_zz_dataOut_payload_0_61 ? dataIn_payload_123 : dataIn_payload_122);
    _zz_dataOut_payload_0_252 <= (_zz_dataOut_payload_0_62 ? dataIn_payload_124 : dataIn_payload_125);
    _zz_dataOut_payload_0_253 <= (_zz_dataOut_payload_0_62 ? dataIn_payload_125 : dataIn_payload_124);
    _zz_dataOut_payload_0_254 <= (_zz_dataOut_payload_0_63 ? dataIn_payload_126 : dataIn_payload_127);
    _zz_dataOut_payload_0_255 <= (_zz_dataOut_payload_0_63 ? dataIn_payload_127 : dataIn_payload_126);
    _zz_dataOut_payload_0_256 <= (_zz_dataOut_payload_0_64 ? dataIn_payload_128 : dataIn_payload_129);
    _zz_dataOut_payload_0_257 <= (_zz_dataOut_payload_0_64 ? dataIn_payload_129 : dataIn_payload_128);
    _zz_dataOut_payload_0_258 <= (_zz_dataOut_payload_0_65 ? dataIn_payload_130 : dataIn_payload_131);
    _zz_dataOut_payload_0_259 <= (_zz_dataOut_payload_0_65 ? dataIn_payload_131 : dataIn_payload_130);
    _zz_dataOut_payload_0_260 <= (_zz_dataOut_payload_0_66 ? dataIn_payload_132 : dataIn_payload_133);
    _zz_dataOut_payload_0_261 <= (_zz_dataOut_payload_0_66 ? dataIn_payload_133 : dataIn_payload_132);
    _zz_dataOut_payload_0_262 <= (_zz_dataOut_payload_0_67 ? dataIn_payload_134 : dataIn_payload_135);
    _zz_dataOut_payload_0_263 <= (_zz_dataOut_payload_0_67 ? dataIn_payload_135 : dataIn_payload_134);
    _zz_dataOut_payload_0_264 <= (_zz_dataOut_payload_0_68 ? dataIn_payload_136 : dataIn_payload_137);
    _zz_dataOut_payload_0_265 <= (_zz_dataOut_payload_0_68 ? dataIn_payload_137 : dataIn_payload_136);
    _zz_dataOut_payload_0_266 <= (_zz_dataOut_payload_0_69 ? dataIn_payload_138 : dataIn_payload_139);
    _zz_dataOut_payload_0_267 <= (_zz_dataOut_payload_0_69 ? dataIn_payload_139 : dataIn_payload_138);
    _zz_dataOut_payload_0_268 <= (_zz_dataOut_payload_0_70 ? dataIn_payload_140 : dataIn_payload_141);
    _zz_dataOut_payload_0_269 <= (_zz_dataOut_payload_0_70 ? dataIn_payload_141 : dataIn_payload_140);
    _zz_dataOut_payload_0_270 <= (_zz_dataOut_payload_0_71 ? dataIn_payload_142 : dataIn_payload_143);
    _zz_dataOut_payload_0_271 <= (_zz_dataOut_payload_0_71 ? dataIn_payload_143 : dataIn_payload_142);
    _zz_dataOut_payload_0_272 <= (_zz_dataOut_payload_0_72 ? dataIn_payload_144 : dataIn_payload_145);
    _zz_dataOut_payload_0_273 <= (_zz_dataOut_payload_0_72 ? dataIn_payload_145 : dataIn_payload_144);
    _zz_dataOut_payload_0_274 <= (_zz_dataOut_payload_0_73 ? dataIn_payload_146 : dataIn_payload_147);
    _zz_dataOut_payload_0_275 <= (_zz_dataOut_payload_0_73 ? dataIn_payload_147 : dataIn_payload_146);
    _zz_dataOut_payload_0_276 <= (_zz_dataOut_payload_0_74 ? dataIn_payload_148 : dataIn_payload_149);
    _zz_dataOut_payload_0_277 <= (_zz_dataOut_payload_0_74 ? dataIn_payload_149 : dataIn_payload_148);
    _zz_dataOut_payload_0_278 <= (_zz_dataOut_payload_0_75 ? dataIn_payload_150 : dataIn_payload_151);
    _zz_dataOut_payload_0_279 <= (_zz_dataOut_payload_0_75 ? dataIn_payload_151 : dataIn_payload_150);
    _zz_dataOut_payload_0_280 <= (_zz_dataOut_payload_0_76 ? dataIn_payload_152 : dataIn_payload_153);
    _zz_dataOut_payload_0_281 <= (_zz_dataOut_payload_0_76 ? dataIn_payload_153 : dataIn_payload_152);
    _zz_dataOut_payload_0_282 <= (_zz_dataOut_payload_0_77 ? dataIn_payload_154 : dataIn_payload_155);
    _zz_dataOut_payload_0_283 <= (_zz_dataOut_payload_0_77 ? dataIn_payload_155 : dataIn_payload_154);
    _zz_dataOut_payload_0_284 <= (_zz_dataOut_payload_0_78 ? dataIn_payload_156 : dataIn_payload_157);
    _zz_dataOut_payload_0_285 <= (_zz_dataOut_payload_0_78 ? dataIn_payload_157 : dataIn_payload_156);
    _zz_dataOut_payload_0_286 <= (_zz_dataOut_payload_0_79 ? dataIn_payload_158 : dataIn_payload_159);
    _zz_dataOut_payload_0_287 <= (_zz_dataOut_payload_0_79 ? dataIn_payload_159 : dataIn_payload_158);
    _zz_dataOut_payload_0_288 <= (_zz_dataOut_payload_0_80 ? dataIn_payload_160 : dataIn_payload_161);
    _zz_dataOut_payload_0_289 <= (_zz_dataOut_payload_0_80 ? dataIn_payload_161 : dataIn_payload_160);
    _zz_dataOut_payload_0_290 <= (_zz_dataOut_payload_0_81 ? dataIn_payload_162 : dataIn_payload_163);
    _zz_dataOut_payload_0_291 <= (_zz_dataOut_payload_0_81 ? dataIn_payload_163 : dataIn_payload_162);
    _zz_dataOut_payload_0_292 <= (_zz_dataOut_payload_0_82 ? dataIn_payload_164 : dataIn_payload_165);
    _zz_dataOut_payload_0_293 <= (_zz_dataOut_payload_0_82 ? dataIn_payload_165 : dataIn_payload_164);
    _zz_dataOut_payload_0_294 <= (_zz_dataOut_payload_0_83 ? dataIn_payload_166 : dataIn_payload_167);
    _zz_dataOut_payload_0_295 <= (_zz_dataOut_payload_0_83 ? dataIn_payload_167 : dataIn_payload_166);
    _zz_dataOut_payload_0_296 <= (_zz_dataOut_payload_0_84 ? dataIn_payload_168 : dataIn_payload_169);
    _zz_dataOut_payload_0_297 <= (_zz_dataOut_payload_0_84 ? dataIn_payload_169 : dataIn_payload_168);
    _zz_dataOut_payload_0_298 <= (_zz_dataOut_payload_0_85 ? dataIn_payload_170 : dataIn_payload_171);
    _zz_dataOut_payload_0_299 <= (_zz_dataOut_payload_0_85 ? dataIn_payload_171 : dataIn_payload_170);
    _zz_dataOut_payload_0_300 <= (_zz_dataOut_payload_0_86 ? dataIn_payload_172 : dataIn_payload_173);
    _zz_dataOut_payload_0_301 <= (_zz_dataOut_payload_0_86 ? dataIn_payload_173 : dataIn_payload_172);
    _zz_dataOut_payload_0_302 <= (_zz_dataOut_payload_0_87 ? dataIn_payload_174 : dataIn_payload_175);
    _zz_dataOut_payload_0_303 <= (_zz_dataOut_payload_0_87 ? dataIn_payload_175 : dataIn_payload_174);
    _zz_dataOut_payload_0_304 <= (_zz_dataOut_payload_0_88 ? dataIn_payload_176 : dataIn_payload_177);
    _zz_dataOut_payload_0_305 <= (_zz_dataOut_payload_0_88 ? dataIn_payload_177 : dataIn_payload_176);
    _zz_dataOut_payload_0_306 <= (_zz_dataOut_payload_0_89 ? dataIn_payload_178 : dataIn_payload_179);
    _zz_dataOut_payload_0_307 <= (_zz_dataOut_payload_0_89 ? dataIn_payload_179 : dataIn_payload_178);
    _zz_dataOut_payload_0_308 <= (_zz_dataOut_payload_0_90 ? dataIn_payload_180 : dataIn_payload_181);
    _zz_dataOut_payload_0_309 <= (_zz_dataOut_payload_0_90 ? dataIn_payload_181 : dataIn_payload_180);
    _zz_dataOut_payload_0_310 <= (_zz_dataOut_payload_0_91 ? dataIn_payload_182 : dataIn_payload_183);
    _zz_dataOut_payload_0_311 <= (_zz_dataOut_payload_0_91 ? dataIn_payload_183 : dataIn_payload_182);
    _zz_dataOut_payload_0_312 <= (_zz_dataOut_payload_0_92 ? dataIn_payload_184 : dataIn_payload_185);
    _zz_dataOut_payload_0_313 <= (_zz_dataOut_payload_0_92 ? dataIn_payload_185 : dataIn_payload_184);
    _zz_dataOut_payload_0_314 <= (_zz_dataOut_payload_0_93 ? dataIn_payload_186 : dataIn_payload_187);
    _zz_dataOut_payload_0_315 <= (_zz_dataOut_payload_0_93 ? dataIn_payload_187 : dataIn_payload_186);
    _zz_dataOut_payload_0_316 <= (_zz_dataOut_payload_0_94 ? dataIn_payload_188 : dataIn_payload_189);
    _zz_dataOut_payload_0_317 <= (_zz_dataOut_payload_0_94 ? dataIn_payload_189 : dataIn_payload_188);
    _zz_dataOut_payload_0_318 <= (_zz_dataOut_payload_0_95 ? dataIn_payload_190 : dataIn_payload_191);
    _zz_dataOut_payload_0_319 <= (_zz_dataOut_payload_0_95 ? dataIn_payload_191 : dataIn_payload_190);
    _zz_dataOut_payload_0_320 <= (_zz_dataOut_payload_0_96 ? dataIn_payload_192 : dataIn_payload_193);
    _zz_dataOut_payload_0_321 <= (_zz_dataOut_payload_0_96 ? dataIn_payload_193 : dataIn_payload_192);
    _zz_dataOut_payload_0_322 <= (_zz_dataOut_payload_0_97 ? dataIn_payload_194 : dataIn_payload_195);
    _zz_dataOut_payload_0_323 <= (_zz_dataOut_payload_0_97 ? dataIn_payload_195 : dataIn_payload_194);
    _zz_dataOut_payload_0_324 <= (_zz_dataOut_payload_0_98 ? dataIn_payload_196 : dataIn_payload_197);
    _zz_dataOut_payload_0_325 <= (_zz_dataOut_payload_0_98 ? dataIn_payload_197 : dataIn_payload_196);
    _zz_dataOut_payload_0_326 <= (_zz_dataOut_payload_0_99 ? dataIn_payload_198 : dataIn_payload_199);
    _zz_dataOut_payload_0_327 <= (_zz_dataOut_payload_0_99 ? dataIn_payload_199 : dataIn_payload_198);
    _zz_dataOut_payload_0_328 <= (_zz_dataOut_payload_0_100 ? dataIn_payload_200 : dataIn_payload_201);
    _zz_dataOut_payload_0_329 <= (_zz_dataOut_payload_0_100 ? dataIn_payload_201 : dataIn_payload_200);
    _zz_dataOut_payload_0_330 <= (_zz_dataOut_payload_0_101 ? dataIn_payload_202 : dataIn_payload_203);
    _zz_dataOut_payload_0_331 <= (_zz_dataOut_payload_0_101 ? dataIn_payload_203 : dataIn_payload_202);
    _zz_dataOut_payload_0_332 <= (_zz_dataOut_payload_0_102 ? dataIn_payload_204 : dataIn_payload_205);
    _zz_dataOut_payload_0_333 <= (_zz_dataOut_payload_0_102 ? dataIn_payload_205 : dataIn_payload_204);
    _zz_dataOut_payload_0_334 <= (_zz_dataOut_payload_0_103 ? dataIn_payload_206 : dataIn_payload_207);
    _zz_dataOut_payload_0_335 <= (_zz_dataOut_payload_0_103 ? dataIn_payload_207 : dataIn_payload_206);
    _zz_dataOut_payload_0_336 <= (_zz_dataOut_payload_0_104 ? dataIn_payload_208 : dataIn_payload_209);
    _zz_dataOut_payload_0_337 <= (_zz_dataOut_payload_0_104 ? dataIn_payload_209 : dataIn_payload_208);
    _zz_dataOut_payload_0_338 <= (_zz_dataOut_payload_0_105 ? dataIn_payload_210 : dataIn_payload_211);
    _zz_dataOut_payload_0_339 <= (_zz_dataOut_payload_0_105 ? dataIn_payload_211 : dataIn_payload_210);
    _zz_dataOut_payload_0_340 <= (_zz_dataOut_payload_0_106 ? dataIn_payload_212 : dataIn_payload_213);
    _zz_dataOut_payload_0_341 <= (_zz_dataOut_payload_0_106 ? dataIn_payload_213 : dataIn_payload_212);
    _zz_dataOut_payload_0_342 <= (_zz_dataOut_payload_0_107 ? dataIn_payload_214 : dataIn_payload_215);
    _zz_dataOut_payload_0_343 <= (_zz_dataOut_payload_0_107 ? dataIn_payload_215 : dataIn_payload_214);
    _zz_dataOut_payload_0_344 <= (_zz_dataOut_payload_0_108 ? dataIn_payload_216 : dataIn_payload_217);
    _zz_dataOut_payload_0_345 <= (_zz_dataOut_payload_0_108 ? dataIn_payload_217 : dataIn_payload_216);
    _zz_dataOut_payload_0_346 <= (_zz_dataOut_payload_0_109 ? dataIn_payload_218 : dataIn_payload_219);
    _zz_dataOut_payload_0_347 <= (_zz_dataOut_payload_0_109 ? dataIn_payload_219 : dataIn_payload_218);
    _zz_dataOut_payload_0_348 <= (_zz_dataOut_payload_0_110 ? dataIn_payload_220 : dataIn_payload_221);
    _zz_dataOut_payload_0_349 <= (_zz_dataOut_payload_0_110 ? dataIn_payload_221 : dataIn_payload_220);
    _zz_dataOut_payload_0_350 <= (_zz_dataOut_payload_0_111 ? dataIn_payload_222 : dataIn_payload_223);
    _zz_dataOut_payload_0_351 <= (_zz_dataOut_payload_0_111 ? dataIn_payload_223 : dataIn_payload_222);
    _zz_dataOut_payload_0_352 <= (_zz_dataOut_payload_0_112 ? dataIn_payload_224 : dataIn_payload_225);
    _zz_dataOut_payload_0_353 <= (_zz_dataOut_payload_0_112 ? dataIn_payload_225 : dataIn_payload_224);
    _zz_dataOut_payload_0_354 <= (_zz_dataOut_payload_0_113 ? dataIn_payload_226 : dataIn_payload_227);
    _zz_dataOut_payload_0_355 <= (_zz_dataOut_payload_0_113 ? dataIn_payload_227 : dataIn_payload_226);
    _zz_dataOut_payload_0_356 <= (_zz_dataOut_payload_0_114 ? dataIn_payload_228 : dataIn_payload_229);
    _zz_dataOut_payload_0_357 <= (_zz_dataOut_payload_0_114 ? dataIn_payload_229 : dataIn_payload_228);
    _zz_dataOut_payload_0_358 <= (_zz_dataOut_payload_0_115 ? dataIn_payload_230 : dataIn_payload_231);
    _zz_dataOut_payload_0_359 <= (_zz_dataOut_payload_0_115 ? dataIn_payload_231 : dataIn_payload_230);
    _zz_dataOut_payload_0_360 <= (_zz_dataOut_payload_0_116 ? dataIn_payload_232 : dataIn_payload_233);
    _zz_dataOut_payload_0_361 <= (_zz_dataOut_payload_0_116 ? dataIn_payload_233 : dataIn_payload_232);
    _zz_dataOut_payload_0_362 <= (_zz_dataOut_payload_0_117 ? dataIn_payload_234 : dataIn_payload_235);
    _zz_dataOut_payload_0_363 <= (_zz_dataOut_payload_0_117 ? dataIn_payload_235 : dataIn_payload_234);
    _zz_dataOut_payload_0_364 <= (_zz_dataOut_payload_0_118 ? dataIn_payload_236 : dataIn_payload_237);
    _zz_dataOut_payload_0_365 <= (_zz_dataOut_payload_0_118 ? dataIn_payload_237 : dataIn_payload_236);
    _zz_dataOut_payload_0_366 <= (_zz_dataOut_payload_0_119 ? dataIn_payload_238 : dataIn_payload_239);
    _zz_dataOut_payload_0_367 <= (_zz_dataOut_payload_0_119 ? dataIn_payload_239 : dataIn_payload_238);
    _zz_dataOut_payload_0_368 <= (_zz_dataOut_payload_0_120 ? dataIn_payload_240 : dataIn_payload_241);
    _zz_dataOut_payload_0_369 <= (_zz_dataOut_payload_0_120 ? dataIn_payload_241 : dataIn_payload_240);
    _zz_dataOut_payload_0_370 <= (_zz_dataOut_payload_0_121 ? dataIn_payload_242 : dataIn_payload_243);
    _zz_dataOut_payload_0_371 <= (_zz_dataOut_payload_0_121 ? dataIn_payload_243 : dataIn_payload_242);
    _zz_dataOut_payload_0_372 <= (_zz_dataOut_payload_0_122 ? dataIn_payload_244 : dataIn_payload_245);
    _zz_dataOut_payload_0_373 <= (_zz_dataOut_payload_0_122 ? dataIn_payload_245 : dataIn_payload_244);
    _zz_dataOut_payload_0_374 <= (_zz_dataOut_payload_0_123 ? dataIn_payload_246 : dataIn_payload_247);
    _zz_dataOut_payload_0_375 <= (_zz_dataOut_payload_0_123 ? dataIn_payload_247 : dataIn_payload_246);
    _zz_dataOut_payload_0_376 <= (_zz_dataOut_payload_0_124 ? dataIn_payload_248 : dataIn_payload_249);
    _zz_dataOut_payload_0_377 <= (_zz_dataOut_payload_0_124 ? dataIn_payload_249 : dataIn_payload_248);
    _zz_dataOut_payload_0_378 <= (_zz_dataOut_payload_0_125 ? dataIn_payload_250 : dataIn_payload_251);
    _zz_dataOut_payload_0_379 <= (_zz_dataOut_payload_0_125 ? dataIn_payload_251 : dataIn_payload_250);
    _zz_dataOut_payload_0_380 <= (_zz_dataOut_payload_0_126 ? dataIn_payload_252 : dataIn_payload_253);
    _zz_dataOut_payload_0_381 <= (_zz_dataOut_payload_0_126 ? dataIn_payload_253 : dataIn_payload_252);
    _zz_dataOut_payload_0_382 <= (_zz_dataOut_payload_0_127 ? dataIn_payload_254 : dataIn_payload_255);
    _zz_dataOut_payload_0_383 <= (_zz_dataOut_payload_0_127 ? dataIn_payload_255 : dataIn_payload_254);
    _zz_dataOut_payload_0_392 <= (_zz_dataOut_payload_0_390 ? _zz_dataOut_payload_0_385 : _zz_dataOut_payload_0_388);
    _zz_dataOut_payload_0_393 <= (_zz_dataOut_payload_0_390 ? _zz_dataOut_payload_0_388 : _zz_dataOut_payload_0_385);
    _zz_dataOut_payload_0_394 <= (_zz_dataOut_payload_0_391 ? _zz_dataOut_payload_0_389 : _zz_dataOut_payload_0_386);
    _zz_dataOut_payload_0_395 <= (_zz_dataOut_payload_0_391 ? _zz_dataOut_payload_0_386 : _zz_dataOut_payload_0_389);
    _zz_dataOut_payload_0_404 <= (_zz_dataOut_payload_0_402 ? _zz_dataOut_payload_0_397 : _zz_dataOut_payload_0_400);
    _zz_dataOut_payload_0_405 <= (_zz_dataOut_payload_0_402 ? _zz_dataOut_payload_0_400 : _zz_dataOut_payload_0_397);
    _zz_dataOut_payload_0_406 <= (_zz_dataOut_payload_0_403 ? _zz_dataOut_payload_0_401 : _zz_dataOut_payload_0_398);
    _zz_dataOut_payload_0_407 <= (_zz_dataOut_payload_0_403 ? _zz_dataOut_payload_0_398 : _zz_dataOut_payload_0_401);
    _zz_dataOut_payload_0_416 <= (_zz_dataOut_payload_0_414 ? _zz_dataOut_payload_0_409 : _zz_dataOut_payload_0_412);
    _zz_dataOut_payload_0_417 <= (_zz_dataOut_payload_0_414 ? _zz_dataOut_payload_0_412 : _zz_dataOut_payload_0_409);
    _zz_dataOut_payload_0_418 <= (_zz_dataOut_payload_0_415 ? _zz_dataOut_payload_0_413 : _zz_dataOut_payload_0_410);
    _zz_dataOut_payload_0_419 <= (_zz_dataOut_payload_0_415 ? _zz_dataOut_payload_0_410 : _zz_dataOut_payload_0_413);
    _zz_dataOut_payload_0_428 <= (_zz_dataOut_payload_0_426 ? _zz_dataOut_payload_0_421 : _zz_dataOut_payload_0_424);
    _zz_dataOut_payload_0_429 <= (_zz_dataOut_payload_0_426 ? _zz_dataOut_payload_0_424 : _zz_dataOut_payload_0_421);
    _zz_dataOut_payload_0_430 <= (_zz_dataOut_payload_0_427 ? _zz_dataOut_payload_0_425 : _zz_dataOut_payload_0_422);
    _zz_dataOut_payload_0_431 <= (_zz_dataOut_payload_0_427 ? _zz_dataOut_payload_0_422 : _zz_dataOut_payload_0_425);
    _zz_dataOut_payload_0_440 <= (_zz_dataOut_payload_0_438 ? _zz_dataOut_payload_0_433 : _zz_dataOut_payload_0_436);
    _zz_dataOut_payload_0_441 <= (_zz_dataOut_payload_0_438 ? _zz_dataOut_payload_0_436 : _zz_dataOut_payload_0_433);
    _zz_dataOut_payload_0_442 <= (_zz_dataOut_payload_0_439 ? _zz_dataOut_payload_0_437 : _zz_dataOut_payload_0_434);
    _zz_dataOut_payload_0_443 <= (_zz_dataOut_payload_0_439 ? _zz_dataOut_payload_0_434 : _zz_dataOut_payload_0_437);
    _zz_dataOut_payload_0_452 <= (_zz_dataOut_payload_0_450 ? _zz_dataOut_payload_0_445 : _zz_dataOut_payload_0_448);
    _zz_dataOut_payload_0_453 <= (_zz_dataOut_payload_0_450 ? _zz_dataOut_payload_0_448 : _zz_dataOut_payload_0_445);
    _zz_dataOut_payload_0_454 <= (_zz_dataOut_payload_0_451 ? _zz_dataOut_payload_0_449 : _zz_dataOut_payload_0_446);
    _zz_dataOut_payload_0_455 <= (_zz_dataOut_payload_0_451 ? _zz_dataOut_payload_0_446 : _zz_dataOut_payload_0_449);
    _zz_dataOut_payload_0_464 <= (_zz_dataOut_payload_0_462 ? _zz_dataOut_payload_0_457 : _zz_dataOut_payload_0_460);
    _zz_dataOut_payload_0_465 <= (_zz_dataOut_payload_0_462 ? _zz_dataOut_payload_0_460 : _zz_dataOut_payload_0_457);
    _zz_dataOut_payload_0_466 <= (_zz_dataOut_payload_0_463 ? _zz_dataOut_payload_0_461 : _zz_dataOut_payload_0_458);
    _zz_dataOut_payload_0_467 <= (_zz_dataOut_payload_0_463 ? _zz_dataOut_payload_0_458 : _zz_dataOut_payload_0_461);
    _zz_dataOut_payload_0_476 <= (_zz_dataOut_payload_0_474 ? _zz_dataOut_payload_0_469 : _zz_dataOut_payload_0_472);
    _zz_dataOut_payload_0_477 <= (_zz_dataOut_payload_0_474 ? _zz_dataOut_payload_0_472 : _zz_dataOut_payload_0_469);
    _zz_dataOut_payload_0_478 <= (_zz_dataOut_payload_0_475 ? _zz_dataOut_payload_0_473 : _zz_dataOut_payload_0_470);
    _zz_dataOut_payload_0_479 <= (_zz_dataOut_payload_0_475 ? _zz_dataOut_payload_0_470 : _zz_dataOut_payload_0_473);
    _zz_dataOut_payload_0_488 <= (_zz_dataOut_payload_0_486 ? _zz_dataOut_payload_0_481 : _zz_dataOut_payload_0_484);
    _zz_dataOut_payload_0_489 <= (_zz_dataOut_payload_0_486 ? _zz_dataOut_payload_0_484 : _zz_dataOut_payload_0_481);
    _zz_dataOut_payload_0_490 <= (_zz_dataOut_payload_0_487 ? _zz_dataOut_payload_0_485 : _zz_dataOut_payload_0_482);
    _zz_dataOut_payload_0_491 <= (_zz_dataOut_payload_0_487 ? _zz_dataOut_payload_0_482 : _zz_dataOut_payload_0_485);
    _zz_dataOut_payload_0_500 <= (_zz_dataOut_payload_0_498 ? _zz_dataOut_payload_0_493 : _zz_dataOut_payload_0_496);
    _zz_dataOut_payload_0_501 <= (_zz_dataOut_payload_0_498 ? _zz_dataOut_payload_0_496 : _zz_dataOut_payload_0_493);
    _zz_dataOut_payload_0_502 <= (_zz_dataOut_payload_0_499 ? _zz_dataOut_payload_0_497 : _zz_dataOut_payload_0_494);
    _zz_dataOut_payload_0_503 <= (_zz_dataOut_payload_0_499 ? _zz_dataOut_payload_0_494 : _zz_dataOut_payload_0_497);
    _zz_dataOut_payload_0_512 <= (_zz_dataOut_payload_0_510 ? _zz_dataOut_payload_0_505 : _zz_dataOut_payload_0_508);
    _zz_dataOut_payload_0_513 <= (_zz_dataOut_payload_0_510 ? _zz_dataOut_payload_0_508 : _zz_dataOut_payload_0_505);
    _zz_dataOut_payload_0_514 <= (_zz_dataOut_payload_0_511 ? _zz_dataOut_payload_0_509 : _zz_dataOut_payload_0_506);
    _zz_dataOut_payload_0_515 <= (_zz_dataOut_payload_0_511 ? _zz_dataOut_payload_0_506 : _zz_dataOut_payload_0_509);
    _zz_dataOut_payload_0_524 <= (_zz_dataOut_payload_0_522 ? _zz_dataOut_payload_0_517 : _zz_dataOut_payload_0_520);
    _zz_dataOut_payload_0_525 <= (_zz_dataOut_payload_0_522 ? _zz_dataOut_payload_0_520 : _zz_dataOut_payload_0_517);
    _zz_dataOut_payload_0_526 <= (_zz_dataOut_payload_0_523 ? _zz_dataOut_payload_0_521 : _zz_dataOut_payload_0_518);
    _zz_dataOut_payload_0_527 <= (_zz_dataOut_payload_0_523 ? _zz_dataOut_payload_0_518 : _zz_dataOut_payload_0_521);
    _zz_dataOut_payload_0_536 <= (_zz_dataOut_payload_0_534 ? _zz_dataOut_payload_0_529 : _zz_dataOut_payload_0_532);
    _zz_dataOut_payload_0_537 <= (_zz_dataOut_payload_0_534 ? _zz_dataOut_payload_0_532 : _zz_dataOut_payload_0_529);
    _zz_dataOut_payload_0_538 <= (_zz_dataOut_payload_0_535 ? _zz_dataOut_payload_0_533 : _zz_dataOut_payload_0_530);
    _zz_dataOut_payload_0_539 <= (_zz_dataOut_payload_0_535 ? _zz_dataOut_payload_0_530 : _zz_dataOut_payload_0_533);
    _zz_dataOut_payload_0_548 <= (_zz_dataOut_payload_0_546 ? _zz_dataOut_payload_0_541 : _zz_dataOut_payload_0_544);
    _zz_dataOut_payload_0_549 <= (_zz_dataOut_payload_0_546 ? _zz_dataOut_payload_0_544 : _zz_dataOut_payload_0_541);
    _zz_dataOut_payload_0_550 <= (_zz_dataOut_payload_0_547 ? _zz_dataOut_payload_0_545 : _zz_dataOut_payload_0_542);
    _zz_dataOut_payload_0_551 <= (_zz_dataOut_payload_0_547 ? _zz_dataOut_payload_0_542 : _zz_dataOut_payload_0_545);
    _zz_dataOut_payload_0_560 <= (_zz_dataOut_payload_0_558 ? _zz_dataOut_payload_0_553 : _zz_dataOut_payload_0_556);
    _zz_dataOut_payload_0_561 <= (_zz_dataOut_payload_0_558 ? _zz_dataOut_payload_0_556 : _zz_dataOut_payload_0_553);
    _zz_dataOut_payload_0_562 <= (_zz_dataOut_payload_0_559 ? _zz_dataOut_payload_0_557 : _zz_dataOut_payload_0_554);
    _zz_dataOut_payload_0_563 <= (_zz_dataOut_payload_0_559 ? _zz_dataOut_payload_0_554 : _zz_dataOut_payload_0_557);
    _zz_dataOut_payload_0_572 <= (_zz_dataOut_payload_0_570 ? _zz_dataOut_payload_0_565 : _zz_dataOut_payload_0_568);
    _zz_dataOut_payload_0_573 <= (_zz_dataOut_payload_0_570 ? _zz_dataOut_payload_0_568 : _zz_dataOut_payload_0_565);
    _zz_dataOut_payload_0_574 <= (_zz_dataOut_payload_0_571 ? _zz_dataOut_payload_0_569 : _zz_dataOut_payload_0_566);
    _zz_dataOut_payload_0_575 <= (_zz_dataOut_payload_0_571 ? _zz_dataOut_payload_0_566 : _zz_dataOut_payload_0_569);
    _zz_dataOut_payload_0_584 <= (_zz_dataOut_payload_0_582 ? _zz_dataOut_payload_0_577 : _zz_dataOut_payload_0_580);
    _zz_dataOut_payload_0_585 <= (_zz_dataOut_payload_0_582 ? _zz_dataOut_payload_0_580 : _zz_dataOut_payload_0_577);
    _zz_dataOut_payload_0_586 <= (_zz_dataOut_payload_0_583 ? _zz_dataOut_payload_0_581 : _zz_dataOut_payload_0_578);
    _zz_dataOut_payload_0_587 <= (_zz_dataOut_payload_0_583 ? _zz_dataOut_payload_0_578 : _zz_dataOut_payload_0_581);
    _zz_dataOut_payload_0_596 <= (_zz_dataOut_payload_0_594 ? _zz_dataOut_payload_0_589 : _zz_dataOut_payload_0_592);
    _zz_dataOut_payload_0_597 <= (_zz_dataOut_payload_0_594 ? _zz_dataOut_payload_0_592 : _zz_dataOut_payload_0_589);
    _zz_dataOut_payload_0_598 <= (_zz_dataOut_payload_0_595 ? _zz_dataOut_payload_0_593 : _zz_dataOut_payload_0_590);
    _zz_dataOut_payload_0_599 <= (_zz_dataOut_payload_0_595 ? _zz_dataOut_payload_0_590 : _zz_dataOut_payload_0_593);
    _zz_dataOut_payload_0_608 <= (_zz_dataOut_payload_0_606 ? _zz_dataOut_payload_0_601 : _zz_dataOut_payload_0_604);
    _zz_dataOut_payload_0_609 <= (_zz_dataOut_payload_0_606 ? _zz_dataOut_payload_0_604 : _zz_dataOut_payload_0_601);
    _zz_dataOut_payload_0_610 <= (_zz_dataOut_payload_0_607 ? _zz_dataOut_payload_0_605 : _zz_dataOut_payload_0_602);
    _zz_dataOut_payload_0_611 <= (_zz_dataOut_payload_0_607 ? _zz_dataOut_payload_0_602 : _zz_dataOut_payload_0_605);
    _zz_dataOut_payload_0_620 <= (_zz_dataOut_payload_0_618 ? _zz_dataOut_payload_0_613 : _zz_dataOut_payload_0_616);
    _zz_dataOut_payload_0_621 <= (_zz_dataOut_payload_0_618 ? _zz_dataOut_payload_0_616 : _zz_dataOut_payload_0_613);
    _zz_dataOut_payload_0_622 <= (_zz_dataOut_payload_0_619 ? _zz_dataOut_payload_0_617 : _zz_dataOut_payload_0_614);
    _zz_dataOut_payload_0_623 <= (_zz_dataOut_payload_0_619 ? _zz_dataOut_payload_0_614 : _zz_dataOut_payload_0_617);
    _zz_dataOut_payload_0_632 <= (_zz_dataOut_payload_0_630 ? _zz_dataOut_payload_0_625 : _zz_dataOut_payload_0_628);
    _zz_dataOut_payload_0_633 <= (_zz_dataOut_payload_0_630 ? _zz_dataOut_payload_0_628 : _zz_dataOut_payload_0_625);
    _zz_dataOut_payload_0_634 <= (_zz_dataOut_payload_0_631 ? _zz_dataOut_payload_0_629 : _zz_dataOut_payload_0_626);
    _zz_dataOut_payload_0_635 <= (_zz_dataOut_payload_0_631 ? _zz_dataOut_payload_0_626 : _zz_dataOut_payload_0_629);
    _zz_dataOut_payload_0_644 <= (_zz_dataOut_payload_0_642 ? _zz_dataOut_payload_0_637 : _zz_dataOut_payload_0_640);
    _zz_dataOut_payload_0_645 <= (_zz_dataOut_payload_0_642 ? _zz_dataOut_payload_0_640 : _zz_dataOut_payload_0_637);
    _zz_dataOut_payload_0_646 <= (_zz_dataOut_payload_0_643 ? _zz_dataOut_payload_0_641 : _zz_dataOut_payload_0_638);
    _zz_dataOut_payload_0_647 <= (_zz_dataOut_payload_0_643 ? _zz_dataOut_payload_0_638 : _zz_dataOut_payload_0_641);
    _zz_dataOut_payload_0_656 <= (_zz_dataOut_payload_0_654 ? _zz_dataOut_payload_0_649 : _zz_dataOut_payload_0_652);
    _zz_dataOut_payload_0_657 <= (_zz_dataOut_payload_0_654 ? _zz_dataOut_payload_0_652 : _zz_dataOut_payload_0_649);
    _zz_dataOut_payload_0_658 <= (_zz_dataOut_payload_0_655 ? _zz_dataOut_payload_0_653 : _zz_dataOut_payload_0_650);
    _zz_dataOut_payload_0_659 <= (_zz_dataOut_payload_0_655 ? _zz_dataOut_payload_0_650 : _zz_dataOut_payload_0_653);
    _zz_dataOut_payload_0_668 <= (_zz_dataOut_payload_0_666 ? _zz_dataOut_payload_0_661 : _zz_dataOut_payload_0_664);
    _zz_dataOut_payload_0_669 <= (_zz_dataOut_payload_0_666 ? _zz_dataOut_payload_0_664 : _zz_dataOut_payload_0_661);
    _zz_dataOut_payload_0_670 <= (_zz_dataOut_payload_0_667 ? _zz_dataOut_payload_0_665 : _zz_dataOut_payload_0_662);
    _zz_dataOut_payload_0_671 <= (_zz_dataOut_payload_0_667 ? _zz_dataOut_payload_0_662 : _zz_dataOut_payload_0_665);
    _zz_dataOut_payload_0_680 <= (_zz_dataOut_payload_0_678 ? _zz_dataOut_payload_0_673 : _zz_dataOut_payload_0_676);
    _zz_dataOut_payload_0_681 <= (_zz_dataOut_payload_0_678 ? _zz_dataOut_payload_0_676 : _zz_dataOut_payload_0_673);
    _zz_dataOut_payload_0_682 <= (_zz_dataOut_payload_0_679 ? _zz_dataOut_payload_0_677 : _zz_dataOut_payload_0_674);
    _zz_dataOut_payload_0_683 <= (_zz_dataOut_payload_0_679 ? _zz_dataOut_payload_0_674 : _zz_dataOut_payload_0_677);
    _zz_dataOut_payload_0_692 <= (_zz_dataOut_payload_0_690 ? _zz_dataOut_payload_0_685 : _zz_dataOut_payload_0_688);
    _zz_dataOut_payload_0_693 <= (_zz_dataOut_payload_0_690 ? _zz_dataOut_payload_0_688 : _zz_dataOut_payload_0_685);
    _zz_dataOut_payload_0_694 <= (_zz_dataOut_payload_0_691 ? _zz_dataOut_payload_0_689 : _zz_dataOut_payload_0_686);
    _zz_dataOut_payload_0_695 <= (_zz_dataOut_payload_0_691 ? _zz_dataOut_payload_0_686 : _zz_dataOut_payload_0_689);
    _zz_dataOut_payload_0_704 <= (_zz_dataOut_payload_0_702 ? _zz_dataOut_payload_0_697 : _zz_dataOut_payload_0_700);
    _zz_dataOut_payload_0_705 <= (_zz_dataOut_payload_0_702 ? _zz_dataOut_payload_0_700 : _zz_dataOut_payload_0_697);
    _zz_dataOut_payload_0_706 <= (_zz_dataOut_payload_0_703 ? _zz_dataOut_payload_0_701 : _zz_dataOut_payload_0_698);
    _zz_dataOut_payload_0_707 <= (_zz_dataOut_payload_0_703 ? _zz_dataOut_payload_0_698 : _zz_dataOut_payload_0_701);
    _zz_dataOut_payload_0_716 <= (_zz_dataOut_payload_0_714 ? _zz_dataOut_payload_0_709 : _zz_dataOut_payload_0_712);
    _zz_dataOut_payload_0_717 <= (_zz_dataOut_payload_0_714 ? _zz_dataOut_payload_0_712 : _zz_dataOut_payload_0_709);
    _zz_dataOut_payload_0_718 <= (_zz_dataOut_payload_0_715 ? _zz_dataOut_payload_0_713 : _zz_dataOut_payload_0_710);
    _zz_dataOut_payload_0_719 <= (_zz_dataOut_payload_0_715 ? _zz_dataOut_payload_0_710 : _zz_dataOut_payload_0_713);
    _zz_dataOut_payload_0_728 <= (_zz_dataOut_payload_0_726 ? _zz_dataOut_payload_0_721 : _zz_dataOut_payload_0_724);
    _zz_dataOut_payload_0_729 <= (_zz_dataOut_payload_0_726 ? _zz_dataOut_payload_0_724 : _zz_dataOut_payload_0_721);
    _zz_dataOut_payload_0_730 <= (_zz_dataOut_payload_0_727 ? _zz_dataOut_payload_0_725 : _zz_dataOut_payload_0_722);
    _zz_dataOut_payload_0_731 <= (_zz_dataOut_payload_0_727 ? _zz_dataOut_payload_0_722 : _zz_dataOut_payload_0_725);
    _zz_dataOut_payload_0_740 <= (_zz_dataOut_payload_0_738 ? _zz_dataOut_payload_0_733 : _zz_dataOut_payload_0_736);
    _zz_dataOut_payload_0_741 <= (_zz_dataOut_payload_0_738 ? _zz_dataOut_payload_0_736 : _zz_dataOut_payload_0_733);
    _zz_dataOut_payload_0_742 <= (_zz_dataOut_payload_0_739 ? _zz_dataOut_payload_0_737 : _zz_dataOut_payload_0_734);
    _zz_dataOut_payload_0_743 <= (_zz_dataOut_payload_0_739 ? _zz_dataOut_payload_0_734 : _zz_dataOut_payload_0_737);
    _zz_dataOut_payload_0_752 <= (_zz_dataOut_payload_0_750 ? _zz_dataOut_payload_0_745 : _zz_dataOut_payload_0_748);
    _zz_dataOut_payload_0_753 <= (_zz_dataOut_payload_0_750 ? _zz_dataOut_payload_0_748 : _zz_dataOut_payload_0_745);
    _zz_dataOut_payload_0_754 <= (_zz_dataOut_payload_0_751 ? _zz_dataOut_payload_0_749 : _zz_dataOut_payload_0_746);
    _zz_dataOut_payload_0_755 <= (_zz_dataOut_payload_0_751 ? _zz_dataOut_payload_0_746 : _zz_dataOut_payload_0_749);
    _zz_dataOut_payload_0_764 <= (_zz_dataOut_payload_0_762 ? _zz_dataOut_payload_0_757 : _zz_dataOut_payload_0_760);
    _zz_dataOut_payload_0_765 <= (_zz_dataOut_payload_0_762 ? _zz_dataOut_payload_0_760 : _zz_dataOut_payload_0_757);
    _zz_dataOut_payload_0_766 <= (_zz_dataOut_payload_0_763 ? _zz_dataOut_payload_0_761 : _zz_dataOut_payload_0_758);
    _zz_dataOut_payload_0_767 <= (_zz_dataOut_payload_0_763 ? _zz_dataOut_payload_0_758 : _zz_dataOut_payload_0_761);
    _zz_dataOut_payload_0_776 <= (_zz_dataOut_payload_0_774 ? _zz_dataOut_payload_0_769 : _zz_dataOut_payload_0_772);
    _zz_dataOut_payload_0_777 <= (_zz_dataOut_payload_0_774 ? _zz_dataOut_payload_0_772 : _zz_dataOut_payload_0_769);
    _zz_dataOut_payload_0_778 <= (_zz_dataOut_payload_0_775 ? _zz_dataOut_payload_0_773 : _zz_dataOut_payload_0_770);
    _zz_dataOut_payload_0_779 <= (_zz_dataOut_payload_0_775 ? _zz_dataOut_payload_0_770 : _zz_dataOut_payload_0_773);
    _zz_dataOut_payload_0_788 <= (_zz_dataOut_payload_0_786 ? _zz_dataOut_payload_0_781 : _zz_dataOut_payload_0_784);
    _zz_dataOut_payload_0_789 <= (_zz_dataOut_payload_0_786 ? _zz_dataOut_payload_0_784 : _zz_dataOut_payload_0_781);
    _zz_dataOut_payload_0_790 <= (_zz_dataOut_payload_0_787 ? _zz_dataOut_payload_0_785 : _zz_dataOut_payload_0_782);
    _zz_dataOut_payload_0_791 <= (_zz_dataOut_payload_0_787 ? _zz_dataOut_payload_0_782 : _zz_dataOut_payload_0_785);
    _zz_dataOut_payload_0_800 <= (_zz_dataOut_payload_0_798 ? _zz_dataOut_payload_0_793 : _zz_dataOut_payload_0_796);
    _zz_dataOut_payload_0_801 <= (_zz_dataOut_payload_0_798 ? _zz_dataOut_payload_0_796 : _zz_dataOut_payload_0_793);
    _zz_dataOut_payload_0_802 <= (_zz_dataOut_payload_0_799 ? _zz_dataOut_payload_0_797 : _zz_dataOut_payload_0_794);
    _zz_dataOut_payload_0_803 <= (_zz_dataOut_payload_0_799 ? _zz_dataOut_payload_0_794 : _zz_dataOut_payload_0_797);
    _zz_dataOut_payload_0_812 <= (_zz_dataOut_payload_0_810 ? _zz_dataOut_payload_0_805 : _zz_dataOut_payload_0_808);
    _zz_dataOut_payload_0_813 <= (_zz_dataOut_payload_0_810 ? _zz_dataOut_payload_0_808 : _zz_dataOut_payload_0_805);
    _zz_dataOut_payload_0_814 <= (_zz_dataOut_payload_0_811 ? _zz_dataOut_payload_0_809 : _zz_dataOut_payload_0_806);
    _zz_dataOut_payload_0_815 <= (_zz_dataOut_payload_0_811 ? _zz_dataOut_payload_0_806 : _zz_dataOut_payload_0_809);
    _zz_dataOut_payload_0_824 <= (_zz_dataOut_payload_0_822 ? _zz_dataOut_payload_0_817 : _zz_dataOut_payload_0_820);
    _zz_dataOut_payload_0_825 <= (_zz_dataOut_payload_0_822 ? _zz_dataOut_payload_0_820 : _zz_dataOut_payload_0_817);
    _zz_dataOut_payload_0_826 <= (_zz_dataOut_payload_0_823 ? _zz_dataOut_payload_0_821 : _zz_dataOut_payload_0_818);
    _zz_dataOut_payload_0_827 <= (_zz_dataOut_payload_0_823 ? _zz_dataOut_payload_0_818 : _zz_dataOut_payload_0_821);
    _zz_dataOut_payload_0_836 <= (_zz_dataOut_payload_0_834 ? _zz_dataOut_payload_0_829 : _zz_dataOut_payload_0_832);
    _zz_dataOut_payload_0_837 <= (_zz_dataOut_payload_0_834 ? _zz_dataOut_payload_0_832 : _zz_dataOut_payload_0_829);
    _zz_dataOut_payload_0_838 <= (_zz_dataOut_payload_0_835 ? _zz_dataOut_payload_0_833 : _zz_dataOut_payload_0_830);
    _zz_dataOut_payload_0_839 <= (_zz_dataOut_payload_0_835 ? _zz_dataOut_payload_0_830 : _zz_dataOut_payload_0_833);
    _zz_dataOut_payload_0_848 <= (_zz_dataOut_payload_0_846 ? _zz_dataOut_payload_0_841 : _zz_dataOut_payload_0_844);
    _zz_dataOut_payload_0_849 <= (_zz_dataOut_payload_0_846 ? _zz_dataOut_payload_0_844 : _zz_dataOut_payload_0_841);
    _zz_dataOut_payload_0_850 <= (_zz_dataOut_payload_0_847 ? _zz_dataOut_payload_0_845 : _zz_dataOut_payload_0_842);
    _zz_dataOut_payload_0_851 <= (_zz_dataOut_payload_0_847 ? _zz_dataOut_payload_0_842 : _zz_dataOut_payload_0_845);
    _zz_dataOut_payload_0_860 <= (_zz_dataOut_payload_0_858 ? _zz_dataOut_payload_0_853 : _zz_dataOut_payload_0_856);
    _zz_dataOut_payload_0_861 <= (_zz_dataOut_payload_0_858 ? _zz_dataOut_payload_0_856 : _zz_dataOut_payload_0_853);
    _zz_dataOut_payload_0_862 <= (_zz_dataOut_payload_0_859 ? _zz_dataOut_payload_0_857 : _zz_dataOut_payload_0_854);
    _zz_dataOut_payload_0_863 <= (_zz_dataOut_payload_0_859 ? _zz_dataOut_payload_0_854 : _zz_dataOut_payload_0_857);
    _zz_dataOut_payload_0_872 <= (_zz_dataOut_payload_0_870 ? _zz_dataOut_payload_0_865 : _zz_dataOut_payload_0_868);
    _zz_dataOut_payload_0_873 <= (_zz_dataOut_payload_0_870 ? _zz_dataOut_payload_0_868 : _zz_dataOut_payload_0_865);
    _zz_dataOut_payload_0_874 <= (_zz_dataOut_payload_0_871 ? _zz_dataOut_payload_0_869 : _zz_dataOut_payload_0_866);
    _zz_dataOut_payload_0_875 <= (_zz_dataOut_payload_0_871 ? _zz_dataOut_payload_0_866 : _zz_dataOut_payload_0_869);
    _zz_dataOut_payload_0_884 <= (_zz_dataOut_payload_0_882 ? _zz_dataOut_payload_0_877 : _zz_dataOut_payload_0_880);
    _zz_dataOut_payload_0_885 <= (_zz_dataOut_payload_0_882 ? _zz_dataOut_payload_0_880 : _zz_dataOut_payload_0_877);
    _zz_dataOut_payload_0_886 <= (_zz_dataOut_payload_0_883 ? _zz_dataOut_payload_0_881 : _zz_dataOut_payload_0_878);
    _zz_dataOut_payload_0_887 <= (_zz_dataOut_payload_0_883 ? _zz_dataOut_payload_0_878 : _zz_dataOut_payload_0_881);
    _zz_dataOut_payload_0_896 <= (_zz_dataOut_payload_0_894 ? _zz_dataOut_payload_0_889 : _zz_dataOut_payload_0_892);
    _zz_dataOut_payload_0_897 <= (_zz_dataOut_payload_0_894 ? _zz_dataOut_payload_0_892 : _zz_dataOut_payload_0_889);
    _zz_dataOut_payload_0_898 <= (_zz_dataOut_payload_0_895 ? _zz_dataOut_payload_0_893 : _zz_dataOut_payload_0_890);
    _zz_dataOut_payload_0_899 <= (_zz_dataOut_payload_0_895 ? _zz_dataOut_payload_0_890 : _zz_dataOut_payload_0_893);
    _zz_dataOut_payload_0_908 <= (_zz_dataOut_payload_0_906 ? _zz_dataOut_payload_0_901 : _zz_dataOut_payload_0_904);
    _zz_dataOut_payload_0_909 <= (_zz_dataOut_payload_0_906 ? _zz_dataOut_payload_0_904 : _zz_dataOut_payload_0_901);
    _zz_dataOut_payload_0_910 <= (_zz_dataOut_payload_0_907 ? _zz_dataOut_payload_0_905 : _zz_dataOut_payload_0_902);
    _zz_dataOut_payload_0_911 <= (_zz_dataOut_payload_0_907 ? _zz_dataOut_payload_0_902 : _zz_dataOut_payload_0_905);
    _zz_dataOut_payload_0_920 <= (_zz_dataOut_payload_0_918 ? _zz_dataOut_payload_0_913 : _zz_dataOut_payload_0_916);
    _zz_dataOut_payload_0_921 <= (_zz_dataOut_payload_0_918 ? _zz_dataOut_payload_0_916 : _zz_dataOut_payload_0_913);
    _zz_dataOut_payload_0_922 <= (_zz_dataOut_payload_0_919 ? _zz_dataOut_payload_0_917 : _zz_dataOut_payload_0_914);
    _zz_dataOut_payload_0_923 <= (_zz_dataOut_payload_0_919 ? _zz_dataOut_payload_0_914 : _zz_dataOut_payload_0_917);
    _zz_dataOut_payload_0_932 <= (_zz_dataOut_payload_0_930 ? _zz_dataOut_payload_0_925 : _zz_dataOut_payload_0_928);
    _zz_dataOut_payload_0_933 <= (_zz_dataOut_payload_0_930 ? _zz_dataOut_payload_0_928 : _zz_dataOut_payload_0_925);
    _zz_dataOut_payload_0_934 <= (_zz_dataOut_payload_0_931 ? _zz_dataOut_payload_0_929 : _zz_dataOut_payload_0_926);
    _zz_dataOut_payload_0_935 <= (_zz_dataOut_payload_0_931 ? _zz_dataOut_payload_0_926 : _zz_dataOut_payload_0_929);
    _zz_dataOut_payload_0_944 <= (_zz_dataOut_payload_0_942 ? _zz_dataOut_payload_0_937 : _zz_dataOut_payload_0_940);
    _zz_dataOut_payload_0_945 <= (_zz_dataOut_payload_0_942 ? _zz_dataOut_payload_0_940 : _zz_dataOut_payload_0_937);
    _zz_dataOut_payload_0_946 <= (_zz_dataOut_payload_0_943 ? _zz_dataOut_payload_0_941 : _zz_dataOut_payload_0_938);
    _zz_dataOut_payload_0_947 <= (_zz_dataOut_payload_0_943 ? _zz_dataOut_payload_0_938 : _zz_dataOut_payload_0_941);
    _zz_dataOut_payload_0_956 <= (_zz_dataOut_payload_0_954 ? _zz_dataOut_payload_0_949 : _zz_dataOut_payload_0_952);
    _zz_dataOut_payload_0_957 <= (_zz_dataOut_payload_0_954 ? _zz_dataOut_payload_0_952 : _zz_dataOut_payload_0_949);
    _zz_dataOut_payload_0_958 <= (_zz_dataOut_payload_0_955 ? _zz_dataOut_payload_0_953 : _zz_dataOut_payload_0_950);
    _zz_dataOut_payload_0_959 <= (_zz_dataOut_payload_0_955 ? _zz_dataOut_payload_0_950 : _zz_dataOut_payload_0_953);
    _zz_dataOut_payload_0_968 <= (_zz_dataOut_payload_0_966 ? _zz_dataOut_payload_0_961 : _zz_dataOut_payload_0_964);
    _zz_dataOut_payload_0_969 <= (_zz_dataOut_payload_0_966 ? _zz_dataOut_payload_0_964 : _zz_dataOut_payload_0_961);
    _zz_dataOut_payload_0_970 <= (_zz_dataOut_payload_0_967 ? _zz_dataOut_payload_0_965 : _zz_dataOut_payload_0_962);
    _zz_dataOut_payload_0_971 <= (_zz_dataOut_payload_0_967 ? _zz_dataOut_payload_0_962 : _zz_dataOut_payload_0_965);
    _zz_dataOut_payload_0_980 <= (_zz_dataOut_payload_0_978 ? _zz_dataOut_payload_0_973 : _zz_dataOut_payload_0_976);
    _zz_dataOut_payload_0_981 <= (_zz_dataOut_payload_0_978 ? _zz_dataOut_payload_0_976 : _zz_dataOut_payload_0_973);
    _zz_dataOut_payload_0_982 <= (_zz_dataOut_payload_0_979 ? _zz_dataOut_payload_0_977 : _zz_dataOut_payload_0_974);
    _zz_dataOut_payload_0_983 <= (_zz_dataOut_payload_0_979 ? _zz_dataOut_payload_0_974 : _zz_dataOut_payload_0_977);
    _zz_dataOut_payload_0_992 <= (_zz_dataOut_payload_0_990 ? _zz_dataOut_payload_0_985 : _zz_dataOut_payload_0_988);
    _zz_dataOut_payload_0_993 <= (_zz_dataOut_payload_0_990 ? _zz_dataOut_payload_0_988 : _zz_dataOut_payload_0_985);
    _zz_dataOut_payload_0_994 <= (_zz_dataOut_payload_0_991 ? _zz_dataOut_payload_0_989 : _zz_dataOut_payload_0_986);
    _zz_dataOut_payload_0_995 <= (_zz_dataOut_payload_0_991 ? _zz_dataOut_payload_0_986 : _zz_dataOut_payload_0_989);
    _zz_dataOut_payload_0_1004 <= (_zz_dataOut_payload_0_1002 ? _zz_dataOut_payload_0_997 : _zz_dataOut_payload_0_1000);
    _zz_dataOut_payload_0_1005 <= (_zz_dataOut_payload_0_1002 ? _zz_dataOut_payload_0_1000 : _zz_dataOut_payload_0_997);
    _zz_dataOut_payload_0_1006 <= (_zz_dataOut_payload_0_1003 ? _zz_dataOut_payload_0_1001 : _zz_dataOut_payload_0_998);
    _zz_dataOut_payload_0_1007 <= (_zz_dataOut_payload_0_1003 ? _zz_dataOut_payload_0_998 : _zz_dataOut_payload_0_1001);
    _zz_dataOut_payload_0_1016 <= (_zz_dataOut_payload_0_1014 ? _zz_dataOut_payload_0_1009 : _zz_dataOut_payload_0_1012);
    _zz_dataOut_payload_0_1017 <= (_zz_dataOut_payload_0_1014 ? _zz_dataOut_payload_0_1012 : _zz_dataOut_payload_0_1009);
    _zz_dataOut_payload_0_1018 <= (_zz_dataOut_payload_0_1015 ? _zz_dataOut_payload_0_1013 : _zz_dataOut_payload_0_1010);
    _zz_dataOut_payload_0_1019 <= (_zz_dataOut_payload_0_1015 ? _zz_dataOut_payload_0_1010 : _zz_dataOut_payload_0_1013);
    _zz_dataOut_payload_0_1028 <= (_zz_dataOut_payload_0_1026 ? _zz_dataOut_payload_0_1021 : _zz_dataOut_payload_0_1024);
    _zz_dataOut_payload_0_1029 <= (_zz_dataOut_payload_0_1026 ? _zz_dataOut_payload_0_1024 : _zz_dataOut_payload_0_1021);
    _zz_dataOut_payload_0_1030 <= (_zz_dataOut_payload_0_1027 ? _zz_dataOut_payload_0_1025 : _zz_dataOut_payload_0_1022);
    _zz_dataOut_payload_0_1031 <= (_zz_dataOut_payload_0_1027 ? _zz_dataOut_payload_0_1022 : _zz_dataOut_payload_0_1025);
    _zz_dataOut_payload_0_1040 <= (_zz_dataOut_payload_0_1038 ? _zz_dataOut_payload_0_1033 : _zz_dataOut_payload_0_1036);
    _zz_dataOut_payload_0_1041 <= (_zz_dataOut_payload_0_1038 ? _zz_dataOut_payload_0_1036 : _zz_dataOut_payload_0_1033);
    _zz_dataOut_payload_0_1042 <= (_zz_dataOut_payload_0_1039 ? _zz_dataOut_payload_0_1037 : _zz_dataOut_payload_0_1034);
    _zz_dataOut_payload_0_1043 <= (_zz_dataOut_payload_0_1039 ? _zz_dataOut_payload_0_1034 : _zz_dataOut_payload_0_1037);
    _zz_dataOut_payload_0_1052 <= (_zz_dataOut_payload_0_1050 ? _zz_dataOut_payload_0_1045 : _zz_dataOut_payload_0_1048);
    _zz_dataOut_payload_0_1053 <= (_zz_dataOut_payload_0_1050 ? _zz_dataOut_payload_0_1048 : _zz_dataOut_payload_0_1045);
    _zz_dataOut_payload_0_1054 <= (_zz_dataOut_payload_0_1051 ? _zz_dataOut_payload_0_1049 : _zz_dataOut_payload_0_1046);
    _zz_dataOut_payload_0_1055 <= (_zz_dataOut_payload_0_1051 ? _zz_dataOut_payload_0_1046 : _zz_dataOut_payload_0_1049);
    _zz_dataOut_payload_0_1064 <= (_zz_dataOut_payload_0_1062 ? _zz_dataOut_payload_0_1057 : _zz_dataOut_payload_0_1060);
    _zz_dataOut_payload_0_1065 <= (_zz_dataOut_payload_0_1062 ? _zz_dataOut_payload_0_1060 : _zz_dataOut_payload_0_1057);
    _zz_dataOut_payload_0_1066 <= (_zz_dataOut_payload_0_1063 ? _zz_dataOut_payload_0_1061 : _zz_dataOut_payload_0_1058);
    _zz_dataOut_payload_0_1067 <= (_zz_dataOut_payload_0_1063 ? _zz_dataOut_payload_0_1058 : _zz_dataOut_payload_0_1061);
    _zz_dataOut_payload_0_1076 <= (_zz_dataOut_payload_0_1074 ? _zz_dataOut_payload_0_1069 : _zz_dataOut_payload_0_1072);
    _zz_dataOut_payload_0_1077 <= (_zz_dataOut_payload_0_1074 ? _zz_dataOut_payload_0_1072 : _zz_dataOut_payload_0_1069);
    _zz_dataOut_payload_0_1078 <= (_zz_dataOut_payload_0_1075 ? _zz_dataOut_payload_0_1073 : _zz_dataOut_payload_0_1070);
    _zz_dataOut_payload_0_1079 <= (_zz_dataOut_payload_0_1075 ? _zz_dataOut_payload_0_1070 : _zz_dataOut_payload_0_1073);
    _zz_dataOut_payload_0_1088 <= (_zz_dataOut_payload_0_1086 ? _zz_dataOut_payload_0_1081 : _zz_dataOut_payload_0_1084);
    _zz_dataOut_payload_0_1089 <= (_zz_dataOut_payload_0_1086 ? _zz_dataOut_payload_0_1084 : _zz_dataOut_payload_0_1081);
    _zz_dataOut_payload_0_1090 <= (_zz_dataOut_payload_0_1087 ? _zz_dataOut_payload_0_1085 : _zz_dataOut_payload_0_1082);
    _zz_dataOut_payload_0_1091 <= (_zz_dataOut_payload_0_1087 ? _zz_dataOut_payload_0_1082 : _zz_dataOut_payload_0_1085);
    _zz_dataOut_payload_0_1100 <= (_zz_dataOut_payload_0_1098 ? _zz_dataOut_payload_0_1093 : _zz_dataOut_payload_0_1096);
    _zz_dataOut_payload_0_1101 <= (_zz_dataOut_payload_0_1098 ? _zz_dataOut_payload_0_1096 : _zz_dataOut_payload_0_1093);
    _zz_dataOut_payload_0_1102 <= (_zz_dataOut_payload_0_1099 ? _zz_dataOut_payload_0_1097 : _zz_dataOut_payload_0_1094);
    _zz_dataOut_payload_0_1103 <= (_zz_dataOut_payload_0_1099 ? _zz_dataOut_payload_0_1094 : _zz_dataOut_payload_0_1097);
    _zz_dataOut_payload_0_1112 <= (_zz_dataOut_payload_0_1110 ? _zz_dataOut_payload_0_1105 : _zz_dataOut_payload_0_1108);
    _zz_dataOut_payload_0_1113 <= (_zz_dataOut_payload_0_1110 ? _zz_dataOut_payload_0_1108 : _zz_dataOut_payload_0_1105);
    _zz_dataOut_payload_0_1114 <= (_zz_dataOut_payload_0_1111 ? _zz_dataOut_payload_0_1109 : _zz_dataOut_payload_0_1106);
    _zz_dataOut_payload_0_1115 <= (_zz_dataOut_payload_0_1111 ? _zz_dataOut_payload_0_1106 : _zz_dataOut_payload_0_1109);
    _zz_dataOut_payload_0_1124 <= (_zz_dataOut_payload_0_1122 ? _zz_dataOut_payload_0_1117 : _zz_dataOut_payload_0_1120);
    _zz_dataOut_payload_0_1125 <= (_zz_dataOut_payload_0_1122 ? _zz_dataOut_payload_0_1120 : _zz_dataOut_payload_0_1117);
    _zz_dataOut_payload_0_1126 <= (_zz_dataOut_payload_0_1123 ? _zz_dataOut_payload_0_1121 : _zz_dataOut_payload_0_1118);
    _zz_dataOut_payload_0_1127 <= (_zz_dataOut_payload_0_1123 ? _zz_dataOut_payload_0_1118 : _zz_dataOut_payload_0_1121);
    _zz_dataOut_payload_0_1136 <= (_zz_dataOut_payload_0_1134 ? _zz_dataOut_payload_0_1129 : _zz_dataOut_payload_0_1132);
    _zz_dataOut_payload_0_1137 <= (_zz_dataOut_payload_0_1134 ? _zz_dataOut_payload_0_1132 : _zz_dataOut_payload_0_1129);
    _zz_dataOut_payload_0_1138 <= (_zz_dataOut_payload_0_1135 ? _zz_dataOut_payload_0_1133 : _zz_dataOut_payload_0_1130);
    _zz_dataOut_payload_0_1139 <= (_zz_dataOut_payload_0_1135 ? _zz_dataOut_payload_0_1130 : _zz_dataOut_payload_0_1133);
    _zz_dataOut_payload_0_1148 <= (_zz_dataOut_payload_0_1146 ? _zz_dataOut_payload_0_1141 : _zz_dataOut_payload_0_1144);
    _zz_dataOut_payload_0_1149 <= (_zz_dataOut_payload_0_1146 ? _zz_dataOut_payload_0_1144 : _zz_dataOut_payload_0_1141);
    _zz_dataOut_payload_0_1150 <= (_zz_dataOut_payload_0_1147 ? _zz_dataOut_payload_0_1145 : _zz_dataOut_payload_0_1142);
    _zz_dataOut_payload_0_1151 <= (_zz_dataOut_payload_0_1147 ? _zz_dataOut_payload_0_1142 : _zz_dataOut_payload_0_1145);
    _zz_dataOut_payload_0_1152 <= _zz_dataOut_payload_0_392;
    _zz_dataOut_payload_0_1153 <= _zz_dataOut_payload_0_393;
    _zz_dataOut_payload_0_1154 <= _zz_dataOut_payload_0_394;
    _zz_dataOut_payload_0_1155 <= _zz_dataOut_payload_0_395;
    _zz_dataOut_payload_0_1156 <= _zz_dataOut_payload_0_404;
    _zz_dataOut_payload_0_1157 <= _zz_dataOut_payload_0_405;
    _zz_dataOut_payload_0_1158 <= _zz_dataOut_payload_0_406;
    _zz_dataOut_payload_0_1159 <= _zz_dataOut_payload_0_407;
    _zz_dataOut_payload_0_1160 <= _zz_dataOut_payload_0_416;
    _zz_dataOut_payload_0_1161 <= _zz_dataOut_payload_0_417;
    _zz_dataOut_payload_0_1162 <= _zz_dataOut_payload_0_418;
    _zz_dataOut_payload_0_1163 <= _zz_dataOut_payload_0_419;
    _zz_dataOut_payload_0_1164 <= _zz_dataOut_payload_0_428;
    _zz_dataOut_payload_0_1165 <= _zz_dataOut_payload_0_429;
    _zz_dataOut_payload_0_1166 <= _zz_dataOut_payload_0_430;
    _zz_dataOut_payload_0_1167 <= _zz_dataOut_payload_0_431;
    _zz_dataOut_payload_0_1168 <= _zz_dataOut_payload_0_440;
    _zz_dataOut_payload_0_1169 <= _zz_dataOut_payload_0_441;
    _zz_dataOut_payload_0_1170 <= _zz_dataOut_payload_0_442;
    _zz_dataOut_payload_0_1171 <= _zz_dataOut_payload_0_443;
    _zz_dataOut_payload_0_1172 <= _zz_dataOut_payload_0_452;
    _zz_dataOut_payload_0_1173 <= _zz_dataOut_payload_0_453;
    _zz_dataOut_payload_0_1174 <= _zz_dataOut_payload_0_454;
    _zz_dataOut_payload_0_1175 <= _zz_dataOut_payload_0_455;
    _zz_dataOut_payload_0_1176 <= _zz_dataOut_payload_0_464;
    _zz_dataOut_payload_0_1177 <= _zz_dataOut_payload_0_465;
    _zz_dataOut_payload_0_1178 <= _zz_dataOut_payload_0_466;
    _zz_dataOut_payload_0_1179 <= _zz_dataOut_payload_0_467;
    _zz_dataOut_payload_0_1180 <= _zz_dataOut_payload_0_476;
    _zz_dataOut_payload_0_1181 <= _zz_dataOut_payload_0_477;
    _zz_dataOut_payload_0_1182 <= _zz_dataOut_payload_0_478;
    _zz_dataOut_payload_0_1183 <= _zz_dataOut_payload_0_479;
    _zz_dataOut_payload_0_1184 <= _zz_dataOut_payload_0_488;
    _zz_dataOut_payload_0_1185 <= _zz_dataOut_payload_0_489;
    _zz_dataOut_payload_0_1186 <= _zz_dataOut_payload_0_490;
    _zz_dataOut_payload_0_1187 <= _zz_dataOut_payload_0_491;
    _zz_dataOut_payload_0_1188 <= _zz_dataOut_payload_0_500;
    _zz_dataOut_payload_0_1189 <= _zz_dataOut_payload_0_501;
    _zz_dataOut_payload_0_1190 <= _zz_dataOut_payload_0_502;
    _zz_dataOut_payload_0_1191 <= _zz_dataOut_payload_0_503;
    _zz_dataOut_payload_0_1192 <= _zz_dataOut_payload_0_512;
    _zz_dataOut_payload_0_1193 <= _zz_dataOut_payload_0_513;
    _zz_dataOut_payload_0_1194 <= _zz_dataOut_payload_0_514;
    _zz_dataOut_payload_0_1195 <= _zz_dataOut_payload_0_515;
    _zz_dataOut_payload_0_1196 <= _zz_dataOut_payload_0_524;
    _zz_dataOut_payload_0_1197 <= _zz_dataOut_payload_0_525;
    _zz_dataOut_payload_0_1198 <= _zz_dataOut_payload_0_526;
    _zz_dataOut_payload_0_1199 <= _zz_dataOut_payload_0_527;
    _zz_dataOut_payload_0_1200 <= _zz_dataOut_payload_0_536;
    _zz_dataOut_payload_0_1201 <= _zz_dataOut_payload_0_537;
    _zz_dataOut_payload_0_1202 <= _zz_dataOut_payload_0_538;
    _zz_dataOut_payload_0_1203 <= _zz_dataOut_payload_0_539;
    _zz_dataOut_payload_0_1204 <= _zz_dataOut_payload_0_548;
    _zz_dataOut_payload_0_1205 <= _zz_dataOut_payload_0_549;
    _zz_dataOut_payload_0_1206 <= _zz_dataOut_payload_0_550;
    _zz_dataOut_payload_0_1207 <= _zz_dataOut_payload_0_551;
    _zz_dataOut_payload_0_1208 <= _zz_dataOut_payload_0_560;
    _zz_dataOut_payload_0_1209 <= _zz_dataOut_payload_0_561;
    _zz_dataOut_payload_0_1210 <= _zz_dataOut_payload_0_562;
    _zz_dataOut_payload_0_1211 <= _zz_dataOut_payload_0_563;
    _zz_dataOut_payload_0_1212 <= _zz_dataOut_payload_0_572;
    _zz_dataOut_payload_0_1213 <= _zz_dataOut_payload_0_573;
    _zz_dataOut_payload_0_1214 <= _zz_dataOut_payload_0_574;
    _zz_dataOut_payload_0_1215 <= _zz_dataOut_payload_0_575;
    _zz_dataOut_payload_0_1216 <= _zz_dataOut_payload_0_584;
    _zz_dataOut_payload_0_1217 <= _zz_dataOut_payload_0_585;
    _zz_dataOut_payload_0_1218 <= _zz_dataOut_payload_0_586;
    _zz_dataOut_payload_0_1219 <= _zz_dataOut_payload_0_587;
    _zz_dataOut_payload_0_1220 <= _zz_dataOut_payload_0_596;
    _zz_dataOut_payload_0_1221 <= _zz_dataOut_payload_0_597;
    _zz_dataOut_payload_0_1222 <= _zz_dataOut_payload_0_598;
    _zz_dataOut_payload_0_1223 <= _zz_dataOut_payload_0_599;
    _zz_dataOut_payload_0_1224 <= _zz_dataOut_payload_0_608;
    _zz_dataOut_payload_0_1225 <= _zz_dataOut_payload_0_609;
    _zz_dataOut_payload_0_1226 <= _zz_dataOut_payload_0_610;
    _zz_dataOut_payload_0_1227 <= _zz_dataOut_payload_0_611;
    _zz_dataOut_payload_0_1228 <= _zz_dataOut_payload_0_620;
    _zz_dataOut_payload_0_1229 <= _zz_dataOut_payload_0_621;
    _zz_dataOut_payload_0_1230 <= _zz_dataOut_payload_0_622;
    _zz_dataOut_payload_0_1231 <= _zz_dataOut_payload_0_623;
    _zz_dataOut_payload_0_1232 <= _zz_dataOut_payload_0_632;
    _zz_dataOut_payload_0_1233 <= _zz_dataOut_payload_0_633;
    _zz_dataOut_payload_0_1234 <= _zz_dataOut_payload_0_634;
    _zz_dataOut_payload_0_1235 <= _zz_dataOut_payload_0_635;
    _zz_dataOut_payload_0_1236 <= _zz_dataOut_payload_0_644;
    _zz_dataOut_payload_0_1237 <= _zz_dataOut_payload_0_645;
    _zz_dataOut_payload_0_1238 <= _zz_dataOut_payload_0_646;
    _zz_dataOut_payload_0_1239 <= _zz_dataOut_payload_0_647;
    _zz_dataOut_payload_0_1240 <= _zz_dataOut_payload_0_656;
    _zz_dataOut_payload_0_1241 <= _zz_dataOut_payload_0_657;
    _zz_dataOut_payload_0_1242 <= _zz_dataOut_payload_0_658;
    _zz_dataOut_payload_0_1243 <= _zz_dataOut_payload_0_659;
    _zz_dataOut_payload_0_1244 <= _zz_dataOut_payload_0_668;
    _zz_dataOut_payload_0_1245 <= _zz_dataOut_payload_0_669;
    _zz_dataOut_payload_0_1246 <= _zz_dataOut_payload_0_670;
    _zz_dataOut_payload_0_1247 <= _zz_dataOut_payload_0_671;
    _zz_dataOut_payload_0_1248 <= _zz_dataOut_payload_0_680;
    _zz_dataOut_payload_0_1249 <= _zz_dataOut_payload_0_681;
    _zz_dataOut_payload_0_1250 <= _zz_dataOut_payload_0_682;
    _zz_dataOut_payload_0_1251 <= _zz_dataOut_payload_0_683;
    _zz_dataOut_payload_0_1252 <= _zz_dataOut_payload_0_692;
    _zz_dataOut_payload_0_1253 <= _zz_dataOut_payload_0_693;
    _zz_dataOut_payload_0_1254 <= _zz_dataOut_payload_0_694;
    _zz_dataOut_payload_0_1255 <= _zz_dataOut_payload_0_695;
    _zz_dataOut_payload_0_1256 <= _zz_dataOut_payload_0_704;
    _zz_dataOut_payload_0_1257 <= _zz_dataOut_payload_0_705;
    _zz_dataOut_payload_0_1258 <= _zz_dataOut_payload_0_706;
    _zz_dataOut_payload_0_1259 <= _zz_dataOut_payload_0_707;
    _zz_dataOut_payload_0_1260 <= _zz_dataOut_payload_0_716;
    _zz_dataOut_payload_0_1261 <= _zz_dataOut_payload_0_717;
    _zz_dataOut_payload_0_1262 <= _zz_dataOut_payload_0_718;
    _zz_dataOut_payload_0_1263 <= _zz_dataOut_payload_0_719;
    _zz_dataOut_payload_0_1264 <= _zz_dataOut_payload_0_728;
    _zz_dataOut_payload_0_1265 <= _zz_dataOut_payload_0_729;
    _zz_dataOut_payload_0_1266 <= _zz_dataOut_payload_0_730;
    _zz_dataOut_payload_0_1267 <= _zz_dataOut_payload_0_731;
    _zz_dataOut_payload_0_1268 <= _zz_dataOut_payload_0_740;
    _zz_dataOut_payload_0_1269 <= _zz_dataOut_payload_0_741;
    _zz_dataOut_payload_0_1270 <= _zz_dataOut_payload_0_742;
    _zz_dataOut_payload_0_1271 <= _zz_dataOut_payload_0_743;
    _zz_dataOut_payload_0_1272 <= _zz_dataOut_payload_0_752;
    _zz_dataOut_payload_0_1273 <= _zz_dataOut_payload_0_753;
    _zz_dataOut_payload_0_1274 <= _zz_dataOut_payload_0_754;
    _zz_dataOut_payload_0_1275 <= _zz_dataOut_payload_0_755;
    _zz_dataOut_payload_0_1276 <= _zz_dataOut_payload_0_764;
    _zz_dataOut_payload_0_1277 <= _zz_dataOut_payload_0_765;
    _zz_dataOut_payload_0_1278 <= _zz_dataOut_payload_0_766;
    _zz_dataOut_payload_0_1279 <= _zz_dataOut_payload_0_767;
    _zz_dataOut_payload_0_1280 <= _zz_dataOut_payload_0_776;
    _zz_dataOut_payload_0_1281 <= _zz_dataOut_payload_0_777;
    _zz_dataOut_payload_0_1282 <= _zz_dataOut_payload_0_778;
    _zz_dataOut_payload_0_1283 <= _zz_dataOut_payload_0_779;
    _zz_dataOut_payload_0_1284 <= _zz_dataOut_payload_0_788;
    _zz_dataOut_payload_0_1285 <= _zz_dataOut_payload_0_789;
    _zz_dataOut_payload_0_1286 <= _zz_dataOut_payload_0_790;
    _zz_dataOut_payload_0_1287 <= _zz_dataOut_payload_0_791;
    _zz_dataOut_payload_0_1288 <= _zz_dataOut_payload_0_800;
    _zz_dataOut_payload_0_1289 <= _zz_dataOut_payload_0_801;
    _zz_dataOut_payload_0_1290 <= _zz_dataOut_payload_0_802;
    _zz_dataOut_payload_0_1291 <= _zz_dataOut_payload_0_803;
    _zz_dataOut_payload_0_1292 <= _zz_dataOut_payload_0_812;
    _zz_dataOut_payload_0_1293 <= _zz_dataOut_payload_0_813;
    _zz_dataOut_payload_0_1294 <= _zz_dataOut_payload_0_814;
    _zz_dataOut_payload_0_1295 <= _zz_dataOut_payload_0_815;
    _zz_dataOut_payload_0_1296 <= _zz_dataOut_payload_0_824;
    _zz_dataOut_payload_0_1297 <= _zz_dataOut_payload_0_825;
    _zz_dataOut_payload_0_1298 <= _zz_dataOut_payload_0_826;
    _zz_dataOut_payload_0_1299 <= _zz_dataOut_payload_0_827;
    _zz_dataOut_payload_0_1300 <= _zz_dataOut_payload_0_836;
    _zz_dataOut_payload_0_1301 <= _zz_dataOut_payload_0_837;
    _zz_dataOut_payload_0_1302 <= _zz_dataOut_payload_0_838;
    _zz_dataOut_payload_0_1303 <= _zz_dataOut_payload_0_839;
    _zz_dataOut_payload_0_1304 <= _zz_dataOut_payload_0_848;
    _zz_dataOut_payload_0_1305 <= _zz_dataOut_payload_0_849;
    _zz_dataOut_payload_0_1306 <= _zz_dataOut_payload_0_850;
    _zz_dataOut_payload_0_1307 <= _zz_dataOut_payload_0_851;
    _zz_dataOut_payload_0_1308 <= _zz_dataOut_payload_0_860;
    _zz_dataOut_payload_0_1309 <= _zz_dataOut_payload_0_861;
    _zz_dataOut_payload_0_1310 <= _zz_dataOut_payload_0_862;
    _zz_dataOut_payload_0_1311 <= _zz_dataOut_payload_0_863;
    _zz_dataOut_payload_0_1312 <= _zz_dataOut_payload_0_872;
    _zz_dataOut_payload_0_1313 <= _zz_dataOut_payload_0_873;
    _zz_dataOut_payload_0_1314 <= _zz_dataOut_payload_0_874;
    _zz_dataOut_payload_0_1315 <= _zz_dataOut_payload_0_875;
    _zz_dataOut_payload_0_1316 <= _zz_dataOut_payload_0_884;
    _zz_dataOut_payload_0_1317 <= _zz_dataOut_payload_0_885;
    _zz_dataOut_payload_0_1318 <= _zz_dataOut_payload_0_886;
    _zz_dataOut_payload_0_1319 <= _zz_dataOut_payload_0_887;
    _zz_dataOut_payload_0_1320 <= _zz_dataOut_payload_0_896;
    _zz_dataOut_payload_0_1321 <= _zz_dataOut_payload_0_897;
    _zz_dataOut_payload_0_1322 <= _zz_dataOut_payload_0_898;
    _zz_dataOut_payload_0_1323 <= _zz_dataOut_payload_0_899;
    _zz_dataOut_payload_0_1324 <= _zz_dataOut_payload_0_908;
    _zz_dataOut_payload_0_1325 <= _zz_dataOut_payload_0_909;
    _zz_dataOut_payload_0_1326 <= _zz_dataOut_payload_0_910;
    _zz_dataOut_payload_0_1327 <= _zz_dataOut_payload_0_911;
    _zz_dataOut_payload_0_1328 <= _zz_dataOut_payload_0_920;
    _zz_dataOut_payload_0_1329 <= _zz_dataOut_payload_0_921;
    _zz_dataOut_payload_0_1330 <= _zz_dataOut_payload_0_922;
    _zz_dataOut_payload_0_1331 <= _zz_dataOut_payload_0_923;
    _zz_dataOut_payload_0_1332 <= _zz_dataOut_payload_0_932;
    _zz_dataOut_payload_0_1333 <= _zz_dataOut_payload_0_933;
    _zz_dataOut_payload_0_1334 <= _zz_dataOut_payload_0_934;
    _zz_dataOut_payload_0_1335 <= _zz_dataOut_payload_0_935;
    _zz_dataOut_payload_0_1336 <= _zz_dataOut_payload_0_944;
    _zz_dataOut_payload_0_1337 <= _zz_dataOut_payload_0_945;
    _zz_dataOut_payload_0_1338 <= _zz_dataOut_payload_0_946;
    _zz_dataOut_payload_0_1339 <= _zz_dataOut_payload_0_947;
    _zz_dataOut_payload_0_1340 <= _zz_dataOut_payload_0_956;
    _zz_dataOut_payload_0_1341 <= _zz_dataOut_payload_0_957;
    _zz_dataOut_payload_0_1342 <= _zz_dataOut_payload_0_958;
    _zz_dataOut_payload_0_1343 <= _zz_dataOut_payload_0_959;
    _zz_dataOut_payload_0_1344 <= _zz_dataOut_payload_0_968;
    _zz_dataOut_payload_0_1345 <= _zz_dataOut_payload_0_969;
    _zz_dataOut_payload_0_1346 <= _zz_dataOut_payload_0_970;
    _zz_dataOut_payload_0_1347 <= _zz_dataOut_payload_0_971;
    _zz_dataOut_payload_0_1348 <= _zz_dataOut_payload_0_980;
    _zz_dataOut_payload_0_1349 <= _zz_dataOut_payload_0_981;
    _zz_dataOut_payload_0_1350 <= _zz_dataOut_payload_0_982;
    _zz_dataOut_payload_0_1351 <= _zz_dataOut_payload_0_983;
    _zz_dataOut_payload_0_1352 <= _zz_dataOut_payload_0_992;
    _zz_dataOut_payload_0_1353 <= _zz_dataOut_payload_0_993;
    _zz_dataOut_payload_0_1354 <= _zz_dataOut_payload_0_994;
    _zz_dataOut_payload_0_1355 <= _zz_dataOut_payload_0_995;
    _zz_dataOut_payload_0_1356 <= _zz_dataOut_payload_0_1004;
    _zz_dataOut_payload_0_1357 <= _zz_dataOut_payload_0_1005;
    _zz_dataOut_payload_0_1358 <= _zz_dataOut_payload_0_1006;
    _zz_dataOut_payload_0_1359 <= _zz_dataOut_payload_0_1007;
    _zz_dataOut_payload_0_1360 <= _zz_dataOut_payload_0_1016;
    _zz_dataOut_payload_0_1361 <= _zz_dataOut_payload_0_1017;
    _zz_dataOut_payload_0_1362 <= _zz_dataOut_payload_0_1018;
    _zz_dataOut_payload_0_1363 <= _zz_dataOut_payload_0_1019;
    _zz_dataOut_payload_0_1364 <= _zz_dataOut_payload_0_1028;
    _zz_dataOut_payload_0_1365 <= _zz_dataOut_payload_0_1029;
    _zz_dataOut_payload_0_1366 <= _zz_dataOut_payload_0_1030;
    _zz_dataOut_payload_0_1367 <= _zz_dataOut_payload_0_1031;
    _zz_dataOut_payload_0_1368 <= _zz_dataOut_payload_0_1040;
    _zz_dataOut_payload_0_1369 <= _zz_dataOut_payload_0_1041;
    _zz_dataOut_payload_0_1370 <= _zz_dataOut_payload_0_1042;
    _zz_dataOut_payload_0_1371 <= _zz_dataOut_payload_0_1043;
    _zz_dataOut_payload_0_1372 <= _zz_dataOut_payload_0_1052;
    _zz_dataOut_payload_0_1373 <= _zz_dataOut_payload_0_1053;
    _zz_dataOut_payload_0_1374 <= _zz_dataOut_payload_0_1054;
    _zz_dataOut_payload_0_1375 <= _zz_dataOut_payload_0_1055;
    _zz_dataOut_payload_0_1376 <= _zz_dataOut_payload_0_1064;
    _zz_dataOut_payload_0_1377 <= _zz_dataOut_payload_0_1065;
    _zz_dataOut_payload_0_1378 <= _zz_dataOut_payload_0_1066;
    _zz_dataOut_payload_0_1379 <= _zz_dataOut_payload_0_1067;
    _zz_dataOut_payload_0_1380 <= _zz_dataOut_payload_0_1076;
    _zz_dataOut_payload_0_1381 <= _zz_dataOut_payload_0_1077;
    _zz_dataOut_payload_0_1382 <= _zz_dataOut_payload_0_1078;
    _zz_dataOut_payload_0_1383 <= _zz_dataOut_payload_0_1079;
    _zz_dataOut_payload_0_1384 <= _zz_dataOut_payload_0_1088;
    _zz_dataOut_payload_0_1385 <= _zz_dataOut_payload_0_1089;
    _zz_dataOut_payload_0_1386 <= _zz_dataOut_payload_0_1090;
    _zz_dataOut_payload_0_1387 <= _zz_dataOut_payload_0_1091;
    _zz_dataOut_payload_0_1388 <= _zz_dataOut_payload_0_1100;
    _zz_dataOut_payload_0_1389 <= _zz_dataOut_payload_0_1101;
    _zz_dataOut_payload_0_1390 <= _zz_dataOut_payload_0_1102;
    _zz_dataOut_payload_0_1391 <= _zz_dataOut_payload_0_1103;
    _zz_dataOut_payload_0_1392 <= _zz_dataOut_payload_0_1112;
    _zz_dataOut_payload_0_1393 <= _zz_dataOut_payload_0_1113;
    _zz_dataOut_payload_0_1394 <= _zz_dataOut_payload_0_1114;
    _zz_dataOut_payload_0_1395 <= _zz_dataOut_payload_0_1115;
    _zz_dataOut_payload_0_1396 <= _zz_dataOut_payload_0_1124;
    _zz_dataOut_payload_0_1397 <= _zz_dataOut_payload_0_1125;
    _zz_dataOut_payload_0_1398 <= _zz_dataOut_payload_0_1126;
    _zz_dataOut_payload_0_1399 <= _zz_dataOut_payload_0_1127;
    _zz_dataOut_payload_0_1400 <= _zz_dataOut_payload_0_1136;
    _zz_dataOut_payload_0_1401 <= _zz_dataOut_payload_0_1137;
    _zz_dataOut_payload_0_1402 <= _zz_dataOut_payload_0_1138;
    _zz_dataOut_payload_0_1403 <= _zz_dataOut_payload_0_1139;
    _zz_dataOut_payload_0_1404 <= _zz_dataOut_payload_0_1148;
    _zz_dataOut_payload_0_1405 <= _zz_dataOut_payload_0_1149;
    _zz_dataOut_payload_0_1406 <= _zz_dataOut_payload_0_1150;
    _zz_dataOut_payload_0_1407 <= _zz_dataOut_payload_0_1151;
    _zz_dataOut_payload_0_1428 <= (_zz_dataOut_payload_0_1426 ? _zz_dataOut_payload_0_1421 : _zz_dataOut_payload_0_1424);
    _zz_dataOut_payload_0_1429 <= (_zz_dataOut_payload_0_1426 ? _zz_dataOut_payload_0_1424 : _zz_dataOut_payload_0_1421);
    _zz_dataOut_payload_0_1430 <= (_zz_dataOut_payload_0_1427 ? _zz_dataOut_payload_0_1422 : _zz_dataOut_payload_0_1425);
    _zz_dataOut_payload_0_1431 <= (_zz_dataOut_payload_0_1427 ? _zz_dataOut_payload_0_1425 : _zz_dataOut_payload_0_1422);
    _zz_dataOut_payload_0_1440 <= (_zz_dataOut_payload_0_1438 ? _zz_dataOut_payload_0_1433 : _zz_dataOut_payload_0_1436);
    _zz_dataOut_payload_0_1441 <= (_zz_dataOut_payload_0_1438 ? _zz_dataOut_payload_0_1436 : _zz_dataOut_payload_0_1433);
    _zz_dataOut_payload_0_1442 <= (_zz_dataOut_payload_0_1439 ? _zz_dataOut_payload_0_1434 : _zz_dataOut_payload_0_1437);
    _zz_dataOut_payload_0_1443 <= (_zz_dataOut_payload_0_1439 ? _zz_dataOut_payload_0_1437 : _zz_dataOut_payload_0_1434);
    _zz_dataOut_payload_0_1444 <= _zz_dataOut_payload_0_1428;
    _zz_dataOut_payload_0_1445 <= _zz_dataOut_payload_0_1429;
    _zz_dataOut_payload_0_1446 <= _zz_dataOut_payload_0_1430;
    _zz_dataOut_payload_0_1447 <= _zz_dataOut_payload_0_1431;
    _zz_dataOut_payload_0_1448 <= _zz_dataOut_payload_0_1440;
    _zz_dataOut_payload_0_1449 <= _zz_dataOut_payload_0_1441;
    _zz_dataOut_payload_0_1450 <= _zz_dataOut_payload_0_1442;
    _zz_dataOut_payload_0_1451 <= _zz_dataOut_payload_0_1443;
    _zz_dataOut_payload_0_1472 <= (_zz_dataOut_payload_0_1470 ? _zz_dataOut_payload_0_1465 : _zz_dataOut_payload_0_1468);
    _zz_dataOut_payload_0_1473 <= (_zz_dataOut_payload_0_1470 ? _zz_dataOut_payload_0_1468 : _zz_dataOut_payload_0_1465);
    _zz_dataOut_payload_0_1474 <= (_zz_dataOut_payload_0_1471 ? _zz_dataOut_payload_0_1466 : _zz_dataOut_payload_0_1469);
    _zz_dataOut_payload_0_1475 <= (_zz_dataOut_payload_0_1471 ? _zz_dataOut_payload_0_1469 : _zz_dataOut_payload_0_1466);
    _zz_dataOut_payload_0_1484 <= (_zz_dataOut_payload_0_1482 ? _zz_dataOut_payload_0_1477 : _zz_dataOut_payload_0_1480);
    _zz_dataOut_payload_0_1485 <= (_zz_dataOut_payload_0_1482 ? _zz_dataOut_payload_0_1480 : _zz_dataOut_payload_0_1477);
    _zz_dataOut_payload_0_1486 <= (_zz_dataOut_payload_0_1483 ? _zz_dataOut_payload_0_1478 : _zz_dataOut_payload_0_1481);
    _zz_dataOut_payload_0_1487 <= (_zz_dataOut_payload_0_1483 ? _zz_dataOut_payload_0_1481 : _zz_dataOut_payload_0_1478);
    _zz_dataOut_payload_0_1488 <= _zz_dataOut_payload_0_1472;
    _zz_dataOut_payload_0_1489 <= _zz_dataOut_payload_0_1473;
    _zz_dataOut_payload_0_1490 <= _zz_dataOut_payload_0_1474;
    _zz_dataOut_payload_0_1491 <= _zz_dataOut_payload_0_1475;
    _zz_dataOut_payload_0_1492 <= _zz_dataOut_payload_0_1484;
    _zz_dataOut_payload_0_1493 <= _zz_dataOut_payload_0_1485;
    _zz_dataOut_payload_0_1494 <= _zz_dataOut_payload_0_1486;
    _zz_dataOut_payload_0_1495 <= _zz_dataOut_payload_0_1487;
    _zz_dataOut_payload_0_1516 <= (_zz_dataOut_payload_0_1514 ? _zz_dataOut_payload_0_1509 : _zz_dataOut_payload_0_1512);
    _zz_dataOut_payload_0_1517 <= (_zz_dataOut_payload_0_1514 ? _zz_dataOut_payload_0_1512 : _zz_dataOut_payload_0_1509);
    _zz_dataOut_payload_0_1518 <= (_zz_dataOut_payload_0_1515 ? _zz_dataOut_payload_0_1510 : _zz_dataOut_payload_0_1513);
    _zz_dataOut_payload_0_1519 <= (_zz_dataOut_payload_0_1515 ? _zz_dataOut_payload_0_1513 : _zz_dataOut_payload_0_1510);
    _zz_dataOut_payload_0_1528 <= (_zz_dataOut_payload_0_1526 ? _zz_dataOut_payload_0_1521 : _zz_dataOut_payload_0_1524);
    _zz_dataOut_payload_0_1529 <= (_zz_dataOut_payload_0_1526 ? _zz_dataOut_payload_0_1524 : _zz_dataOut_payload_0_1521);
    _zz_dataOut_payload_0_1530 <= (_zz_dataOut_payload_0_1527 ? _zz_dataOut_payload_0_1522 : _zz_dataOut_payload_0_1525);
    _zz_dataOut_payload_0_1531 <= (_zz_dataOut_payload_0_1527 ? _zz_dataOut_payload_0_1525 : _zz_dataOut_payload_0_1522);
    _zz_dataOut_payload_0_1532 <= _zz_dataOut_payload_0_1516;
    _zz_dataOut_payload_0_1533 <= _zz_dataOut_payload_0_1517;
    _zz_dataOut_payload_0_1534 <= _zz_dataOut_payload_0_1518;
    _zz_dataOut_payload_0_1535 <= _zz_dataOut_payload_0_1519;
    _zz_dataOut_payload_0_1536 <= _zz_dataOut_payload_0_1528;
    _zz_dataOut_payload_0_1537 <= _zz_dataOut_payload_0_1529;
    _zz_dataOut_payload_0_1538 <= _zz_dataOut_payload_0_1530;
    _zz_dataOut_payload_0_1539 <= _zz_dataOut_payload_0_1531;
    _zz_dataOut_payload_0_1560 <= (_zz_dataOut_payload_0_1558 ? _zz_dataOut_payload_0_1553 : _zz_dataOut_payload_0_1556);
    _zz_dataOut_payload_0_1561 <= (_zz_dataOut_payload_0_1558 ? _zz_dataOut_payload_0_1556 : _zz_dataOut_payload_0_1553);
    _zz_dataOut_payload_0_1562 <= (_zz_dataOut_payload_0_1559 ? _zz_dataOut_payload_0_1554 : _zz_dataOut_payload_0_1557);
    _zz_dataOut_payload_0_1563 <= (_zz_dataOut_payload_0_1559 ? _zz_dataOut_payload_0_1557 : _zz_dataOut_payload_0_1554);
    _zz_dataOut_payload_0_1572 <= (_zz_dataOut_payload_0_1570 ? _zz_dataOut_payload_0_1565 : _zz_dataOut_payload_0_1568);
    _zz_dataOut_payload_0_1573 <= (_zz_dataOut_payload_0_1570 ? _zz_dataOut_payload_0_1568 : _zz_dataOut_payload_0_1565);
    _zz_dataOut_payload_0_1574 <= (_zz_dataOut_payload_0_1571 ? _zz_dataOut_payload_0_1566 : _zz_dataOut_payload_0_1569);
    _zz_dataOut_payload_0_1575 <= (_zz_dataOut_payload_0_1571 ? _zz_dataOut_payload_0_1569 : _zz_dataOut_payload_0_1566);
    _zz_dataOut_payload_0_1576 <= _zz_dataOut_payload_0_1560;
    _zz_dataOut_payload_0_1577 <= _zz_dataOut_payload_0_1561;
    _zz_dataOut_payload_0_1578 <= _zz_dataOut_payload_0_1562;
    _zz_dataOut_payload_0_1579 <= _zz_dataOut_payload_0_1563;
    _zz_dataOut_payload_0_1580 <= _zz_dataOut_payload_0_1572;
    _zz_dataOut_payload_0_1581 <= _zz_dataOut_payload_0_1573;
    _zz_dataOut_payload_0_1582 <= _zz_dataOut_payload_0_1574;
    _zz_dataOut_payload_0_1583 <= _zz_dataOut_payload_0_1575;
    _zz_dataOut_payload_0_1604 <= (_zz_dataOut_payload_0_1602 ? _zz_dataOut_payload_0_1597 : _zz_dataOut_payload_0_1600);
    _zz_dataOut_payload_0_1605 <= (_zz_dataOut_payload_0_1602 ? _zz_dataOut_payload_0_1600 : _zz_dataOut_payload_0_1597);
    _zz_dataOut_payload_0_1606 <= (_zz_dataOut_payload_0_1603 ? _zz_dataOut_payload_0_1598 : _zz_dataOut_payload_0_1601);
    _zz_dataOut_payload_0_1607 <= (_zz_dataOut_payload_0_1603 ? _zz_dataOut_payload_0_1601 : _zz_dataOut_payload_0_1598);
    _zz_dataOut_payload_0_1616 <= (_zz_dataOut_payload_0_1614 ? _zz_dataOut_payload_0_1609 : _zz_dataOut_payload_0_1612);
    _zz_dataOut_payload_0_1617 <= (_zz_dataOut_payload_0_1614 ? _zz_dataOut_payload_0_1612 : _zz_dataOut_payload_0_1609);
    _zz_dataOut_payload_0_1618 <= (_zz_dataOut_payload_0_1615 ? _zz_dataOut_payload_0_1610 : _zz_dataOut_payload_0_1613);
    _zz_dataOut_payload_0_1619 <= (_zz_dataOut_payload_0_1615 ? _zz_dataOut_payload_0_1613 : _zz_dataOut_payload_0_1610);
    _zz_dataOut_payload_0_1620 <= _zz_dataOut_payload_0_1604;
    _zz_dataOut_payload_0_1621 <= _zz_dataOut_payload_0_1605;
    _zz_dataOut_payload_0_1622 <= _zz_dataOut_payload_0_1606;
    _zz_dataOut_payload_0_1623 <= _zz_dataOut_payload_0_1607;
    _zz_dataOut_payload_0_1624 <= _zz_dataOut_payload_0_1616;
    _zz_dataOut_payload_0_1625 <= _zz_dataOut_payload_0_1617;
    _zz_dataOut_payload_0_1626 <= _zz_dataOut_payload_0_1618;
    _zz_dataOut_payload_0_1627 <= _zz_dataOut_payload_0_1619;
    _zz_dataOut_payload_0_1648 <= (_zz_dataOut_payload_0_1646 ? _zz_dataOut_payload_0_1641 : _zz_dataOut_payload_0_1644);
    _zz_dataOut_payload_0_1649 <= (_zz_dataOut_payload_0_1646 ? _zz_dataOut_payload_0_1644 : _zz_dataOut_payload_0_1641);
    _zz_dataOut_payload_0_1650 <= (_zz_dataOut_payload_0_1647 ? _zz_dataOut_payload_0_1642 : _zz_dataOut_payload_0_1645);
    _zz_dataOut_payload_0_1651 <= (_zz_dataOut_payload_0_1647 ? _zz_dataOut_payload_0_1645 : _zz_dataOut_payload_0_1642);
    _zz_dataOut_payload_0_1660 <= (_zz_dataOut_payload_0_1658 ? _zz_dataOut_payload_0_1653 : _zz_dataOut_payload_0_1656);
    _zz_dataOut_payload_0_1661 <= (_zz_dataOut_payload_0_1658 ? _zz_dataOut_payload_0_1656 : _zz_dataOut_payload_0_1653);
    _zz_dataOut_payload_0_1662 <= (_zz_dataOut_payload_0_1659 ? _zz_dataOut_payload_0_1654 : _zz_dataOut_payload_0_1657);
    _zz_dataOut_payload_0_1663 <= (_zz_dataOut_payload_0_1659 ? _zz_dataOut_payload_0_1657 : _zz_dataOut_payload_0_1654);
    _zz_dataOut_payload_0_1664 <= _zz_dataOut_payload_0_1648;
    _zz_dataOut_payload_0_1665 <= _zz_dataOut_payload_0_1649;
    _zz_dataOut_payload_0_1666 <= _zz_dataOut_payload_0_1650;
    _zz_dataOut_payload_0_1667 <= _zz_dataOut_payload_0_1651;
    _zz_dataOut_payload_0_1668 <= _zz_dataOut_payload_0_1660;
    _zz_dataOut_payload_0_1669 <= _zz_dataOut_payload_0_1661;
    _zz_dataOut_payload_0_1670 <= _zz_dataOut_payload_0_1662;
    _zz_dataOut_payload_0_1671 <= _zz_dataOut_payload_0_1663;
    _zz_dataOut_payload_0_1692 <= (_zz_dataOut_payload_0_1690 ? _zz_dataOut_payload_0_1685 : _zz_dataOut_payload_0_1688);
    _zz_dataOut_payload_0_1693 <= (_zz_dataOut_payload_0_1690 ? _zz_dataOut_payload_0_1688 : _zz_dataOut_payload_0_1685);
    _zz_dataOut_payload_0_1694 <= (_zz_dataOut_payload_0_1691 ? _zz_dataOut_payload_0_1686 : _zz_dataOut_payload_0_1689);
    _zz_dataOut_payload_0_1695 <= (_zz_dataOut_payload_0_1691 ? _zz_dataOut_payload_0_1689 : _zz_dataOut_payload_0_1686);
    _zz_dataOut_payload_0_1704 <= (_zz_dataOut_payload_0_1702 ? _zz_dataOut_payload_0_1697 : _zz_dataOut_payload_0_1700);
    _zz_dataOut_payload_0_1705 <= (_zz_dataOut_payload_0_1702 ? _zz_dataOut_payload_0_1700 : _zz_dataOut_payload_0_1697);
    _zz_dataOut_payload_0_1706 <= (_zz_dataOut_payload_0_1703 ? _zz_dataOut_payload_0_1698 : _zz_dataOut_payload_0_1701);
    _zz_dataOut_payload_0_1707 <= (_zz_dataOut_payload_0_1703 ? _zz_dataOut_payload_0_1701 : _zz_dataOut_payload_0_1698);
    _zz_dataOut_payload_0_1708 <= _zz_dataOut_payload_0_1692;
    _zz_dataOut_payload_0_1709 <= _zz_dataOut_payload_0_1693;
    _zz_dataOut_payload_0_1710 <= _zz_dataOut_payload_0_1694;
    _zz_dataOut_payload_0_1711 <= _zz_dataOut_payload_0_1695;
    _zz_dataOut_payload_0_1712 <= _zz_dataOut_payload_0_1704;
    _zz_dataOut_payload_0_1713 <= _zz_dataOut_payload_0_1705;
    _zz_dataOut_payload_0_1714 <= _zz_dataOut_payload_0_1706;
    _zz_dataOut_payload_0_1715 <= _zz_dataOut_payload_0_1707;
    _zz_dataOut_payload_0_1736 <= (_zz_dataOut_payload_0_1734 ? _zz_dataOut_payload_0_1729 : _zz_dataOut_payload_0_1732);
    _zz_dataOut_payload_0_1737 <= (_zz_dataOut_payload_0_1734 ? _zz_dataOut_payload_0_1732 : _zz_dataOut_payload_0_1729);
    _zz_dataOut_payload_0_1738 <= (_zz_dataOut_payload_0_1735 ? _zz_dataOut_payload_0_1730 : _zz_dataOut_payload_0_1733);
    _zz_dataOut_payload_0_1739 <= (_zz_dataOut_payload_0_1735 ? _zz_dataOut_payload_0_1733 : _zz_dataOut_payload_0_1730);
    _zz_dataOut_payload_0_1748 <= (_zz_dataOut_payload_0_1746 ? _zz_dataOut_payload_0_1741 : _zz_dataOut_payload_0_1744);
    _zz_dataOut_payload_0_1749 <= (_zz_dataOut_payload_0_1746 ? _zz_dataOut_payload_0_1744 : _zz_dataOut_payload_0_1741);
    _zz_dataOut_payload_0_1750 <= (_zz_dataOut_payload_0_1747 ? _zz_dataOut_payload_0_1742 : _zz_dataOut_payload_0_1745);
    _zz_dataOut_payload_0_1751 <= (_zz_dataOut_payload_0_1747 ? _zz_dataOut_payload_0_1745 : _zz_dataOut_payload_0_1742);
    _zz_dataOut_payload_0_1752 <= _zz_dataOut_payload_0_1736;
    _zz_dataOut_payload_0_1753 <= _zz_dataOut_payload_0_1737;
    _zz_dataOut_payload_0_1754 <= _zz_dataOut_payload_0_1738;
    _zz_dataOut_payload_0_1755 <= _zz_dataOut_payload_0_1739;
    _zz_dataOut_payload_0_1756 <= _zz_dataOut_payload_0_1748;
    _zz_dataOut_payload_0_1757 <= _zz_dataOut_payload_0_1749;
    _zz_dataOut_payload_0_1758 <= _zz_dataOut_payload_0_1750;
    _zz_dataOut_payload_0_1759 <= _zz_dataOut_payload_0_1751;
    _zz_dataOut_payload_0_1780 <= (_zz_dataOut_payload_0_1778 ? _zz_dataOut_payload_0_1773 : _zz_dataOut_payload_0_1776);
    _zz_dataOut_payload_0_1781 <= (_zz_dataOut_payload_0_1778 ? _zz_dataOut_payload_0_1776 : _zz_dataOut_payload_0_1773);
    _zz_dataOut_payload_0_1782 <= (_zz_dataOut_payload_0_1779 ? _zz_dataOut_payload_0_1774 : _zz_dataOut_payload_0_1777);
    _zz_dataOut_payload_0_1783 <= (_zz_dataOut_payload_0_1779 ? _zz_dataOut_payload_0_1777 : _zz_dataOut_payload_0_1774);
    _zz_dataOut_payload_0_1792 <= (_zz_dataOut_payload_0_1790 ? _zz_dataOut_payload_0_1785 : _zz_dataOut_payload_0_1788);
    _zz_dataOut_payload_0_1793 <= (_zz_dataOut_payload_0_1790 ? _zz_dataOut_payload_0_1788 : _zz_dataOut_payload_0_1785);
    _zz_dataOut_payload_0_1794 <= (_zz_dataOut_payload_0_1791 ? _zz_dataOut_payload_0_1786 : _zz_dataOut_payload_0_1789);
    _zz_dataOut_payload_0_1795 <= (_zz_dataOut_payload_0_1791 ? _zz_dataOut_payload_0_1789 : _zz_dataOut_payload_0_1786);
    _zz_dataOut_payload_0_1796 <= _zz_dataOut_payload_0_1780;
    _zz_dataOut_payload_0_1797 <= _zz_dataOut_payload_0_1781;
    _zz_dataOut_payload_0_1798 <= _zz_dataOut_payload_0_1782;
    _zz_dataOut_payload_0_1799 <= _zz_dataOut_payload_0_1783;
    _zz_dataOut_payload_0_1800 <= _zz_dataOut_payload_0_1792;
    _zz_dataOut_payload_0_1801 <= _zz_dataOut_payload_0_1793;
    _zz_dataOut_payload_0_1802 <= _zz_dataOut_payload_0_1794;
    _zz_dataOut_payload_0_1803 <= _zz_dataOut_payload_0_1795;
    _zz_dataOut_payload_0_1824 <= (_zz_dataOut_payload_0_1822 ? _zz_dataOut_payload_0_1817 : _zz_dataOut_payload_0_1820);
    _zz_dataOut_payload_0_1825 <= (_zz_dataOut_payload_0_1822 ? _zz_dataOut_payload_0_1820 : _zz_dataOut_payload_0_1817);
    _zz_dataOut_payload_0_1826 <= (_zz_dataOut_payload_0_1823 ? _zz_dataOut_payload_0_1818 : _zz_dataOut_payload_0_1821);
    _zz_dataOut_payload_0_1827 <= (_zz_dataOut_payload_0_1823 ? _zz_dataOut_payload_0_1821 : _zz_dataOut_payload_0_1818);
    _zz_dataOut_payload_0_1836 <= (_zz_dataOut_payload_0_1834 ? _zz_dataOut_payload_0_1829 : _zz_dataOut_payload_0_1832);
    _zz_dataOut_payload_0_1837 <= (_zz_dataOut_payload_0_1834 ? _zz_dataOut_payload_0_1832 : _zz_dataOut_payload_0_1829);
    _zz_dataOut_payload_0_1838 <= (_zz_dataOut_payload_0_1835 ? _zz_dataOut_payload_0_1830 : _zz_dataOut_payload_0_1833);
    _zz_dataOut_payload_0_1839 <= (_zz_dataOut_payload_0_1835 ? _zz_dataOut_payload_0_1833 : _zz_dataOut_payload_0_1830);
    _zz_dataOut_payload_0_1840 <= _zz_dataOut_payload_0_1824;
    _zz_dataOut_payload_0_1841 <= _zz_dataOut_payload_0_1825;
    _zz_dataOut_payload_0_1842 <= _zz_dataOut_payload_0_1826;
    _zz_dataOut_payload_0_1843 <= _zz_dataOut_payload_0_1827;
    _zz_dataOut_payload_0_1844 <= _zz_dataOut_payload_0_1836;
    _zz_dataOut_payload_0_1845 <= _zz_dataOut_payload_0_1837;
    _zz_dataOut_payload_0_1846 <= _zz_dataOut_payload_0_1838;
    _zz_dataOut_payload_0_1847 <= _zz_dataOut_payload_0_1839;
    _zz_dataOut_payload_0_1868 <= (_zz_dataOut_payload_0_1866 ? _zz_dataOut_payload_0_1861 : _zz_dataOut_payload_0_1864);
    _zz_dataOut_payload_0_1869 <= (_zz_dataOut_payload_0_1866 ? _zz_dataOut_payload_0_1864 : _zz_dataOut_payload_0_1861);
    _zz_dataOut_payload_0_1870 <= (_zz_dataOut_payload_0_1867 ? _zz_dataOut_payload_0_1862 : _zz_dataOut_payload_0_1865);
    _zz_dataOut_payload_0_1871 <= (_zz_dataOut_payload_0_1867 ? _zz_dataOut_payload_0_1865 : _zz_dataOut_payload_0_1862);
    _zz_dataOut_payload_0_1880 <= (_zz_dataOut_payload_0_1878 ? _zz_dataOut_payload_0_1873 : _zz_dataOut_payload_0_1876);
    _zz_dataOut_payload_0_1881 <= (_zz_dataOut_payload_0_1878 ? _zz_dataOut_payload_0_1876 : _zz_dataOut_payload_0_1873);
    _zz_dataOut_payload_0_1882 <= (_zz_dataOut_payload_0_1879 ? _zz_dataOut_payload_0_1874 : _zz_dataOut_payload_0_1877);
    _zz_dataOut_payload_0_1883 <= (_zz_dataOut_payload_0_1879 ? _zz_dataOut_payload_0_1877 : _zz_dataOut_payload_0_1874);
    _zz_dataOut_payload_0_1884 <= _zz_dataOut_payload_0_1868;
    _zz_dataOut_payload_0_1885 <= _zz_dataOut_payload_0_1869;
    _zz_dataOut_payload_0_1886 <= _zz_dataOut_payload_0_1870;
    _zz_dataOut_payload_0_1887 <= _zz_dataOut_payload_0_1871;
    _zz_dataOut_payload_0_1888 <= _zz_dataOut_payload_0_1880;
    _zz_dataOut_payload_0_1889 <= _zz_dataOut_payload_0_1881;
    _zz_dataOut_payload_0_1890 <= _zz_dataOut_payload_0_1882;
    _zz_dataOut_payload_0_1891 <= _zz_dataOut_payload_0_1883;
    _zz_dataOut_payload_0_1912 <= (_zz_dataOut_payload_0_1910 ? _zz_dataOut_payload_0_1905 : _zz_dataOut_payload_0_1908);
    _zz_dataOut_payload_0_1913 <= (_zz_dataOut_payload_0_1910 ? _zz_dataOut_payload_0_1908 : _zz_dataOut_payload_0_1905);
    _zz_dataOut_payload_0_1914 <= (_zz_dataOut_payload_0_1911 ? _zz_dataOut_payload_0_1906 : _zz_dataOut_payload_0_1909);
    _zz_dataOut_payload_0_1915 <= (_zz_dataOut_payload_0_1911 ? _zz_dataOut_payload_0_1909 : _zz_dataOut_payload_0_1906);
    _zz_dataOut_payload_0_1924 <= (_zz_dataOut_payload_0_1922 ? _zz_dataOut_payload_0_1917 : _zz_dataOut_payload_0_1920);
    _zz_dataOut_payload_0_1925 <= (_zz_dataOut_payload_0_1922 ? _zz_dataOut_payload_0_1920 : _zz_dataOut_payload_0_1917);
    _zz_dataOut_payload_0_1926 <= (_zz_dataOut_payload_0_1923 ? _zz_dataOut_payload_0_1918 : _zz_dataOut_payload_0_1921);
    _zz_dataOut_payload_0_1927 <= (_zz_dataOut_payload_0_1923 ? _zz_dataOut_payload_0_1921 : _zz_dataOut_payload_0_1918);
    _zz_dataOut_payload_0_1928 <= _zz_dataOut_payload_0_1912;
    _zz_dataOut_payload_0_1929 <= _zz_dataOut_payload_0_1913;
    _zz_dataOut_payload_0_1930 <= _zz_dataOut_payload_0_1914;
    _zz_dataOut_payload_0_1931 <= _zz_dataOut_payload_0_1915;
    _zz_dataOut_payload_0_1932 <= _zz_dataOut_payload_0_1924;
    _zz_dataOut_payload_0_1933 <= _zz_dataOut_payload_0_1925;
    _zz_dataOut_payload_0_1934 <= _zz_dataOut_payload_0_1926;
    _zz_dataOut_payload_0_1935 <= _zz_dataOut_payload_0_1927;
    _zz_dataOut_payload_0_1956 <= (_zz_dataOut_payload_0_1954 ? _zz_dataOut_payload_0_1949 : _zz_dataOut_payload_0_1952);
    _zz_dataOut_payload_0_1957 <= (_zz_dataOut_payload_0_1954 ? _zz_dataOut_payload_0_1952 : _zz_dataOut_payload_0_1949);
    _zz_dataOut_payload_0_1958 <= (_zz_dataOut_payload_0_1955 ? _zz_dataOut_payload_0_1950 : _zz_dataOut_payload_0_1953);
    _zz_dataOut_payload_0_1959 <= (_zz_dataOut_payload_0_1955 ? _zz_dataOut_payload_0_1953 : _zz_dataOut_payload_0_1950);
    _zz_dataOut_payload_0_1968 <= (_zz_dataOut_payload_0_1966 ? _zz_dataOut_payload_0_1961 : _zz_dataOut_payload_0_1964);
    _zz_dataOut_payload_0_1969 <= (_zz_dataOut_payload_0_1966 ? _zz_dataOut_payload_0_1964 : _zz_dataOut_payload_0_1961);
    _zz_dataOut_payload_0_1970 <= (_zz_dataOut_payload_0_1967 ? _zz_dataOut_payload_0_1962 : _zz_dataOut_payload_0_1965);
    _zz_dataOut_payload_0_1971 <= (_zz_dataOut_payload_0_1967 ? _zz_dataOut_payload_0_1965 : _zz_dataOut_payload_0_1962);
    _zz_dataOut_payload_0_1972 <= _zz_dataOut_payload_0_1956;
    _zz_dataOut_payload_0_1973 <= _zz_dataOut_payload_0_1957;
    _zz_dataOut_payload_0_1974 <= _zz_dataOut_payload_0_1958;
    _zz_dataOut_payload_0_1975 <= _zz_dataOut_payload_0_1959;
    _zz_dataOut_payload_0_1976 <= _zz_dataOut_payload_0_1968;
    _zz_dataOut_payload_0_1977 <= _zz_dataOut_payload_0_1969;
    _zz_dataOut_payload_0_1978 <= _zz_dataOut_payload_0_1970;
    _zz_dataOut_payload_0_1979 <= _zz_dataOut_payload_0_1971;
    _zz_dataOut_payload_0_2000 <= (_zz_dataOut_payload_0_1998 ? _zz_dataOut_payload_0_1993 : _zz_dataOut_payload_0_1996);
    _zz_dataOut_payload_0_2001 <= (_zz_dataOut_payload_0_1998 ? _zz_dataOut_payload_0_1996 : _zz_dataOut_payload_0_1993);
    _zz_dataOut_payload_0_2002 <= (_zz_dataOut_payload_0_1999 ? _zz_dataOut_payload_0_1994 : _zz_dataOut_payload_0_1997);
    _zz_dataOut_payload_0_2003 <= (_zz_dataOut_payload_0_1999 ? _zz_dataOut_payload_0_1997 : _zz_dataOut_payload_0_1994);
    _zz_dataOut_payload_0_2012 <= (_zz_dataOut_payload_0_2010 ? _zz_dataOut_payload_0_2005 : _zz_dataOut_payload_0_2008);
    _zz_dataOut_payload_0_2013 <= (_zz_dataOut_payload_0_2010 ? _zz_dataOut_payload_0_2008 : _zz_dataOut_payload_0_2005);
    _zz_dataOut_payload_0_2014 <= (_zz_dataOut_payload_0_2011 ? _zz_dataOut_payload_0_2006 : _zz_dataOut_payload_0_2009);
    _zz_dataOut_payload_0_2015 <= (_zz_dataOut_payload_0_2011 ? _zz_dataOut_payload_0_2009 : _zz_dataOut_payload_0_2006);
    _zz_dataOut_payload_0_2016 <= _zz_dataOut_payload_0_2000;
    _zz_dataOut_payload_0_2017 <= _zz_dataOut_payload_0_2001;
    _zz_dataOut_payload_0_2018 <= _zz_dataOut_payload_0_2002;
    _zz_dataOut_payload_0_2019 <= _zz_dataOut_payload_0_2003;
    _zz_dataOut_payload_0_2020 <= _zz_dataOut_payload_0_2012;
    _zz_dataOut_payload_0_2021 <= _zz_dataOut_payload_0_2013;
    _zz_dataOut_payload_0_2022 <= _zz_dataOut_payload_0_2014;
    _zz_dataOut_payload_0_2023 <= _zz_dataOut_payload_0_2015;
    _zz_dataOut_payload_0_2044 <= (_zz_dataOut_payload_0_2042 ? _zz_dataOut_payload_0_2037 : _zz_dataOut_payload_0_2040);
    _zz_dataOut_payload_0_2045 <= (_zz_dataOut_payload_0_2042 ? _zz_dataOut_payload_0_2040 : _zz_dataOut_payload_0_2037);
    _zz_dataOut_payload_0_2046 <= (_zz_dataOut_payload_0_2043 ? _zz_dataOut_payload_0_2038 : _zz_dataOut_payload_0_2041);
    _zz_dataOut_payload_0_2047 <= (_zz_dataOut_payload_0_2043 ? _zz_dataOut_payload_0_2041 : _zz_dataOut_payload_0_2038);
    _zz_dataOut_payload_0_2056 <= (_zz_dataOut_payload_0_2054 ? _zz_dataOut_payload_0_2049 : _zz_dataOut_payload_0_2052);
    _zz_dataOut_payload_0_2057 <= (_zz_dataOut_payload_0_2054 ? _zz_dataOut_payload_0_2052 : _zz_dataOut_payload_0_2049);
    _zz_dataOut_payload_0_2058 <= (_zz_dataOut_payload_0_2055 ? _zz_dataOut_payload_0_2050 : _zz_dataOut_payload_0_2053);
    _zz_dataOut_payload_0_2059 <= (_zz_dataOut_payload_0_2055 ? _zz_dataOut_payload_0_2053 : _zz_dataOut_payload_0_2050);
    _zz_dataOut_payload_0_2060 <= _zz_dataOut_payload_0_2044;
    _zz_dataOut_payload_0_2061 <= _zz_dataOut_payload_0_2045;
    _zz_dataOut_payload_0_2062 <= _zz_dataOut_payload_0_2046;
    _zz_dataOut_payload_0_2063 <= _zz_dataOut_payload_0_2047;
    _zz_dataOut_payload_0_2064 <= _zz_dataOut_payload_0_2056;
    _zz_dataOut_payload_0_2065 <= _zz_dataOut_payload_0_2057;
    _zz_dataOut_payload_0_2066 <= _zz_dataOut_payload_0_2058;
    _zz_dataOut_payload_0_2067 <= _zz_dataOut_payload_0_2059;
    _zz_dataOut_payload_0_2088 <= (_zz_dataOut_payload_0_2086 ? _zz_dataOut_payload_0_2081 : _zz_dataOut_payload_0_2084);
    _zz_dataOut_payload_0_2089 <= (_zz_dataOut_payload_0_2086 ? _zz_dataOut_payload_0_2084 : _zz_dataOut_payload_0_2081);
    _zz_dataOut_payload_0_2090 <= (_zz_dataOut_payload_0_2087 ? _zz_dataOut_payload_0_2082 : _zz_dataOut_payload_0_2085);
    _zz_dataOut_payload_0_2091 <= (_zz_dataOut_payload_0_2087 ? _zz_dataOut_payload_0_2085 : _zz_dataOut_payload_0_2082);
    _zz_dataOut_payload_0_2100 <= (_zz_dataOut_payload_0_2098 ? _zz_dataOut_payload_0_2093 : _zz_dataOut_payload_0_2096);
    _zz_dataOut_payload_0_2101 <= (_zz_dataOut_payload_0_2098 ? _zz_dataOut_payload_0_2096 : _zz_dataOut_payload_0_2093);
    _zz_dataOut_payload_0_2102 <= (_zz_dataOut_payload_0_2099 ? _zz_dataOut_payload_0_2094 : _zz_dataOut_payload_0_2097);
    _zz_dataOut_payload_0_2103 <= (_zz_dataOut_payload_0_2099 ? _zz_dataOut_payload_0_2097 : _zz_dataOut_payload_0_2094);
    _zz_dataOut_payload_0_2104 <= _zz_dataOut_payload_0_2088;
    _zz_dataOut_payload_0_2105 <= _zz_dataOut_payload_0_2089;
    _zz_dataOut_payload_0_2106 <= _zz_dataOut_payload_0_2090;
    _zz_dataOut_payload_0_2107 <= _zz_dataOut_payload_0_2091;
    _zz_dataOut_payload_0_2108 <= _zz_dataOut_payload_0_2100;
    _zz_dataOut_payload_0_2109 <= _zz_dataOut_payload_0_2101;
    _zz_dataOut_payload_0_2110 <= _zz_dataOut_payload_0_2102;
    _zz_dataOut_payload_0_2111 <= _zz_dataOut_payload_0_2103;
    _zz_dataOut_payload_0_2132 <= (_zz_dataOut_payload_0_2130 ? _zz_dataOut_payload_0_2125 : _zz_dataOut_payload_0_2128);
    _zz_dataOut_payload_0_2133 <= (_zz_dataOut_payload_0_2130 ? _zz_dataOut_payload_0_2128 : _zz_dataOut_payload_0_2125);
    _zz_dataOut_payload_0_2134 <= (_zz_dataOut_payload_0_2131 ? _zz_dataOut_payload_0_2126 : _zz_dataOut_payload_0_2129);
    _zz_dataOut_payload_0_2135 <= (_zz_dataOut_payload_0_2131 ? _zz_dataOut_payload_0_2129 : _zz_dataOut_payload_0_2126);
    _zz_dataOut_payload_0_2144 <= (_zz_dataOut_payload_0_2142 ? _zz_dataOut_payload_0_2137 : _zz_dataOut_payload_0_2140);
    _zz_dataOut_payload_0_2145 <= (_zz_dataOut_payload_0_2142 ? _zz_dataOut_payload_0_2140 : _zz_dataOut_payload_0_2137);
    _zz_dataOut_payload_0_2146 <= (_zz_dataOut_payload_0_2143 ? _zz_dataOut_payload_0_2138 : _zz_dataOut_payload_0_2141);
    _zz_dataOut_payload_0_2147 <= (_zz_dataOut_payload_0_2143 ? _zz_dataOut_payload_0_2141 : _zz_dataOut_payload_0_2138);
    _zz_dataOut_payload_0_2148 <= _zz_dataOut_payload_0_2132;
    _zz_dataOut_payload_0_2149 <= _zz_dataOut_payload_0_2133;
    _zz_dataOut_payload_0_2150 <= _zz_dataOut_payload_0_2134;
    _zz_dataOut_payload_0_2151 <= _zz_dataOut_payload_0_2135;
    _zz_dataOut_payload_0_2152 <= _zz_dataOut_payload_0_2144;
    _zz_dataOut_payload_0_2153 <= _zz_dataOut_payload_0_2145;
    _zz_dataOut_payload_0_2154 <= _zz_dataOut_payload_0_2146;
    _zz_dataOut_payload_0_2155 <= _zz_dataOut_payload_0_2147;
    _zz_dataOut_payload_0_2176 <= (_zz_dataOut_payload_0_2174 ? _zz_dataOut_payload_0_2169 : _zz_dataOut_payload_0_2172);
    _zz_dataOut_payload_0_2177 <= (_zz_dataOut_payload_0_2174 ? _zz_dataOut_payload_0_2172 : _zz_dataOut_payload_0_2169);
    _zz_dataOut_payload_0_2178 <= (_zz_dataOut_payload_0_2175 ? _zz_dataOut_payload_0_2170 : _zz_dataOut_payload_0_2173);
    _zz_dataOut_payload_0_2179 <= (_zz_dataOut_payload_0_2175 ? _zz_dataOut_payload_0_2173 : _zz_dataOut_payload_0_2170);
    _zz_dataOut_payload_0_2188 <= (_zz_dataOut_payload_0_2186 ? _zz_dataOut_payload_0_2181 : _zz_dataOut_payload_0_2184);
    _zz_dataOut_payload_0_2189 <= (_zz_dataOut_payload_0_2186 ? _zz_dataOut_payload_0_2184 : _zz_dataOut_payload_0_2181);
    _zz_dataOut_payload_0_2190 <= (_zz_dataOut_payload_0_2187 ? _zz_dataOut_payload_0_2182 : _zz_dataOut_payload_0_2185);
    _zz_dataOut_payload_0_2191 <= (_zz_dataOut_payload_0_2187 ? _zz_dataOut_payload_0_2185 : _zz_dataOut_payload_0_2182);
    _zz_dataOut_payload_0_2192 <= _zz_dataOut_payload_0_2176;
    _zz_dataOut_payload_0_2193 <= _zz_dataOut_payload_0_2177;
    _zz_dataOut_payload_0_2194 <= _zz_dataOut_payload_0_2178;
    _zz_dataOut_payload_0_2195 <= _zz_dataOut_payload_0_2179;
    _zz_dataOut_payload_0_2196 <= _zz_dataOut_payload_0_2188;
    _zz_dataOut_payload_0_2197 <= _zz_dataOut_payload_0_2189;
    _zz_dataOut_payload_0_2198 <= _zz_dataOut_payload_0_2190;
    _zz_dataOut_payload_0_2199 <= _zz_dataOut_payload_0_2191;
    _zz_dataOut_payload_0_2220 <= (_zz_dataOut_payload_0_2218 ? _zz_dataOut_payload_0_2213 : _zz_dataOut_payload_0_2216);
    _zz_dataOut_payload_0_2221 <= (_zz_dataOut_payload_0_2218 ? _zz_dataOut_payload_0_2216 : _zz_dataOut_payload_0_2213);
    _zz_dataOut_payload_0_2222 <= (_zz_dataOut_payload_0_2219 ? _zz_dataOut_payload_0_2214 : _zz_dataOut_payload_0_2217);
    _zz_dataOut_payload_0_2223 <= (_zz_dataOut_payload_0_2219 ? _zz_dataOut_payload_0_2217 : _zz_dataOut_payload_0_2214);
    _zz_dataOut_payload_0_2232 <= (_zz_dataOut_payload_0_2230 ? _zz_dataOut_payload_0_2225 : _zz_dataOut_payload_0_2228);
    _zz_dataOut_payload_0_2233 <= (_zz_dataOut_payload_0_2230 ? _zz_dataOut_payload_0_2228 : _zz_dataOut_payload_0_2225);
    _zz_dataOut_payload_0_2234 <= (_zz_dataOut_payload_0_2231 ? _zz_dataOut_payload_0_2226 : _zz_dataOut_payload_0_2229);
    _zz_dataOut_payload_0_2235 <= (_zz_dataOut_payload_0_2231 ? _zz_dataOut_payload_0_2229 : _zz_dataOut_payload_0_2226);
    _zz_dataOut_payload_0_2236 <= _zz_dataOut_payload_0_2220;
    _zz_dataOut_payload_0_2237 <= _zz_dataOut_payload_0_2221;
    _zz_dataOut_payload_0_2238 <= _zz_dataOut_payload_0_2222;
    _zz_dataOut_payload_0_2239 <= _zz_dataOut_payload_0_2223;
    _zz_dataOut_payload_0_2240 <= _zz_dataOut_payload_0_2232;
    _zz_dataOut_payload_0_2241 <= _zz_dataOut_payload_0_2233;
    _zz_dataOut_payload_0_2242 <= _zz_dataOut_payload_0_2234;
    _zz_dataOut_payload_0_2243 <= _zz_dataOut_payload_0_2235;
    _zz_dataOut_payload_0_2264 <= (_zz_dataOut_payload_0_2262 ? _zz_dataOut_payload_0_2257 : _zz_dataOut_payload_0_2260);
    _zz_dataOut_payload_0_2265 <= (_zz_dataOut_payload_0_2262 ? _zz_dataOut_payload_0_2260 : _zz_dataOut_payload_0_2257);
    _zz_dataOut_payload_0_2266 <= (_zz_dataOut_payload_0_2263 ? _zz_dataOut_payload_0_2258 : _zz_dataOut_payload_0_2261);
    _zz_dataOut_payload_0_2267 <= (_zz_dataOut_payload_0_2263 ? _zz_dataOut_payload_0_2261 : _zz_dataOut_payload_0_2258);
    _zz_dataOut_payload_0_2276 <= (_zz_dataOut_payload_0_2274 ? _zz_dataOut_payload_0_2269 : _zz_dataOut_payload_0_2272);
    _zz_dataOut_payload_0_2277 <= (_zz_dataOut_payload_0_2274 ? _zz_dataOut_payload_0_2272 : _zz_dataOut_payload_0_2269);
    _zz_dataOut_payload_0_2278 <= (_zz_dataOut_payload_0_2275 ? _zz_dataOut_payload_0_2270 : _zz_dataOut_payload_0_2273);
    _zz_dataOut_payload_0_2279 <= (_zz_dataOut_payload_0_2275 ? _zz_dataOut_payload_0_2273 : _zz_dataOut_payload_0_2270);
    _zz_dataOut_payload_0_2280 <= _zz_dataOut_payload_0_2264;
    _zz_dataOut_payload_0_2281 <= _zz_dataOut_payload_0_2265;
    _zz_dataOut_payload_0_2282 <= _zz_dataOut_payload_0_2266;
    _zz_dataOut_payload_0_2283 <= _zz_dataOut_payload_0_2267;
    _zz_dataOut_payload_0_2284 <= _zz_dataOut_payload_0_2276;
    _zz_dataOut_payload_0_2285 <= _zz_dataOut_payload_0_2277;
    _zz_dataOut_payload_0_2286 <= _zz_dataOut_payload_0_2278;
    _zz_dataOut_payload_0_2287 <= _zz_dataOut_payload_0_2279;
    _zz_dataOut_payload_0_2308 <= (_zz_dataOut_payload_0_2306 ? _zz_dataOut_payload_0_2301 : _zz_dataOut_payload_0_2304);
    _zz_dataOut_payload_0_2309 <= (_zz_dataOut_payload_0_2306 ? _zz_dataOut_payload_0_2304 : _zz_dataOut_payload_0_2301);
    _zz_dataOut_payload_0_2310 <= (_zz_dataOut_payload_0_2307 ? _zz_dataOut_payload_0_2302 : _zz_dataOut_payload_0_2305);
    _zz_dataOut_payload_0_2311 <= (_zz_dataOut_payload_0_2307 ? _zz_dataOut_payload_0_2305 : _zz_dataOut_payload_0_2302);
    _zz_dataOut_payload_0_2320 <= (_zz_dataOut_payload_0_2318 ? _zz_dataOut_payload_0_2313 : _zz_dataOut_payload_0_2316);
    _zz_dataOut_payload_0_2321 <= (_zz_dataOut_payload_0_2318 ? _zz_dataOut_payload_0_2316 : _zz_dataOut_payload_0_2313);
    _zz_dataOut_payload_0_2322 <= (_zz_dataOut_payload_0_2319 ? _zz_dataOut_payload_0_2314 : _zz_dataOut_payload_0_2317);
    _zz_dataOut_payload_0_2323 <= (_zz_dataOut_payload_0_2319 ? _zz_dataOut_payload_0_2317 : _zz_dataOut_payload_0_2314);
    _zz_dataOut_payload_0_2324 <= _zz_dataOut_payload_0_2308;
    _zz_dataOut_payload_0_2325 <= _zz_dataOut_payload_0_2309;
    _zz_dataOut_payload_0_2326 <= _zz_dataOut_payload_0_2310;
    _zz_dataOut_payload_0_2327 <= _zz_dataOut_payload_0_2311;
    _zz_dataOut_payload_0_2328 <= _zz_dataOut_payload_0_2320;
    _zz_dataOut_payload_0_2329 <= _zz_dataOut_payload_0_2321;
    _zz_dataOut_payload_0_2330 <= _zz_dataOut_payload_0_2322;
    _zz_dataOut_payload_0_2331 <= _zz_dataOut_payload_0_2323;
    _zz_dataOut_payload_0_2352 <= (_zz_dataOut_payload_0_2350 ? _zz_dataOut_payload_0_2345 : _zz_dataOut_payload_0_2348);
    _zz_dataOut_payload_0_2353 <= (_zz_dataOut_payload_0_2350 ? _zz_dataOut_payload_0_2348 : _zz_dataOut_payload_0_2345);
    _zz_dataOut_payload_0_2354 <= (_zz_dataOut_payload_0_2351 ? _zz_dataOut_payload_0_2346 : _zz_dataOut_payload_0_2349);
    _zz_dataOut_payload_0_2355 <= (_zz_dataOut_payload_0_2351 ? _zz_dataOut_payload_0_2349 : _zz_dataOut_payload_0_2346);
    _zz_dataOut_payload_0_2364 <= (_zz_dataOut_payload_0_2362 ? _zz_dataOut_payload_0_2357 : _zz_dataOut_payload_0_2360);
    _zz_dataOut_payload_0_2365 <= (_zz_dataOut_payload_0_2362 ? _zz_dataOut_payload_0_2360 : _zz_dataOut_payload_0_2357);
    _zz_dataOut_payload_0_2366 <= (_zz_dataOut_payload_0_2363 ? _zz_dataOut_payload_0_2358 : _zz_dataOut_payload_0_2361);
    _zz_dataOut_payload_0_2367 <= (_zz_dataOut_payload_0_2363 ? _zz_dataOut_payload_0_2361 : _zz_dataOut_payload_0_2358);
    _zz_dataOut_payload_0_2368 <= _zz_dataOut_payload_0_2352;
    _zz_dataOut_payload_0_2369 <= _zz_dataOut_payload_0_2353;
    _zz_dataOut_payload_0_2370 <= _zz_dataOut_payload_0_2354;
    _zz_dataOut_payload_0_2371 <= _zz_dataOut_payload_0_2355;
    _zz_dataOut_payload_0_2372 <= _zz_dataOut_payload_0_2364;
    _zz_dataOut_payload_0_2373 <= _zz_dataOut_payload_0_2365;
    _zz_dataOut_payload_0_2374 <= _zz_dataOut_payload_0_2366;
    _zz_dataOut_payload_0_2375 <= _zz_dataOut_payload_0_2367;
    _zz_dataOut_payload_0_2396 <= (_zz_dataOut_payload_0_2394 ? _zz_dataOut_payload_0_2389 : _zz_dataOut_payload_0_2392);
    _zz_dataOut_payload_0_2397 <= (_zz_dataOut_payload_0_2394 ? _zz_dataOut_payload_0_2392 : _zz_dataOut_payload_0_2389);
    _zz_dataOut_payload_0_2398 <= (_zz_dataOut_payload_0_2395 ? _zz_dataOut_payload_0_2390 : _zz_dataOut_payload_0_2393);
    _zz_dataOut_payload_0_2399 <= (_zz_dataOut_payload_0_2395 ? _zz_dataOut_payload_0_2393 : _zz_dataOut_payload_0_2390);
    _zz_dataOut_payload_0_2408 <= (_zz_dataOut_payload_0_2406 ? _zz_dataOut_payload_0_2401 : _zz_dataOut_payload_0_2404);
    _zz_dataOut_payload_0_2409 <= (_zz_dataOut_payload_0_2406 ? _zz_dataOut_payload_0_2404 : _zz_dataOut_payload_0_2401);
    _zz_dataOut_payload_0_2410 <= (_zz_dataOut_payload_0_2407 ? _zz_dataOut_payload_0_2402 : _zz_dataOut_payload_0_2405);
    _zz_dataOut_payload_0_2411 <= (_zz_dataOut_payload_0_2407 ? _zz_dataOut_payload_0_2405 : _zz_dataOut_payload_0_2402);
    _zz_dataOut_payload_0_2412 <= _zz_dataOut_payload_0_2396;
    _zz_dataOut_payload_0_2413 <= _zz_dataOut_payload_0_2397;
    _zz_dataOut_payload_0_2414 <= _zz_dataOut_payload_0_2398;
    _zz_dataOut_payload_0_2415 <= _zz_dataOut_payload_0_2399;
    _zz_dataOut_payload_0_2416 <= _zz_dataOut_payload_0_2408;
    _zz_dataOut_payload_0_2417 <= _zz_dataOut_payload_0_2409;
    _zz_dataOut_payload_0_2418 <= _zz_dataOut_payload_0_2410;
    _zz_dataOut_payload_0_2419 <= _zz_dataOut_payload_0_2411;
    _zz_dataOut_payload_0_2440 <= (_zz_dataOut_payload_0_2438 ? _zz_dataOut_payload_0_2433 : _zz_dataOut_payload_0_2436);
    _zz_dataOut_payload_0_2441 <= (_zz_dataOut_payload_0_2438 ? _zz_dataOut_payload_0_2436 : _zz_dataOut_payload_0_2433);
    _zz_dataOut_payload_0_2442 <= (_zz_dataOut_payload_0_2439 ? _zz_dataOut_payload_0_2434 : _zz_dataOut_payload_0_2437);
    _zz_dataOut_payload_0_2443 <= (_zz_dataOut_payload_0_2439 ? _zz_dataOut_payload_0_2437 : _zz_dataOut_payload_0_2434);
    _zz_dataOut_payload_0_2452 <= (_zz_dataOut_payload_0_2450 ? _zz_dataOut_payload_0_2445 : _zz_dataOut_payload_0_2448);
    _zz_dataOut_payload_0_2453 <= (_zz_dataOut_payload_0_2450 ? _zz_dataOut_payload_0_2448 : _zz_dataOut_payload_0_2445);
    _zz_dataOut_payload_0_2454 <= (_zz_dataOut_payload_0_2451 ? _zz_dataOut_payload_0_2446 : _zz_dataOut_payload_0_2449);
    _zz_dataOut_payload_0_2455 <= (_zz_dataOut_payload_0_2451 ? _zz_dataOut_payload_0_2449 : _zz_dataOut_payload_0_2446);
    _zz_dataOut_payload_0_2456 <= _zz_dataOut_payload_0_2440;
    _zz_dataOut_payload_0_2457 <= _zz_dataOut_payload_0_2441;
    _zz_dataOut_payload_0_2458 <= _zz_dataOut_payload_0_2442;
    _zz_dataOut_payload_0_2459 <= _zz_dataOut_payload_0_2443;
    _zz_dataOut_payload_0_2460 <= _zz_dataOut_payload_0_2452;
    _zz_dataOut_payload_0_2461 <= _zz_dataOut_payload_0_2453;
    _zz_dataOut_payload_0_2462 <= _zz_dataOut_payload_0_2454;
    _zz_dataOut_payload_0_2463 <= _zz_dataOut_payload_0_2455;
    _zz_dataOut_payload_0_2484 <= (_zz_dataOut_payload_0_2482 ? _zz_dataOut_payload_0_2477 : _zz_dataOut_payload_0_2480);
    _zz_dataOut_payload_0_2485 <= (_zz_dataOut_payload_0_2482 ? _zz_dataOut_payload_0_2480 : _zz_dataOut_payload_0_2477);
    _zz_dataOut_payload_0_2486 <= (_zz_dataOut_payload_0_2483 ? _zz_dataOut_payload_0_2478 : _zz_dataOut_payload_0_2481);
    _zz_dataOut_payload_0_2487 <= (_zz_dataOut_payload_0_2483 ? _zz_dataOut_payload_0_2481 : _zz_dataOut_payload_0_2478);
    _zz_dataOut_payload_0_2496 <= (_zz_dataOut_payload_0_2494 ? _zz_dataOut_payload_0_2489 : _zz_dataOut_payload_0_2492);
    _zz_dataOut_payload_0_2497 <= (_zz_dataOut_payload_0_2494 ? _zz_dataOut_payload_0_2492 : _zz_dataOut_payload_0_2489);
    _zz_dataOut_payload_0_2498 <= (_zz_dataOut_payload_0_2495 ? _zz_dataOut_payload_0_2490 : _zz_dataOut_payload_0_2493);
    _zz_dataOut_payload_0_2499 <= (_zz_dataOut_payload_0_2495 ? _zz_dataOut_payload_0_2493 : _zz_dataOut_payload_0_2490);
    _zz_dataOut_payload_0_2500 <= _zz_dataOut_payload_0_2484;
    _zz_dataOut_payload_0_2501 <= _zz_dataOut_payload_0_2485;
    _zz_dataOut_payload_0_2502 <= _zz_dataOut_payload_0_2486;
    _zz_dataOut_payload_0_2503 <= _zz_dataOut_payload_0_2487;
    _zz_dataOut_payload_0_2504 <= _zz_dataOut_payload_0_2496;
    _zz_dataOut_payload_0_2505 <= _zz_dataOut_payload_0_2497;
    _zz_dataOut_payload_0_2506 <= _zz_dataOut_payload_0_2498;
    _zz_dataOut_payload_0_2507 <= _zz_dataOut_payload_0_2499;
    _zz_dataOut_payload_0_2528 <= (_zz_dataOut_payload_0_2526 ? _zz_dataOut_payload_0_2521 : _zz_dataOut_payload_0_2524);
    _zz_dataOut_payload_0_2529 <= (_zz_dataOut_payload_0_2526 ? _zz_dataOut_payload_0_2524 : _zz_dataOut_payload_0_2521);
    _zz_dataOut_payload_0_2530 <= (_zz_dataOut_payload_0_2527 ? _zz_dataOut_payload_0_2522 : _zz_dataOut_payload_0_2525);
    _zz_dataOut_payload_0_2531 <= (_zz_dataOut_payload_0_2527 ? _zz_dataOut_payload_0_2525 : _zz_dataOut_payload_0_2522);
    _zz_dataOut_payload_0_2540 <= (_zz_dataOut_payload_0_2538 ? _zz_dataOut_payload_0_2533 : _zz_dataOut_payload_0_2536);
    _zz_dataOut_payload_0_2541 <= (_zz_dataOut_payload_0_2538 ? _zz_dataOut_payload_0_2536 : _zz_dataOut_payload_0_2533);
    _zz_dataOut_payload_0_2542 <= (_zz_dataOut_payload_0_2539 ? _zz_dataOut_payload_0_2534 : _zz_dataOut_payload_0_2537);
    _zz_dataOut_payload_0_2543 <= (_zz_dataOut_payload_0_2539 ? _zz_dataOut_payload_0_2537 : _zz_dataOut_payload_0_2534);
    _zz_dataOut_payload_0_2544 <= _zz_dataOut_payload_0_2528;
    _zz_dataOut_payload_0_2545 <= _zz_dataOut_payload_0_2529;
    _zz_dataOut_payload_0_2546 <= _zz_dataOut_payload_0_2530;
    _zz_dataOut_payload_0_2547 <= _zz_dataOut_payload_0_2531;
    _zz_dataOut_payload_0_2548 <= _zz_dataOut_payload_0_2540;
    _zz_dataOut_payload_0_2549 <= _zz_dataOut_payload_0_2541;
    _zz_dataOut_payload_0_2550 <= _zz_dataOut_payload_0_2542;
    _zz_dataOut_payload_0_2551 <= _zz_dataOut_payload_0_2543;
    _zz_dataOut_payload_0_2572 <= (_zz_dataOut_payload_0_2570 ? _zz_dataOut_payload_0_2565 : _zz_dataOut_payload_0_2568);
    _zz_dataOut_payload_0_2573 <= (_zz_dataOut_payload_0_2570 ? _zz_dataOut_payload_0_2568 : _zz_dataOut_payload_0_2565);
    _zz_dataOut_payload_0_2574 <= (_zz_dataOut_payload_0_2571 ? _zz_dataOut_payload_0_2566 : _zz_dataOut_payload_0_2569);
    _zz_dataOut_payload_0_2575 <= (_zz_dataOut_payload_0_2571 ? _zz_dataOut_payload_0_2569 : _zz_dataOut_payload_0_2566);
    _zz_dataOut_payload_0_2584 <= (_zz_dataOut_payload_0_2582 ? _zz_dataOut_payload_0_2577 : _zz_dataOut_payload_0_2580);
    _zz_dataOut_payload_0_2585 <= (_zz_dataOut_payload_0_2582 ? _zz_dataOut_payload_0_2580 : _zz_dataOut_payload_0_2577);
    _zz_dataOut_payload_0_2586 <= (_zz_dataOut_payload_0_2583 ? _zz_dataOut_payload_0_2578 : _zz_dataOut_payload_0_2581);
    _zz_dataOut_payload_0_2587 <= (_zz_dataOut_payload_0_2583 ? _zz_dataOut_payload_0_2581 : _zz_dataOut_payload_0_2578);
    _zz_dataOut_payload_0_2588 <= _zz_dataOut_payload_0_2572;
    _zz_dataOut_payload_0_2589 <= _zz_dataOut_payload_0_2573;
    _zz_dataOut_payload_0_2590 <= _zz_dataOut_payload_0_2574;
    _zz_dataOut_payload_0_2591 <= _zz_dataOut_payload_0_2575;
    _zz_dataOut_payload_0_2592 <= _zz_dataOut_payload_0_2584;
    _zz_dataOut_payload_0_2593 <= _zz_dataOut_payload_0_2585;
    _zz_dataOut_payload_0_2594 <= _zz_dataOut_payload_0_2586;
    _zz_dataOut_payload_0_2595 <= _zz_dataOut_payload_0_2587;
    _zz_dataOut_payload_0_2616 <= (_zz_dataOut_payload_0_2614 ? _zz_dataOut_payload_0_2609 : _zz_dataOut_payload_0_2612);
    _zz_dataOut_payload_0_2617 <= (_zz_dataOut_payload_0_2614 ? _zz_dataOut_payload_0_2612 : _zz_dataOut_payload_0_2609);
    _zz_dataOut_payload_0_2618 <= (_zz_dataOut_payload_0_2615 ? _zz_dataOut_payload_0_2610 : _zz_dataOut_payload_0_2613);
    _zz_dataOut_payload_0_2619 <= (_zz_dataOut_payload_0_2615 ? _zz_dataOut_payload_0_2613 : _zz_dataOut_payload_0_2610);
    _zz_dataOut_payload_0_2628 <= (_zz_dataOut_payload_0_2626 ? _zz_dataOut_payload_0_2621 : _zz_dataOut_payload_0_2624);
    _zz_dataOut_payload_0_2629 <= (_zz_dataOut_payload_0_2626 ? _zz_dataOut_payload_0_2624 : _zz_dataOut_payload_0_2621);
    _zz_dataOut_payload_0_2630 <= (_zz_dataOut_payload_0_2627 ? _zz_dataOut_payload_0_2622 : _zz_dataOut_payload_0_2625);
    _zz_dataOut_payload_0_2631 <= (_zz_dataOut_payload_0_2627 ? _zz_dataOut_payload_0_2625 : _zz_dataOut_payload_0_2622);
    _zz_dataOut_payload_0_2632 <= _zz_dataOut_payload_0_2616;
    _zz_dataOut_payload_0_2633 <= _zz_dataOut_payload_0_2617;
    _zz_dataOut_payload_0_2634 <= _zz_dataOut_payload_0_2618;
    _zz_dataOut_payload_0_2635 <= _zz_dataOut_payload_0_2619;
    _zz_dataOut_payload_0_2636 <= _zz_dataOut_payload_0_2628;
    _zz_dataOut_payload_0_2637 <= _zz_dataOut_payload_0_2629;
    _zz_dataOut_payload_0_2638 <= _zz_dataOut_payload_0_2630;
    _zz_dataOut_payload_0_2639 <= _zz_dataOut_payload_0_2631;
    _zz_dataOut_payload_0_2660 <= (_zz_dataOut_payload_0_2658 ? _zz_dataOut_payload_0_2653 : _zz_dataOut_payload_0_2656);
    _zz_dataOut_payload_0_2661 <= (_zz_dataOut_payload_0_2658 ? _zz_dataOut_payload_0_2656 : _zz_dataOut_payload_0_2653);
    _zz_dataOut_payload_0_2662 <= (_zz_dataOut_payload_0_2659 ? _zz_dataOut_payload_0_2654 : _zz_dataOut_payload_0_2657);
    _zz_dataOut_payload_0_2663 <= (_zz_dataOut_payload_0_2659 ? _zz_dataOut_payload_0_2657 : _zz_dataOut_payload_0_2654);
    _zz_dataOut_payload_0_2672 <= (_zz_dataOut_payload_0_2670 ? _zz_dataOut_payload_0_2665 : _zz_dataOut_payload_0_2668);
    _zz_dataOut_payload_0_2673 <= (_zz_dataOut_payload_0_2670 ? _zz_dataOut_payload_0_2668 : _zz_dataOut_payload_0_2665);
    _zz_dataOut_payload_0_2674 <= (_zz_dataOut_payload_0_2671 ? _zz_dataOut_payload_0_2666 : _zz_dataOut_payload_0_2669);
    _zz_dataOut_payload_0_2675 <= (_zz_dataOut_payload_0_2671 ? _zz_dataOut_payload_0_2669 : _zz_dataOut_payload_0_2666);
    _zz_dataOut_payload_0_2676 <= _zz_dataOut_payload_0_2660;
    _zz_dataOut_payload_0_2677 <= _zz_dataOut_payload_0_2661;
    _zz_dataOut_payload_0_2678 <= _zz_dataOut_payload_0_2662;
    _zz_dataOut_payload_0_2679 <= _zz_dataOut_payload_0_2663;
    _zz_dataOut_payload_0_2680 <= _zz_dataOut_payload_0_2672;
    _zz_dataOut_payload_0_2681 <= _zz_dataOut_payload_0_2673;
    _zz_dataOut_payload_0_2682 <= _zz_dataOut_payload_0_2674;
    _zz_dataOut_payload_0_2683 <= _zz_dataOut_payload_0_2675;
    _zz_dataOut_payload_0_2704 <= (_zz_dataOut_payload_0_2702 ? _zz_dataOut_payload_0_2697 : _zz_dataOut_payload_0_2700);
    _zz_dataOut_payload_0_2705 <= (_zz_dataOut_payload_0_2702 ? _zz_dataOut_payload_0_2700 : _zz_dataOut_payload_0_2697);
    _zz_dataOut_payload_0_2706 <= (_zz_dataOut_payload_0_2703 ? _zz_dataOut_payload_0_2698 : _zz_dataOut_payload_0_2701);
    _zz_dataOut_payload_0_2707 <= (_zz_dataOut_payload_0_2703 ? _zz_dataOut_payload_0_2701 : _zz_dataOut_payload_0_2698);
    _zz_dataOut_payload_0_2716 <= (_zz_dataOut_payload_0_2714 ? _zz_dataOut_payload_0_2709 : _zz_dataOut_payload_0_2712);
    _zz_dataOut_payload_0_2717 <= (_zz_dataOut_payload_0_2714 ? _zz_dataOut_payload_0_2712 : _zz_dataOut_payload_0_2709);
    _zz_dataOut_payload_0_2718 <= (_zz_dataOut_payload_0_2715 ? _zz_dataOut_payload_0_2710 : _zz_dataOut_payload_0_2713);
    _zz_dataOut_payload_0_2719 <= (_zz_dataOut_payload_0_2715 ? _zz_dataOut_payload_0_2713 : _zz_dataOut_payload_0_2710);
    _zz_dataOut_payload_0_2720 <= _zz_dataOut_payload_0_2704;
    _zz_dataOut_payload_0_2721 <= _zz_dataOut_payload_0_2705;
    _zz_dataOut_payload_0_2722 <= _zz_dataOut_payload_0_2706;
    _zz_dataOut_payload_0_2723 <= _zz_dataOut_payload_0_2707;
    _zz_dataOut_payload_0_2724 <= _zz_dataOut_payload_0_2716;
    _zz_dataOut_payload_0_2725 <= _zz_dataOut_payload_0_2717;
    _zz_dataOut_payload_0_2726 <= _zz_dataOut_payload_0_2718;
    _zz_dataOut_payload_0_2727 <= _zz_dataOut_payload_0_2719;
    _zz_dataOut_payload_0_2748 <= (_zz_dataOut_payload_0_2746 ? _zz_dataOut_payload_0_2741 : _zz_dataOut_payload_0_2744);
    _zz_dataOut_payload_0_2749 <= (_zz_dataOut_payload_0_2746 ? _zz_dataOut_payload_0_2744 : _zz_dataOut_payload_0_2741);
    _zz_dataOut_payload_0_2750 <= (_zz_dataOut_payload_0_2747 ? _zz_dataOut_payload_0_2742 : _zz_dataOut_payload_0_2745);
    _zz_dataOut_payload_0_2751 <= (_zz_dataOut_payload_0_2747 ? _zz_dataOut_payload_0_2745 : _zz_dataOut_payload_0_2742);
    _zz_dataOut_payload_0_2760 <= (_zz_dataOut_payload_0_2758 ? _zz_dataOut_payload_0_2753 : _zz_dataOut_payload_0_2756);
    _zz_dataOut_payload_0_2761 <= (_zz_dataOut_payload_0_2758 ? _zz_dataOut_payload_0_2756 : _zz_dataOut_payload_0_2753);
    _zz_dataOut_payload_0_2762 <= (_zz_dataOut_payload_0_2759 ? _zz_dataOut_payload_0_2754 : _zz_dataOut_payload_0_2757);
    _zz_dataOut_payload_0_2763 <= (_zz_dataOut_payload_0_2759 ? _zz_dataOut_payload_0_2757 : _zz_dataOut_payload_0_2754);
    _zz_dataOut_payload_0_2764 <= _zz_dataOut_payload_0_2748;
    _zz_dataOut_payload_0_2765 <= _zz_dataOut_payload_0_2749;
    _zz_dataOut_payload_0_2766 <= _zz_dataOut_payload_0_2750;
    _zz_dataOut_payload_0_2767 <= _zz_dataOut_payload_0_2751;
    _zz_dataOut_payload_0_2768 <= _zz_dataOut_payload_0_2760;
    _zz_dataOut_payload_0_2769 <= _zz_dataOut_payload_0_2761;
    _zz_dataOut_payload_0_2770 <= _zz_dataOut_payload_0_2762;
    _zz_dataOut_payload_0_2771 <= _zz_dataOut_payload_0_2763;
    _zz_dataOut_payload_0_2792 <= (_zz_dataOut_payload_0_2790 ? _zz_dataOut_payload_0_2785 : _zz_dataOut_payload_0_2788);
    _zz_dataOut_payload_0_2793 <= (_zz_dataOut_payload_0_2790 ? _zz_dataOut_payload_0_2788 : _zz_dataOut_payload_0_2785);
    _zz_dataOut_payload_0_2794 <= (_zz_dataOut_payload_0_2791 ? _zz_dataOut_payload_0_2786 : _zz_dataOut_payload_0_2789);
    _zz_dataOut_payload_0_2795 <= (_zz_dataOut_payload_0_2791 ? _zz_dataOut_payload_0_2789 : _zz_dataOut_payload_0_2786);
    _zz_dataOut_payload_0_2804 <= (_zz_dataOut_payload_0_2802 ? _zz_dataOut_payload_0_2797 : _zz_dataOut_payload_0_2800);
    _zz_dataOut_payload_0_2805 <= (_zz_dataOut_payload_0_2802 ? _zz_dataOut_payload_0_2800 : _zz_dataOut_payload_0_2797);
    _zz_dataOut_payload_0_2806 <= (_zz_dataOut_payload_0_2803 ? _zz_dataOut_payload_0_2798 : _zz_dataOut_payload_0_2801);
    _zz_dataOut_payload_0_2807 <= (_zz_dataOut_payload_0_2803 ? _zz_dataOut_payload_0_2801 : _zz_dataOut_payload_0_2798);
    _zz_dataOut_payload_0_2808 <= _zz_dataOut_payload_0_2792;
    _zz_dataOut_payload_0_2809 <= _zz_dataOut_payload_0_2793;
    _zz_dataOut_payload_0_2810 <= _zz_dataOut_payload_0_2794;
    _zz_dataOut_payload_0_2811 <= _zz_dataOut_payload_0_2795;
    _zz_dataOut_payload_0_2812 <= _zz_dataOut_payload_0_2804;
    _zz_dataOut_payload_0_2813 <= _zz_dataOut_payload_0_2805;
    _zz_dataOut_payload_0_2814 <= _zz_dataOut_payload_0_2806;
    _zz_dataOut_payload_0_2815 <= _zz_dataOut_payload_0_2807;
    _zz_dataOut_payload_0_2816 <= _zz_dataOut_payload_0_1444;
    _zz_dataOut_payload_0_2817 <= _zz_dataOut_payload_0_1445;
    _zz_dataOut_payload_0_2818 <= _zz_dataOut_payload_0_1446;
    _zz_dataOut_payload_0_2819 <= _zz_dataOut_payload_0_1447;
    _zz_dataOut_payload_0_2820 <= _zz_dataOut_payload_0_1448;
    _zz_dataOut_payload_0_2821 <= _zz_dataOut_payload_0_1449;
    _zz_dataOut_payload_0_2822 <= _zz_dataOut_payload_0_1450;
    _zz_dataOut_payload_0_2823 <= _zz_dataOut_payload_0_1451;
    _zz_dataOut_payload_0_2824 <= _zz_dataOut_payload_0_1488;
    _zz_dataOut_payload_0_2825 <= _zz_dataOut_payload_0_1489;
    _zz_dataOut_payload_0_2826 <= _zz_dataOut_payload_0_1490;
    _zz_dataOut_payload_0_2827 <= _zz_dataOut_payload_0_1491;
    _zz_dataOut_payload_0_2828 <= _zz_dataOut_payload_0_1492;
    _zz_dataOut_payload_0_2829 <= _zz_dataOut_payload_0_1493;
    _zz_dataOut_payload_0_2830 <= _zz_dataOut_payload_0_1494;
    _zz_dataOut_payload_0_2831 <= _zz_dataOut_payload_0_1495;
    _zz_dataOut_payload_0_2832 <= _zz_dataOut_payload_0_1532;
    _zz_dataOut_payload_0_2833 <= _zz_dataOut_payload_0_1533;
    _zz_dataOut_payload_0_2834 <= _zz_dataOut_payload_0_1534;
    _zz_dataOut_payload_0_2835 <= _zz_dataOut_payload_0_1535;
    _zz_dataOut_payload_0_2836 <= _zz_dataOut_payload_0_1536;
    _zz_dataOut_payload_0_2837 <= _zz_dataOut_payload_0_1537;
    _zz_dataOut_payload_0_2838 <= _zz_dataOut_payload_0_1538;
    _zz_dataOut_payload_0_2839 <= _zz_dataOut_payload_0_1539;
    _zz_dataOut_payload_0_2840 <= _zz_dataOut_payload_0_1576;
    _zz_dataOut_payload_0_2841 <= _zz_dataOut_payload_0_1577;
    _zz_dataOut_payload_0_2842 <= _zz_dataOut_payload_0_1578;
    _zz_dataOut_payload_0_2843 <= _zz_dataOut_payload_0_1579;
    _zz_dataOut_payload_0_2844 <= _zz_dataOut_payload_0_1580;
    _zz_dataOut_payload_0_2845 <= _zz_dataOut_payload_0_1581;
    _zz_dataOut_payload_0_2846 <= _zz_dataOut_payload_0_1582;
    _zz_dataOut_payload_0_2847 <= _zz_dataOut_payload_0_1583;
    _zz_dataOut_payload_0_2848 <= _zz_dataOut_payload_0_1620;
    _zz_dataOut_payload_0_2849 <= _zz_dataOut_payload_0_1621;
    _zz_dataOut_payload_0_2850 <= _zz_dataOut_payload_0_1622;
    _zz_dataOut_payload_0_2851 <= _zz_dataOut_payload_0_1623;
    _zz_dataOut_payload_0_2852 <= _zz_dataOut_payload_0_1624;
    _zz_dataOut_payload_0_2853 <= _zz_dataOut_payload_0_1625;
    _zz_dataOut_payload_0_2854 <= _zz_dataOut_payload_0_1626;
    _zz_dataOut_payload_0_2855 <= _zz_dataOut_payload_0_1627;
    _zz_dataOut_payload_0_2856 <= _zz_dataOut_payload_0_1664;
    _zz_dataOut_payload_0_2857 <= _zz_dataOut_payload_0_1665;
    _zz_dataOut_payload_0_2858 <= _zz_dataOut_payload_0_1666;
    _zz_dataOut_payload_0_2859 <= _zz_dataOut_payload_0_1667;
    _zz_dataOut_payload_0_2860 <= _zz_dataOut_payload_0_1668;
    _zz_dataOut_payload_0_2861 <= _zz_dataOut_payload_0_1669;
    _zz_dataOut_payload_0_2862 <= _zz_dataOut_payload_0_1670;
    _zz_dataOut_payload_0_2863 <= _zz_dataOut_payload_0_1671;
    _zz_dataOut_payload_0_2864 <= _zz_dataOut_payload_0_1708;
    _zz_dataOut_payload_0_2865 <= _zz_dataOut_payload_0_1709;
    _zz_dataOut_payload_0_2866 <= _zz_dataOut_payload_0_1710;
    _zz_dataOut_payload_0_2867 <= _zz_dataOut_payload_0_1711;
    _zz_dataOut_payload_0_2868 <= _zz_dataOut_payload_0_1712;
    _zz_dataOut_payload_0_2869 <= _zz_dataOut_payload_0_1713;
    _zz_dataOut_payload_0_2870 <= _zz_dataOut_payload_0_1714;
    _zz_dataOut_payload_0_2871 <= _zz_dataOut_payload_0_1715;
    _zz_dataOut_payload_0_2872 <= _zz_dataOut_payload_0_1752;
    _zz_dataOut_payload_0_2873 <= _zz_dataOut_payload_0_1753;
    _zz_dataOut_payload_0_2874 <= _zz_dataOut_payload_0_1754;
    _zz_dataOut_payload_0_2875 <= _zz_dataOut_payload_0_1755;
    _zz_dataOut_payload_0_2876 <= _zz_dataOut_payload_0_1756;
    _zz_dataOut_payload_0_2877 <= _zz_dataOut_payload_0_1757;
    _zz_dataOut_payload_0_2878 <= _zz_dataOut_payload_0_1758;
    _zz_dataOut_payload_0_2879 <= _zz_dataOut_payload_0_1759;
    _zz_dataOut_payload_0_2880 <= _zz_dataOut_payload_0_1796;
    _zz_dataOut_payload_0_2881 <= _zz_dataOut_payload_0_1797;
    _zz_dataOut_payload_0_2882 <= _zz_dataOut_payload_0_1798;
    _zz_dataOut_payload_0_2883 <= _zz_dataOut_payload_0_1799;
    _zz_dataOut_payload_0_2884 <= _zz_dataOut_payload_0_1800;
    _zz_dataOut_payload_0_2885 <= _zz_dataOut_payload_0_1801;
    _zz_dataOut_payload_0_2886 <= _zz_dataOut_payload_0_1802;
    _zz_dataOut_payload_0_2887 <= _zz_dataOut_payload_0_1803;
    _zz_dataOut_payload_0_2888 <= _zz_dataOut_payload_0_1840;
    _zz_dataOut_payload_0_2889 <= _zz_dataOut_payload_0_1841;
    _zz_dataOut_payload_0_2890 <= _zz_dataOut_payload_0_1842;
    _zz_dataOut_payload_0_2891 <= _zz_dataOut_payload_0_1843;
    _zz_dataOut_payload_0_2892 <= _zz_dataOut_payload_0_1844;
    _zz_dataOut_payload_0_2893 <= _zz_dataOut_payload_0_1845;
    _zz_dataOut_payload_0_2894 <= _zz_dataOut_payload_0_1846;
    _zz_dataOut_payload_0_2895 <= _zz_dataOut_payload_0_1847;
    _zz_dataOut_payload_0_2896 <= _zz_dataOut_payload_0_1884;
    _zz_dataOut_payload_0_2897 <= _zz_dataOut_payload_0_1885;
    _zz_dataOut_payload_0_2898 <= _zz_dataOut_payload_0_1886;
    _zz_dataOut_payload_0_2899 <= _zz_dataOut_payload_0_1887;
    _zz_dataOut_payload_0_2900 <= _zz_dataOut_payload_0_1888;
    _zz_dataOut_payload_0_2901 <= _zz_dataOut_payload_0_1889;
    _zz_dataOut_payload_0_2902 <= _zz_dataOut_payload_0_1890;
    _zz_dataOut_payload_0_2903 <= _zz_dataOut_payload_0_1891;
    _zz_dataOut_payload_0_2904 <= _zz_dataOut_payload_0_1928;
    _zz_dataOut_payload_0_2905 <= _zz_dataOut_payload_0_1929;
    _zz_dataOut_payload_0_2906 <= _zz_dataOut_payload_0_1930;
    _zz_dataOut_payload_0_2907 <= _zz_dataOut_payload_0_1931;
    _zz_dataOut_payload_0_2908 <= _zz_dataOut_payload_0_1932;
    _zz_dataOut_payload_0_2909 <= _zz_dataOut_payload_0_1933;
    _zz_dataOut_payload_0_2910 <= _zz_dataOut_payload_0_1934;
    _zz_dataOut_payload_0_2911 <= _zz_dataOut_payload_0_1935;
    _zz_dataOut_payload_0_2912 <= _zz_dataOut_payload_0_1972;
    _zz_dataOut_payload_0_2913 <= _zz_dataOut_payload_0_1973;
    _zz_dataOut_payload_0_2914 <= _zz_dataOut_payload_0_1974;
    _zz_dataOut_payload_0_2915 <= _zz_dataOut_payload_0_1975;
    _zz_dataOut_payload_0_2916 <= _zz_dataOut_payload_0_1976;
    _zz_dataOut_payload_0_2917 <= _zz_dataOut_payload_0_1977;
    _zz_dataOut_payload_0_2918 <= _zz_dataOut_payload_0_1978;
    _zz_dataOut_payload_0_2919 <= _zz_dataOut_payload_0_1979;
    _zz_dataOut_payload_0_2920 <= _zz_dataOut_payload_0_2016;
    _zz_dataOut_payload_0_2921 <= _zz_dataOut_payload_0_2017;
    _zz_dataOut_payload_0_2922 <= _zz_dataOut_payload_0_2018;
    _zz_dataOut_payload_0_2923 <= _zz_dataOut_payload_0_2019;
    _zz_dataOut_payload_0_2924 <= _zz_dataOut_payload_0_2020;
    _zz_dataOut_payload_0_2925 <= _zz_dataOut_payload_0_2021;
    _zz_dataOut_payload_0_2926 <= _zz_dataOut_payload_0_2022;
    _zz_dataOut_payload_0_2927 <= _zz_dataOut_payload_0_2023;
    _zz_dataOut_payload_0_2928 <= _zz_dataOut_payload_0_2060;
    _zz_dataOut_payload_0_2929 <= _zz_dataOut_payload_0_2061;
    _zz_dataOut_payload_0_2930 <= _zz_dataOut_payload_0_2062;
    _zz_dataOut_payload_0_2931 <= _zz_dataOut_payload_0_2063;
    _zz_dataOut_payload_0_2932 <= _zz_dataOut_payload_0_2064;
    _zz_dataOut_payload_0_2933 <= _zz_dataOut_payload_0_2065;
    _zz_dataOut_payload_0_2934 <= _zz_dataOut_payload_0_2066;
    _zz_dataOut_payload_0_2935 <= _zz_dataOut_payload_0_2067;
    _zz_dataOut_payload_0_2936 <= _zz_dataOut_payload_0_2104;
    _zz_dataOut_payload_0_2937 <= _zz_dataOut_payload_0_2105;
    _zz_dataOut_payload_0_2938 <= _zz_dataOut_payload_0_2106;
    _zz_dataOut_payload_0_2939 <= _zz_dataOut_payload_0_2107;
    _zz_dataOut_payload_0_2940 <= _zz_dataOut_payload_0_2108;
    _zz_dataOut_payload_0_2941 <= _zz_dataOut_payload_0_2109;
    _zz_dataOut_payload_0_2942 <= _zz_dataOut_payload_0_2110;
    _zz_dataOut_payload_0_2943 <= _zz_dataOut_payload_0_2111;
    _zz_dataOut_payload_0_2944 <= _zz_dataOut_payload_0_2148;
    _zz_dataOut_payload_0_2945 <= _zz_dataOut_payload_0_2149;
    _zz_dataOut_payload_0_2946 <= _zz_dataOut_payload_0_2150;
    _zz_dataOut_payload_0_2947 <= _zz_dataOut_payload_0_2151;
    _zz_dataOut_payload_0_2948 <= _zz_dataOut_payload_0_2152;
    _zz_dataOut_payload_0_2949 <= _zz_dataOut_payload_0_2153;
    _zz_dataOut_payload_0_2950 <= _zz_dataOut_payload_0_2154;
    _zz_dataOut_payload_0_2951 <= _zz_dataOut_payload_0_2155;
    _zz_dataOut_payload_0_2952 <= _zz_dataOut_payload_0_2192;
    _zz_dataOut_payload_0_2953 <= _zz_dataOut_payload_0_2193;
    _zz_dataOut_payload_0_2954 <= _zz_dataOut_payload_0_2194;
    _zz_dataOut_payload_0_2955 <= _zz_dataOut_payload_0_2195;
    _zz_dataOut_payload_0_2956 <= _zz_dataOut_payload_0_2196;
    _zz_dataOut_payload_0_2957 <= _zz_dataOut_payload_0_2197;
    _zz_dataOut_payload_0_2958 <= _zz_dataOut_payload_0_2198;
    _zz_dataOut_payload_0_2959 <= _zz_dataOut_payload_0_2199;
    _zz_dataOut_payload_0_2960 <= _zz_dataOut_payload_0_2236;
    _zz_dataOut_payload_0_2961 <= _zz_dataOut_payload_0_2237;
    _zz_dataOut_payload_0_2962 <= _zz_dataOut_payload_0_2238;
    _zz_dataOut_payload_0_2963 <= _zz_dataOut_payload_0_2239;
    _zz_dataOut_payload_0_2964 <= _zz_dataOut_payload_0_2240;
    _zz_dataOut_payload_0_2965 <= _zz_dataOut_payload_0_2241;
    _zz_dataOut_payload_0_2966 <= _zz_dataOut_payload_0_2242;
    _zz_dataOut_payload_0_2967 <= _zz_dataOut_payload_0_2243;
    _zz_dataOut_payload_0_2968 <= _zz_dataOut_payload_0_2280;
    _zz_dataOut_payload_0_2969 <= _zz_dataOut_payload_0_2281;
    _zz_dataOut_payload_0_2970 <= _zz_dataOut_payload_0_2282;
    _zz_dataOut_payload_0_2971 <= _zz_dataOut_payload_0_2283;
    _zz_dataOut_payload_0_2972 <= _zz_dataOut_payload_0_2284;
    _zz_dataOut_payload_0_2973 <= _zz_dataOut_payload_0_2285;
    _zz_dataOut_payload_0_2974 <= _zz_dataOut_payload_0_2286;
    _zz_dataOut_payload_0_2975 <= _zz_dataOut_payload_0_2287;
    _zz_dataOut_payload_0_2976 <= _zz_dataOut_payload_0_2324;
    _zz_dataOut_payload_0_2977 <= _zz_dataOut_payload_0_2325;
    _zz_dataOut_payload_0_2978 <= _zz_dataOut_payload_0_2326;
    _zz_dataOut_payload_0_2979 <= _zz_dataOut_payload_0_2327;
    _zz_dataOut_payload_0_2980 <= _zz_dataOut_payload_0_2328;
    _zz_dataOut_payload_0_2981 <= _zz_dataOut_payload_0_2329;
    _zz_dataOut_payload_0_2982 <= _zz_dataOut_payload_0_2330;
    _zz_dataOut_payload_0_2983 <= _zz_dataOut_payload_0_2331;
    _zz_dataOut_payload_0_2984 <= _zz_dataOut_payload_0_2368;
    _zz_dataOut_payload_0_2985 <= _zz_dataOut_payload_0_2369;
    _zz_dataOut_payload_0_2986 <= _zz_dataOut_payload_0_2370;
    _zz_dataOut_payload_0_2987 <= _zz_dataOut_payload_0_2371;
    _zz_dataOut_payload_0_2988 <= _zz_dataOut_payload_0_2372;
    _zz_dataOut_payload_0_2989 <= _zz_dataOut_payload_0_2373;
    _zz_dataOut_payload_0_2990 <= _zz_dataOut_payload_0_2374;
    _zz_dataOut_payload_0_2991 <= _zz_dataOut_payload_0_2375;
    _zz_dataOut_payload_0_2992 <= _zz_dataOut_payload_0_2412;
    _zz_dataOut_payload_0_2993 <= _zz_dataOut_payload_0_2413;
    _zz_dataOut_payload_0_2994 <= _zz_dataOut_payload_0_2414;
    _zz_dataOut_payload_0_2995 <= _zz_dataOut_payload_0_2415;
    _zz_dataOut_payload_0_2996 <= _zz_dataOut_payload_0_2416;
    _zz_dataOut_payload_0_2997 <= _zz_dataOut_payload_0_2417;
    _zz_dataOut_payload_0_2998 <= _zz_dataOut_payload_0_2418;
    _zz_dataOut_payload_0_2999 <= _zz_dataOut_payload_0_2419;
    _zz_dataOut_payload_0_3000 <= _zz_dataOut_payload_0_2456;
    _zz_dataOut_payload_0_3001 <= _zz_dataOut_payload_0_2457;
    _zz_dataOut_payload_0_3002 <= _zz_dataOut_payload_0_2458;
    _zz_dataOut_payload_0_3003 <= _zz_dataOut_payload_0_2459;
    _zz_dataOut_payload_0_3004 <= _zz_dataOut_payload_0_2460;
    _zz_dataOut_payload_0_3005 <= _zz_dataOut_payload_0_2461;
    _zz_dataOut_payload_0_3006 <= _zz_dataOut_payload_0_2462;
    _zz_dataOut_payload_0_3007 <= _zz_dataOut_payload_0_2463;
    _zz_dataOut_payload_0_3008 <= _zz_dataOut_payload_0_2500;
    _zz_dataOut_payload_0_3009 <= _zz_dataOut_payload_0_2501;
    _zz_dataOut_payload_0_3010 <= _zz_dataOut_payload_0_2502;
    _zz_dataOut_payload_0_3011 <= _zz_dataOut_payload_0_2503;
    _zz_dataOut_payload_0_3012 <= _zz_dataOut_payload_0_2504;
    _zz_dataOut_payload_0_3013 <= _zz_dataOut_payload_0_2505;
    _zz_dataOut_payload_0_3014 <= _zz_dataOut_payload_0_2506;
    _zz_dataOut_payload_0_3015 <= _zz_dataOut_payload_0_2507;
    _zz_dataOut_payload_0_3016 <= _zz_dataOut_payload_0_2544;
    _zz_dataOut_payload_0_3017 <= _zz_dataOut_payload_0_2545;
    _zz_dataOut_payload_0_3018 <= _zz_dataOut_payload_0_2546;
    _zz_dataOut_payload_0_3019 <= _zz_dataOut_payload_0_2547;
    _zz_dataOut_payload_0_3020 <= _zz_dataOut_payload_0_2548;
    _zz_dataOut_payload_0_3021 <= _zz_dataOut_payload_0_2549;
    _zz_dataOut_payload_0_3022 <= _zz_dataOut_payload_0_2550;
    _zz_dataOut_payload_0_3023 <= _zz_dataOut_payload_0_2551;
    _zz_dataOut_payload_0_3024 <= _zz_dataOut_payload_0_2588;
    _zz_dataOut_payload_0_3025 <= _zz_dataOut_payload_0_2589;
    _zz_dataOut_payload_0_3026 <= _zz_dataOut_payload_0_2590;
    _zz_dataOut_payload_0_3027 <= _zz_dataOut_payload_0_2591;
    _zz_dataOut_payload_0_3028 <= _zz_dataOut_payload_0_2592;
    _zz_dataOut_payload_0_3029 <= _zz_dataOut_payload_0_2593;
    _zz_dataOut_payload_0_3030 <= _zz_dataOut_payload_0_2594;
    _zz_dataOut_payload_0_3031 <= _zz_dataOut_payload_0_2595;
    _zz_dataOut_payload_0_3032 <= _zz_dataOut_payload_0_2632;
    _zz_dataOut_payload_0_3033 <= _zz_dataOut_payload_0_2633;
    _zz_dataOut_payload_0_3034 <= _zz_dataOut_payload_0_2634;
    _zz_dataOut_payload_0_3035 <= _zz_dataOut_payload_0_2635;
    _zz_dataOut_payload_0_3036 <= _zz_dataOut_payload_0_2636;
    _zz_dataOut_payload_0_3037 <= _zz_dataOut_payload_0_2637;
    _zz_dataOut_payload_0_3038 <= _zz_dataOut_payload_0_2638;
    _zz_dataOut_payload_0_3039 <= _zz_dataOut_payload_0_2639;
    _zz_dataOut_payload_0_3040 <= _zz_dataOut_payload_0_2676;
    _zz_dataOut_payload_0_3041 <= _zz_dataOut_payload_0_2677;
    _zz_dataOut_payload_0_3042 <= _zz_dataOut_payload_0_2678;
    _zz_dataOut_payload_0_3043 <= _zz_dataOut_payload_0_2679;
    _zz_dataOut_payload_0_3044 <= _zz_dataOut_payload_0_2680;
    _zz_dataOut_payload_0_3045 <= _zz_dataOut_payload_0_2681;
    _zz_dataOut_payload_0_3046 <= _zz_dataOut_payload_0_2682;
    _zz_dataOut_payload_0_3047 <= _zz_dataOut_payload_0_2683;
    _zz_dataOut_payload_0_3048 <= _zz_dataOut_payload_0_2720;
    _zz_dataOut_payload_0_3049 <= _zz_dataOut_payload_0_2721;
    _zz_dataOut_payload_0_3050 <= _zz_dataOut_payload_0_2722;
    _zz_dataOut_payload_0_3051 <= _zz_dataOut_payload_0_2723;
    _zz_dataOut_payload_0_3052 <= _zz_dataOut_payload_0_2724;
    _zz_dataOut_payload_0_3053 <= _zz_dataOut_payload_0_2725;
    _zz_dataOut_payload_0_3054 <= _zz_dataOut_payload_0_2726;
    _zz_dataOut_payload_0_3055 <= _zz_dataOut_payload_0_2727;
    _zz_dataOut_payload_0_3056 <= _zz_dataOut_payload_0_2764;
    _zz_dataOut_payload_0_3057 <= _zz_dataOut_payload_0_2765;
    _zz_dataOut_payload_0_3058 <= _zz_dataOut_payload_0_2766;
    _zz_dataOut_payload_0_3059 <= _zz_dataOut_payload_0_2767;
    _zz_dataOut_payload_0_3060 <= _zz_dataOut_payload_0_2768;
    _zz_dataOut_payload_0_3061 <= _zz_dataOut_payload_0_2769;
    _zz_dataOut_payload_0_3062 <= _zz_dataOut_payload_0_2770;
    _zz_dataOut_payload_0_3063 <= _zz_dataOut_payload_0_2771;
    _zz_dataOut_payload_0_3064 <= _zz_dataOut_payload_0_2808;
    _zz_dataOut_payload_0_3065 <= _zz_dataOut_payload_0_2809;
    _zz_dataOut_payload_0_3066 <= _zz_dataOut_payload_0_2810;
    _zz_dataOut_payload_0_3067 <= _zz_dataOut_payload_0_2811;
    _zz_dataOut_payload_0_3068 <= _zz_dataOut_payload_0_2812;
    _zz_dataOut_payload_0_3069 <= _zz_dataOut_payload_0_2813;
    _zz_dataOut_payload_0_3070 <= _zz_dataOut_payload_0_2814;
    _zz_dataOut_payload_0_3071 <= _zz_dataOut_payload_0_2815;
    _zz_dataOut_payload_0_3116 <= (_zz_dataOut_payload_0_3114 ? _zz_dataOut_payload_0_3109 : _zz_dataOut_payload_0_3112);
    _zz_dataOut_payload_0_3117 <= (_zz_dataOut_payload_0_3114 ? _zz_dataOut_payload_0_3112 : _zz_dataOut_payload_0_3109);
    _zz_dataOut_payload_0_3118 <= (_zz_dataOut_payload_0_3115 ? _zz_dataOut_payload_0_3110 : _zz_dataOut_payload_0_3113);
    _zz_dataOut_payload_0_3119 <= (_zz_dataOut_payload_0_3115 ? _zz_dataOut_payload_0_3113 : _zz_dataOut_payload_0_3110);
    _zz_dataOut_payload_0_3128 <= (_zz_dataOut_payload_0_3126 ? _zz_dataOut_payload_0_3121 : _zz_dataOut_payload_0_3124);
    _zz_dataOut_payload_0_3129 <= (_zz_dataOut_payload_0_3126 ? _zz_dataOut_payload_0_3124 : _zz_dataOut_payload_0_3121);
    _zz_dataOut_payload_0_3130 <= (_zz_dataOut_payload_0_3127 ? _zz_dataOut_payload_0_3122 : _zz_dataOut_payload_0_3125);
    _zz_dataOut_payload_0_3131 <= (_zz_dataOut_payload_0_3127 ? _zz_dataOut_payload_0_3125 : _zz_dataOut_payload_0_3122);
    _zz_dataOut_payload_0_3132 <= _zz_dataOut_payload_0_3116;
    _zz_dataOut_payload_0_3133 <= _zz_dataOut_payload_0_3117;
    _zz_dataOut_payload_0_3134 <= _zz_dataOut_payload_0_3118;
    _zz_dataOut_payload_0_3135 <= _zz_dataOut_payload_0_3119;
    _zz_dataOut_payload_0_3136 <= _zz_dataOut_payload_0_3128;
    _zz_dataOut_payload_0_3137 <= _zz_dataOut_payload_0_3129;
    _zz_dataOut_payload_0_3138 <= _zz_dataOut_payload_0_3130;
    _zz_dataOut_payload_0_3139 <= _zz_dataOut_payload_0_3131;
    _zz_dataOut_payload_0_3160 <= (_zz_dataOut_payload_0_3158 ? _zz_dataOut_payload_0_3153 : _zz_dataOut_payload_0_3156);
    _zz_dataOut_payload_0_3161 <= (_zz_dataOut_payload_0_3158 ? _zz_dataOut_payload_0_3156 : _zz_dataOut_payload_0_3153);
    _zz_dataOut_payload_0_3162 <= (_zz_dataOut_payload_0_3159 ? _zz_dataOut_payload_0_3154 : _zz_dataOut_payload_0_3157);
    _zz_dataOut_payload_0_3163 <= (_zz_dataOut_payload_0_3159 ? _zz_dataOut_payload_0_3157 : _zz_dataOut_payload_0_3154);
    _zz_dataOut_payload_0_3172 <= (_zz_dataOut_payload_0_3170 ? _zz_dataOut_payload_0_3165 : _zz_dataOut_payload_0_3168);
    _zz_dataOut_payload_0_3173 <= (_zz_dataOut_payload_0_3170 ? _zz_dataOut_payload_0_3168 : _zz_dataOut_payload_0_3165);
    _zz_dataOut_payload_0_3174 <= (_zz_dataOut_payload_0_3171 ? _zz_dataOut_payload_0_3166 : _zz_dataOut_payload_0_3169);
    _zz_dataOut_payload_0_3175 <= (_zz_dataOut_payload_0_3171 ? _zz_dataOut_payload_0_3169 : _zz_dataOut_payload_0_3166);
    _zz_dataOut_payload_0_3176 <= _zz_dataOut_payload_0_3160;
    _zz_dataOut_payload_0_3177 <= _zz_dataOut_payload_0_3161;
    _zz_dataOut_payload_0_3178 <= _zz_dataOut_payload_0_3162;
    _zz_dataOut_payload_0_3179 <= _zz_dataOut_payload_0_3163;
    _zz_dataOut_payload_0_3180 <= _zz_dataOut_payload_0_3172;
    _zz_dataOut_payload_0_3181 <= _zz_dataOut_payload_0_3173;
    _zz_dataOut_payload_0_3182 <= _zz_dataOut_payload_0_3174;
    _zz_dataOut_payload_0_3183 <= _zz_dataOut_payload_0_3175;
    _zz_dataOut_payload_0_3184 <= _zz_dataOut_payload_0_3132;
    _zz_dataOut_payload_0_3185 <= _zz_dataOut_payload_0_3133;
    _zz_dataOut_payload_0_3186 <= _zz_dataOut_payload_0_3134;
    _zz_dataOut_payload_0_3187 <= _zz_dataOut_payload_0_3135;
    _zz_dataOut_payload_0_3188 <= _zz_dataOut_payload_0_3136;
    _zz_dataOut_payload_0_3189 <= _zz_dataOut_payload_0_3137;
    _zz_dataOut_payload_0_3190 <= _zz_dataOut_payload_0_3138;
    _zz_dataOut_payload_0_3191 <= _zz_dataOut_payload_0_3139;
    _zz_dataOut_payload_0_3192 <= _zz_dataOut_payload_0_3176;
    _zz_dataOut_payload_0_3193 <= _zz_dataOut_payload_0_3177;
    _zz_dataOut_payload_0_3194 <= _zz_dataOut_payload_0_3178;
    _zz_dataOut_payload_0_3195 <= _zz_dataOut_payload_0_3179;
    _zz_dataOut_payload_0_3196 <= _zz_dataOut_payload_0_3180;
    _zz_dataOut_payload_0_3197 <= _zz_dataOut_payload_0_3181;
    _zz_dataOut_payload_0_3198 <= _zz_dataOut_payload_0_3182;
    _zz_dataOut_payload_0_3199 <= _zz_dataOut_payload_0_3183;
    _zz_dataOut_payload_0_3244 <= (_zz_dataOut_payload_0_3242 ? _zz_dataOut_payload_0_3237 : _zz_dataOut_payload_0_3240);
    _zz_dataOut_payload_0_3245 <= (_zz_dataOut_payload_0_3242 ? _zz_dataOut_payload_0_3240 : _zz_dataOut_payload_0_3237);
    _zz_dataOut_payload_0_3246 <= (_zz_dataOut_payload_0_3243 ? _zz_dataOut_payload_0_3238 : _zz_dataOut_payload_0_3241);
    _zz_dataOut_payload_0_3247 <= (_zz_dataOut_payload_0_3243 ? _zz_dataOut_payload_0_3241 : _zz_dataOut_payload_0_3238);
    _zz_dataOut_payload_0_3256 <= (_zz_dataOut_payload_0_3254 ? _zz_dataOut_payload_0_3249 : _zz_dataOut_payload_0_3252);
    _zz_dataOut_payload_0_3257 <= (_zz_dataOut_payload_0_3254 ? _zz_dataOut_payload_0_3252 : _zz_dataOut_payload_0_3249);
    _zz_dataOut_payload_0_3258 <= (_zz_dataOut_payload_0_3255 ? _zz_dataOut_payload_0_3250 : _zz_dataOut_payload_0_3253);
    _zz_dataOut_payload_0_3259 <= (_zz_dataOut_payload_0_3255 ? _zz_dataOut_payload_0_3253 : _zz_dataOut_payload_0_3250);
    _zz_dataOut_payload_0_3260 <= _zz_dataOut_payload_0_3244;
    _zz_dataOut_payload_0_3261 <= _zz_dataOut_payload_0_3245;
    _zz_dataOut_payload_0_3262 <= _zz_dataOut_payload_0_3246;
    _zz_dataOut_payload_0_3263 <= _zz_dataOut_payload_0_3247;
    _zz_dataOut_payload_0_3264 <= _zz_dataOut_payload_0_3256;
    _zz_dataOut_payload_0_3265 <= _zz_dataOut_payload_0_3257;
    _zz_dataOut_payload_0_3266 <= _zz_dataOut_payload_0_3258;
    _zz_dataOut_payload_0_3267 <= _zz_dataOut_payload_0_3259;
    _zz_dataOut_payload_0_3288 <= (_zz_dataOut_payload_0_3286 ? _zz_dataOut_payload_0_3281 : _zz_dataOut_payload_0_3284);
    _zz_dataOut_payload_0_3289 <= (_zz_dataOut_payload_0_3286 ? _zz_dataOut_payload_0_3284 : _zz_dataOut_payload_0_3281);
    _zz_dataOut_payload_0_3290 <= (_zz_dataOut_payload_0_3287 ? _zz_dataOut_payload_0_3282 : _zz_dataOut_payload_0_3285);
    _zz_dataOut_payload_0_3291 <= (_zz_dataOut_payload_0_3287 ? _zz_dataOut_payload_0_3285 : _zz_dataOut_payload_0_3282);
    _zz_dataOut_payload_0_3300 <= (_zz_dataOut_payload_0_3298 ? _zz_dataOut_payload_0_3293 : _zz_dataOut_payload_0_3296);
    _zz_dataOut_payload_0_3301 <= (_zz_dataOut_payload_0_3298 ? _zz_dataOut_payload_0_3296 : _zz_dataOut_payload_0_3293);
    _zz_dataOut_payload_0_3302 <= (_zz_dataOut_payload_0_3299 ? _zz_dataOut_payload_0_3294 : _zz_dataOut_payload_0_3297);
    _zz_dataOut_payload_0_3303 <= (_zz_dataOut_payload_0_3299 ? _zz_dataOut_payload_0_3297 : _zz_dataOut_payload_0_3294);
    _zz_dataOut_payload_0_3304 <= _zz_dataOut_payload_0_3288;
    _zz_dataOut_payload_0_3305 <= _zz_dataOut_payload_0_3289;
    _zz_dataOut_payload_0_3306 <= _zz_dataOut_payload_0_3290;
    _zz_dataOut_payload_0_3307 <= _zz_dataOut_payload_0_3291;
    _zz_dataOut_payload_0_3308 <= _zz_dataOut_payload_0_3300;
    _zz_dataOut_payload_0_3309 <= _zz_dataOut_payload_0_3301;
    _zz_dataOut_payload_0_3310 <= _zz_dataOut_payload_0_3302;
    _zz_dataOut_payload_0_3311 <= _zz_dataOut_payload_0_3303;
    _zz_dataOut_payload_0_3312 <= _zz_dataOut_payload_0_3260;
    _zz_dataOut_payload_0_3313 <= _zz_dataOut_payload_0_3261;
    _zz_dataOut_payload_0_3314 <= _zz_dataOut_payload_0_3262;
    _zz_dataOut_payload_0_3315 <= _zz_dataOut_payload_0_3263;
    _zz_dataOut_payload_0_3316 <= _zz_dataOut_payload_0_3264;
    _zz_dataOut_payload_0_3317 <= _zz_dataOut_payload_0_3265;
    _zz_dataOut_payload_0_3318 <= _zz_dataOut_payload_0_3266;
    _zz_dataOut_payload_0_3319 <= _zz_dataOut_payload_0_3267;
    _zz_dataOut_payload_0_3320 <= _zz_dataOut_payload_0_3304;
    _zz_dataOut_payload_0_3321 <= _zz_dataOut_payload_0_3305;
    _zz_dataOut_payload_0_3322 <= _zz_dataOut_payload_0_3306;
    _zz_dataOut_payload_0_3323 <= _zz_dataOut_payload_0_3307;
    _zz_dataOut_payload_0_3324 <= _zz_dataOut_payload_0_3308;
    _zz_dataOut_payload_0_3325 <= _zz_dataOut_payload_0_3309;
    _zz_dataOut_payload_0_3326 <= _zz_dataOut_payload_0_3310;
    _zz_dataOut_payload_0_3327 <= _zz_dataOut_payload_0_3311;
    _zz_dataOut_payload_0_3372 <= (_zz_dataOut_payload_0_3370 ? _zz_dataOut_payload_0_3365 : _zz_dataOut_payload_0_3368);
    _zz_dataOut_payload_0_3373 <= (_zz_dataOut_payload_0_3370 ? _zz_dataOut_payload_0_3368 : _zz_dataOut_payload_0_3365);
    _zz_dataOut_payload_0_3374 <= (_zz_dataOut_payload_0_3371 ? _zz_dataOut_payload_0_3366 : _zz_dataOut_payload_0_3369);
    _zz_dataOut_payload_0_3375 <= (_zz_dataOut_payload_0_3371 ? _zz_dataOut_payload_0_3369 : _zz_dataOut_payload_0_3366);
    _zz_dataOut_payload_0_3384 <= (_zz_dataOut_payload_0_3382 ? _zz_dataOut_payload_0_3377 : _zz_dataOut_payload_0_3380);
    _zz_dataOut_payload_0_3385 <= (_zz_dataOut_payload_0_3382 ? _zz_dataOut_payload_0_3380 : _zz_dataOut_payload_0_3377);
    _zz_dataOut_payload_0_3386 <= (_zz_dataOut_payload_0_3383 ? _zz_dataOut_payload_0_3378 : _zz_dataOut_payload_0_3381);
    _zz_dataOut_payload_0_3387 <= (_zz_dataOut_payload_0_3383 ? _zz_dataOut_payload_0_3381 : _zz_dataOut_payload_0_3378);
    _zz_dataOut_payload_0_3388 <= _zz_dataOut_payload_0_3372;
    _zz_dataOut_payload_0_3389 <= _zz_dataOut_payload_0_3373;
    _zz_dataOut_payload_0_3390 <= _zz_dataOut_payload_0_3374;
    _zz_dataOut_payload_0_3391 <= _zz_dataOut_payload_0_3375;
    _zz_dataOut_payload_0_3392 <= _zz_dataOut_payload_0_3384;
    _zz_dataOut_payload_0_3393 <= _zz_dataOut_payload_0_3385;
    _zz_dataOut_payload_0_3394 <= _zz_dataOut_payload_0_3386;
    _zz_dataOut_payload_0_3395 <= _zz_dataOut_payload_0_3387;
    _zz_dataOut_payload_0_3416 <= (_zz_dataOut_payload_0_3414 ? _zz_dataOut_payload_0_3409 : _zz_dataOut_payload_0_3412);
    _zz_dataOut_payload_0_3417 <= (_zz_dataOut_payload_0_3414 ? _zz_dataOut_payload_0_3412 : _zz_dataOut_payload_0_3409);
    _zz_dataOut_payload_0_3418 <= (_zz_dataOut_payload_0_3415 ? _zz_dataOut_payload_0_3410 : _zz_dataOut_payload_0_3413);
    _zz_dataOut_payload_0_3419 <= (_zz_dataOut_payload_0_3415 ? _zz_dataOut_payload_0_3413 : _zz_dataOut_payload_0_3410);
    _zz_dataOut_payload_0_3428 <= (_zz_dataOut_payload_0_3426 ? _zz_dataOut_payload_0_3421 : _zz_dataOut_payload_0_3424);
    _zz_dataOut_payload_0_3429 <= (_zz_dataOut_payload_0_3426 ? _zz_dataOut_payload_0_3424 : _zz_dataOut_payload_0_3421);
    _zz_dataOut_payload_0_3430 <= (_zz_dataOut_payload_0_3427 ? _zz_dataOut_payload_0_3422 : _zz_dataOut_payload_0_3425);
    _zz_dataOut_payload_0_3431 <= (_zz_dataOut_payload_0_3427 ? _zz_dataOut_payload_0_3425 : _zz_dataOut_payload_0_3422);
    _zz_dataOut_payload_0_3432 <= _zz_dataOut_payload_0_3416;
    _zz_dataOut_payload_0_3433 <= _zz_dataOut_payload_0_3417;
    _zz_dataOut_payload_0_3434 <= _zz_dataOut_payload_0_3418;
    _zz_dataOut_payload_0_3435 <= _zz_dataOut_payload_0_3419;
    _zz_dataOut_payload_0_3436 <= _zz_dataOut_payload_0_3428;
    _zz_dataOut_payload_0_3437 <= _zz_dataOut_payload_0_3429;
    _zz_dataOut_payload_0_3438 <= _zz_dataOut_payload_0_3430;
    _zz_dataOut_payload_0_3439 <= _zz_dataOut_payload_0_3431;
    _zz_dataOut_payload_0_3440 <= _zz_dataOut_payload_0_3388;
    _zz_dataOut_payload_0_3441 <= _zz_dataOut_payload_0_3389;
    _zz_dataOut_payload_0_3442 <= _zz_dataOut_payload_0_3390;
    _zz_dataOut_payload_0_3443 <= _zz_dataOut_payload_0_3391;
    _zz_dataOut_payload_0_3444 <= _zz_dataOut_payload_0_3392;
    _zz_dataOut_payload_0_3445 <= _zz_dataOut_payload_0_3393;
    _zz_dataOut_payload_0_3446 <= _zz_dataOut_payload_0_3394;
    _zz_dataOut_payload_0_3447 <= _zz_dataOut_payload_0_3395;
    _zz_dataOut_payload_0_3448 <= _zz_dataOut_payload_0_3432;
    _zz_dataOut_payload_0_3449 <= _zz_dataOut_payload_0_3433;
    _zz_dataOut_payload_0_3450 <= _zz_dataOut_payload_0_3434;
    _zz_dataOut_payload_0_3451 <= _zz_dataOut_payload_0_3435;
    _zz_dataOut_payload_0_3452 <= _zz_dataOut_payload_0_3436;
    _zz_dataOut_payload_0_3453 <= _zz_dataOut_payload_0_3437;
    _zz_dataOut_payload_0_3454 <= _zz_dataOut_payload_0_3438;
    _zz_dataOut_payload_0_3455 <= _zz_dataOut_payload_0_3439;
    _zz_dataOut_payload_0_3500 <= (_zz_dataOut_payload_0_3498 ? _zz_dataOut_payload_0_3493 : _zz_dataOut_payload_0_3496);
    _zz_dataOut_payload_0_3501 <= (_zz_dataOut_payload_0_3498 ? _zz_dataOut_payload_0_3496 : _zz_dataOut_payload_0_3493);
    _zz_dataOut_payload_0_3502 <= (_zz_dataOut_payload_0_3499 ? _zz_dataOut_payload_0_3494 : _zz_dataOut_payload_0_3497);
    _zz_dataOut_payload_0_3503 <= (_zz_dataOut_payload_0_3499 ? _zz_dataOut_payload_0_3497 : _zz_dataOut_payload_0_3494);
    _zz_dataOut_payload_0_3512 <= (_zz_dataOut_payload_0_3510 ? _zz_dataOut_payload_0_3505 : _zz_dataOut_payload_0_3508);
    _zz_dataOut_payload_0_3513 <= (_zz_dataOut_payload_0_3510 ? _zz_dataOut_payload_0_3508 : _zz_dataOut_payload_0_3505);
    _zz_dataOut_payload_0_3514 <= (_zz_dataOut_payload_0_3511 ? _zz_dataOut_payload_0_3506 : _zz_dataOut_payload_0_3509);
    _zz_dataOut_payload_0_3515 <= (_zz_dataOut_payload_0_3511 ? _zz_dataOut_payload_0_3509 : _zz_dataOut_payload_0_3506);
    _zz_dataOut_payload_0_3516 <= _zz_dataOut_payload_0_3500;
    _zz_dataOut_payload_0_3517 <= _zz_dataOut_payload_0_3501;
    _zz_dataOut_payload_0_3518 <= _zz_dataOut_payload_0_3502;
    _zz_dataOut_payload_0_3519 <= _zz_dataOut_payload_0_3503;
    _zz_dataOut_payload_0_3520 <= _zz_dataOut_payload_0_3512;
    _zz_dataOut_payload_0_3521 <= _zz_dataOut_payload_0_3513;
    _zz_dataOut_payload_0_3522 <= _zz_dataOut_payload_0_3514;
    _zz_dataOut_payload_0_3523 <= _zz_dataOut_payload_0_3515;
    _zz_dataOut_payload_0_3544 <= (_zz_dataOut_payload_0_3542 ? _zz_dataOut_payload_0_3537 : _zz_dataOut_payload_0_3540);
    _zz_dataOut_payload_0_3545 <= (_zz_dataOut_payload_0_3542 ? _zz_dataOut_payload_0_3540 : _zz_dataOut_payload_0_3537);
    _zz_dataOut_payload_0_3546 <= (_zz_dataOut_payload_0_3543 ? _zz_dataOut_payload_0_3538 : _zz_dataOut_payload_0_3541);
    _zz_dataOut_payload_0_3547 <= (_zz_dataOut_payload_0_3543 ? _zz_dataOut_payload_0_3541 : _zz_dataOut_payload_0_3538);
    _zz_dataOut_payload_0_3556 <= (_zz_dataOut_payload_0_3554 ? _zz_dataOut_payload_0_3549 : _zz_dataOut_payload_0_3552);
    _zz_dataOut_payload_0_3557 <= (_zz_dataOut_payload_0_3554 ? _zz_dataOut_payload_0_3552 : _zz_dataOut_payload_0_3549);
    _zz_dataOut_payload_0_3558 <= (_zz_dataOut_payload_0_3555 ? _zz_dataOut_payload_0_3550 : _zz_dataOut_payload_0_3553);
    _zz_dataOut_payload_0_3559 <= (_zz_dataOut_payload_0_3555 ? _zz_dataOut_payload_0_3553 : _zz_dataOut_payload_0_3550);
    _zz_dataOut_payload_0_3560 <= _zz_dataOut_payload_0_3544;
    _zz_dataOut_payload_0_3561 <= _zz_dataOut_payload_0_3545;
    _zz_dataOut_payload_0_3562 <= _zz_dataOut_payload_0_3546;
    _zz_dataOut_payload_0_3563 <= _zz_dataOut_payload_0_3547;
    _zz_dataOut_payload_0_3564 <= _zz_dataOut_payload_0_3556;
    _zz_dataOut_payload_0_3565 <= _zz_dataOut_payload_0_3557;
    _zz_dataOut_payload_0_3566 <= _zz_dataOut_payload_0_3558;
    _zz_dataOut_payload_0_3567 <= _zz_dataOut_payload_0_3559;
    _zz_dataOut_payload_0_3568 <= _zz_dataOut_payload_0_3516;
    _zz_dataOut_payload_0_3569 <= _zz_dataOut_payload_0_3517;
    _zz_dataOut_payload_0_3570 <= _zz_dataOut_payload_0_3518;
    _zz_dataOut_payload_0_3571 <= _zz_dataOut_payload_0_3519;
    _zz_dataOut_payload_0_3572 <= _zz_dataOut_payload_0_3520;
    _zz_dataOut_payload_0_3573 <= _zz_dataOut_payload_0_3521;
    _zz_dataOut_payload_0_3574 <= _zz_dataOut_payload_0_3522;
    _zz_dataOut_payload_0_3575 <= _zz_dataOut_payload_0_3523;
    _zz_dataOut_payload_0_3576 <= _zz_dataOut_payload_0_3560;
    _zz_dataOut_payload_0_3577 <= _zz_dataOut_payload_0_3561;
    _zz_dataOut_payload_0_3578 <= _zz_dataOut_payload_0_3562;
    _zz_dataOut_payload_0_3579 <= _zz_dataOut_payload_0_3563;
    _zz_dataOut_payload_0_3580 <= _zz_dataOut_payload_0_3564;
    _zz_dataOut_payload_0_3581 <= _zz_dataOut_payload_0_3565;
    _zz_dataOut_payload_0_3582 <= _zz_dataOut_payload_0_3566;
    _zz_dataOut_payload_0_3583 <= _zz_dataOut_payload_0_3567;
    _zz_dataOut_payload_0_3628 <= (_zz_dataOut_payload_0_3626 ? _zz_dataOut_payload_0_3621 : _zz_dataOut_payload_0_3624);
    _zz_dataOut_payload_0_3629 <= (_zz_dataOut_payload_0_3626 ? _zz_dataOut_payload_0_3624 : _zz_dataOut_payload_0_3621);
    _zz_dataOut_payload_0_3630 <= (_zz_dataOut_payload_0_3627 ? _zz_dataOut_payload_0_3622 : _zz_dataOut_payload_0_3625);
    _zz_dataOut_payload_0_3631 <= (_zz_dataOut_payload_0_3627 ? _zz_dataOut_payload_0_3625 : _zz_dataOut_payload_0_3622);
    _zz_dataOut_payload_0_3640 <= (_zz_dataOut_payload_0_3638 ? _zz_dataOut_payload_0_3633 : _zz_dataOut_payload_0_3636);
    _zz_dataOut_payload_0_3641 <= (_zz_dataOut_payload_0_3638 ? _zz_dataOut_payload_0_3636 : _zz_dataOut_payload_0_3633);
    _zz_dataOut_payload_0_3642 <= (_zz_dataOut_payload_0_3639 ? _zz_dataOut_payload_0_3634 : _zz_dataOut_payload_0_3637);
    _zz_dataOut_payload_0_3643 <= (_zz_dataOut_payload_0_3639 ? _zz_dataOut_payload_0_3637 : _zz_dataOut_payload_0_3634);
    _zz_dataOut_payload_0_3644 <= _zz_dataOut_payload_0_3628;
    _zz_dataOut_payload_0_3645 <= _zz_dataOut_payload_0_3629;
    _zz_dataOut_payload_0_3646 <= _zz_dataOut_payload_0_3630;
    _zz_dataOut_payload_0_3647 <= _zz_dataOut_payload_0_3631;
    _zz_dataOut_payload_0_3648 <= _zz_dataOut_payload_0_3640;
    _zz_dataOut_payload_0_3649 <= _zz_dataOut_payload_0_3641;
    _zz_dataOut_payload_0_3650 <= _zz_dataOut_payload_0_3642;
    _zz_dataOut_payload_0_3651 <= _zz_dataOut_payload_0_3643;
    _zz_dataOut_payload_0_3672 <= (_zz_dataOut_payload_0_3670 ? _zz_dataOut_payload_0_3665 : _zz_dataOut_payload_0_3668);
    _zz_dataOut_payload_0_3673 <= (_zz_dataOut_payload_0_3670 ? _zz_dataOut_payload_0_3668 : _zz_dataOut_payload_0_3665);
    _zz_dataOut_payload_0_3674 <= (_zz_dataOut_payload_0_3671 ? _zz_dataOut_payload_0_3666 : _zz_dataOut_payload_0_3669);
    _zz_dataOut_payload_0_3675 <= (_zz_dataOut_payload_0_3671 ? _zz_dataOut_payload_0_3669 : _zz_dataOut_payload_0_3666);
    _zz_dataOut_payload_0_3684 <= (_zz_dataOut_payload_0_3682 ? _zz_dataOut_payload_0_3677 : _zz_dataOut_payload_0_3680);
    _zz_dataOut_payload_0_3685 <= (_zz_dataOut_payload_0_3682 ? _zz_dataOut_payload_0_3680 : _zz_dataOut_payload_0_3677);
    _zz_dataOut_payload_0_3686 <= (_zz_dataOut_payload_0_3683 ? _zz_dataOut_payload_0_3678 : _zz_dataOut_payload_0_3681);
    _zz_dataOut_payload_0_3687 <= (_zz_dataOut_payload_0_3683 ? _zz_dataOut_payload_0_3681 : _zz_dataOut_payload_0_3678);
    _zz_dataOut_payload_0_3688 <= _zz_dataOut_payload_0_3672;
    _zz_dataOut_payload_0_3689 <= _zz_dataOut_payload_0_3673;
    _zz_dataOut_payload_0_3690 <= _zz_dataOut_payload_0_3674;
    _zz_dataOut_payload_0_3691 <= _zz_dataOut_payload_0_3675;
    _zz_dataOut_payload_0_3692 <= _zz_dataOut_payload_0_3684;
    _zz_dataOut_payload_0_3693 <= _zz_dataOut_payload_0_3685;
    _zz_dataOut_payload_0_3694 <= _zz_dataOut_payload_0_3686;
    _zz_dataOut_payload_0_3695 <= _zz_dataOut_payload_0_3687;
    _zz_dataOut_payload_0_3696 <= _zz_dataOut_payload_0_3644;
    _zz_dataOut_payload_0_3697 <= _zz_dataOut_payload_0_3645;
    _zz_dataOut_payload_0_3698 <= _zz_dataOut_payload_0_3646;
    _zz_dataOut_payload_0_3699 <= _zz_dataOut_payload_0_3647;
    _zz_dataOut_payload_0_3700 <= _zz_dataOut_payload_0_3648;
    _zz_dataOut_payload_0_3701 <= _zz_dataOut_payload_0_3649;
    _zz_dataOut_payload_0_3702 <= _zz_dataOut_payload_0_3650;
    _zz_dataOut_payload_0_3703 <= _zz_dataOut_payload_0_3651;
    _zz_dataOut_payload_0_3704 <= _zz_dataOut_payload_0_3688;
    _zz_dataOut_payload_0_3705 <= _zz_dataOut_payload_0_3689;
    _zz_dataOut_payload_0_3706 <= _zz_dataOut_payload_0_3690;
    _zz_dataOut_payload_0_3707 <= _zz_dataOut_payload_0_3691;
    _zz_dataOut_payload_0_3708 <= _zz_dataOut_payload_0_3692;
    _zz_dataOut_payload_0_3709 <= _zz_dataOut_payload_0_3693;
    _zz_dataOut_payload_0_3710 <= _zz_dataOut_payload_0_3694;
    _zz_dataOut_payload_0_3711 <= _zz_dataOut_payload_0_3695;
    _zz_dataOut_payload_0_3756 <= (_zz_dataOut_payload_0_3754 ? _zz_dataOut_payload_0_3749 : _zz_dataOut_payload_0_3752);
    _zz_dataOut_payload_0_3757 <= (_zz_dataOut_payload_0_3754 ? _zz_dataOut_payload_0_3752 : _zz_dataOut_payload_0_3749);
    _zz_dataOut_payload_0_3758 <= (_zz_dataOut_payload_0_3755 ? _zz_dataOut_payload_0_3750 : _zz_dataOut_payload_0_3753);
    _zz_dataOut_payload_0_3759 <= (_zz_dataOut_payload_0_3755 ? _zz_dataOut_payload_0_3753 : _zz_dataOut_payload_0_3750);
    _zz_dataOut_payload_0_3768 <= (_zz_dataOut_payload_0_3766 ? _zz_dataOut_payload_0_3761 : _zz_dataOut_payload_0_3764);
    _zz_dataOut_payload_0_3769 <= (_zz_dataOut_payload_0_3766 ? _zz_dataOut_payload_0_3764 : _zz_dataOut_payload_0_3761);
    _zz_dataOut_payload_0_3770 <= (_zz_dataOut_payload_0_3767 ? _zz_dataOut_payload_0_3762 : _zz_dataOut_payload_0_3765);
    _zz_dataOut_payload_0_3771 <= (_zz_dataOut_payload_0_3767 ? _zz_dataOut_payload_0_3765 : _zz_dataOut_payload_0_3762);
    _zz_dataOut_payload_0_3772 <= _zz_dataOut_payload_0_3756;
    _zz_dataOut_payload_0_3773 <= _zz_dataOut_payload_0_3757;
    _zz_dataOut_payload_0_3774 <= _zz_dataOut_payload_0_3758;
    _zz_dataOut_payload_0_3775 <= _zz_dataOut_payload_0_3759;
    _zz_dataOut_payload_0_3776 <= _zz_dataOut_payload_0_3768;
    _zz_dataOut_payload_0_3777 <= _zz_dataOut_payload_0_3769;
    _zz_dataOut_payload_0_3778 <= _zz_dataOut_payload_0_3770;
    _zz_dataOut_payload_0_3779 <= _zz_dataOut_payload_0_3771;
    _zz_dataOut_payload_0_3800 <= (_zz_dataOut_payload_0_3798 ? _zz_dataOut_payload_0_3793 : _zz_dataOut_payload_0_3796);
    _zz_dataOut_payload_0_3801 <= (_zz_dataOut_payload_0_3798 ? _zz_dataOut_payload_0_3796 : _zz_dataOut_payload_0_3793);
    _zz_dataOut_payload_0_3802 <= (_zz_dataOut_payload_0_3799 ? _zz_dataOut_payload_0_3794 : _zz_dataOut_payload_0_3797);
    _zz_dataOut_payload_0_3803 <= (_zz_dataOut_payload_0_3799 ? _zz_dataOut_payload_0_3797 : _zz_dataOut_payload_0_3794);
    _zz_dataOut_payload_0_3812 <= (_zz_dataOut_payload_0_3810 ? _zz_dataOut_payload_0_3805 : _zz_dataOut_payload_0_3808);
    _zz_dataOut_payload_0_3813 <= (_zz_dataOut_payload_0_3810 ? _zz_dataOut_payload_0_3808 : _zz_dataOut_payload_0_3805);
    _zz_dataOut_payload_0_3814 <= (_zz_dataOut_payload_0_3811 ? _zz_dataOut_payload_0_3806 : _zz_dataOut_payload_0_3809);
    _zz_dataOut_payload_0_3815 <= (_zz_dataOut_payload_0_3811 ? _zz_dataOut_payload_0_3809 : _zz_dataOut_payload_0_3806);
    _zz_dataOut_payload_0_3816 <= _zz_dataOut_payload_0_3800;
    _zz_dataOut_payload_0_3817 <= _zz_dataOut_payload_0_3801;
    _zz_dataOut_payload_0_3818 <= _zz_dataOut_payload_0_3802;
    _zz_dataOut_payload_0_3819 <= _zz_dataOut_payload_0_3803;
    _zz_dataOut_payload_0_3820 <= _zz_dataOut_payload_0_3812;
    _zz_dataOut_payload_0_3821 <= _zz_dataOut_payload_0_3813;
    _zz_dataOut_payload_0_3822 <= _zz_dataOut_payload_0_3814;
    _zz_dataOut_payload_0_3823 <= _zz_dataOut_payload_0_3815;
    _zz_dataOut_payload_0_3824 <= _zz_dataOut_payload_0_3772;
    _zz_dataOut_payload_0_3825 <= _zz_dataOut_payload_0_3773;
    _zz_dataOut_payload_0_3826 <= _zz_dataOut_payload_0_3774;
    _zz_dataOut_payload_0_3827 <= _zz_dataOut_payload_0_3775;
    _zz_dataOut_payload_0_3828 <= _zz_dataOut_payload_0_3776;
    _zz_dataOut_payload_0_3829 <= _zz_dataOut_payload_0_3777;
    _zz_dataOut_payload_0_3830 <= _zz_dataOut_payload_0_3778;
    _zz_dataOut_payload_0_3831 <= _zz_dataOut_payload_0_3779;
    _zz_dataOut_payload_0_3832 <= _zz_dataOut_payload_0_3816;
    _zz_dataOut_payload_0_3833 <= _zz_dataOut_payload_0_3817;
    _zz_dataOut_payload_0_3834 <= _zz_dataOut_payload_0_3818;
    _zz_dataOut_payload_0_3835 <= _zz_dataOut_payload_0_3819;
    _zz_dataOut_payload_0_3836 <= _zz_dataOut_payload_0_3820;
    _zz_dataOut_payload_0_3837 <= _zz_dataOut_payload_0_3821;
    _zz_dataOut_payload_0_3838 <= _zz_dataOut_payload_0_3822;
    _zz_dataOut_payload_0_3839 <= _zz_dataOut_payload_0_3823;
    _zz_dataOut_payload_0_3884 <= (_zz_dataOut_payload_0_3882 ? _zz_dataOut_payload_0_3877 : _zz_dataOut_payload_0_3880);
    _zz_dataOut_payload_0_3885 <= (_zz_dataOut_payload_0_3882 ? _zz_dataOut_payload_0_3880 : _zz_dataOut_payload_0_3877);
    _zz_dataOut_payload_0_3886 <= (_zz_dataOut_payload_0_3883 ? _zz_dataOut_payload_0_3878 : _zz_dataOut_payload_0_3881);
    _zz_dataOut_payload_0_3887 <= (_zz_dataOut_payload_0_3883 ? _zz_dataOut_payload_0_3881 : _zz_dataOut_payload_0_3878);
    _zz_dataOut_payload_0_3896 <= (_zz_dataOut_payload_0_3894 ? _zz_dataOut_payload_0_3889 : _zz_dataOut_payload_0_3892);
    _zz_dataOut_payload_0_3897 <= (_zz_dataOut_payload_0_3894 ? _zz_dataOut_payload_0_3892 : _zz_dataOut_payload_0_3889);
    _zz_dataOut_payload_0_3898 <= (_zz_dataOut_payload_0_3895 ? _zz_dataOut_payload_0_3890 : _zz_dataOut_payload_0_3893);
    _zz_dataOut_payload_0_3899 <= (_zz_dataOut_payload_0_3895 ? _zz_dataOut_payload_0_3893 : _zz_dataOut_payload_0_3890);
    _zz_dataOut_payload_0_3900 <= _zz_dataOut_payload_0_3884;
    _zz_dataOut_payload_0_3901 <= _zz_dataOut_payload_0_3885;
    _zz_dataOut_payload_0_3902 <= _zz_dataOut_payload_0_3886;
    _zz_dataOut_payload_0_3903 <= _zz_dataOut_payload_0_3887;
    _zz_dataOut_payload_0_3904 <= _zz_dataOut_payload_0_3896;
    _zz_dataOut_payload_0_3905 <= _zz_dataOut_payload_0_3897;
    _zz_dataOut_payload_0_3906 <= _zz_dataOut_payload_0_3898;
    _zz_dataOut_payload_0_3907 <= _zz_dataOut_payload_0_3899;
    _zz_dataOut_payload_0_3928 <= (_zz_dataOut_payload_0_3926 ? _zz_dataOut_payload_0_3921 : _zz_dataOut_payload_0_3924);
    _zz_dataOut_payload_0_3929 <= (_zz_dataOut_payload_0_3926 ? _zz_dataOut_payload_0_3924 : _zz_dataOut_payload_0_3921);
    _zz_dataOut_payload_0_3930 <= (_zz_dataOut_payload_0_3927 ? _zz_dataOut_payload_0_3922 : _zz_dataOut_payload_0_3925);
    _zz_dataOut_payload_0_3931 <= (_zz_dataOut_payload_0_3927 ? _zz_dataOut_payload_0_3925 : _zz_dataOut_payload_0_3922);
    _zz_dataOut_payload_0_3940 <= (_zz_dataOut_payload_0_3938 ? _zz_dataOut_payload_0_3933 : _zz_dataOut_payload_0_3936);
    _zz_dataOut_payload_0_3941 <= (_zz_dataOut_payload_0_3938 ? _zz_dataOut_payload_0_3936 : _zz_dataOut_payload_0_3933);
    _zz_dataOut_payload_0_3942 <= (_zz_dataOut_payload_0_3939 ? _zz_dataOut_payload_0_3934 : _zz_dataOut_payload_0_3937);
    _zz_dataOut_payload_0_3943 <= (_zz_dataOut_payload_0_3939 ? _zz_dataOut_payload_0_3937 : _zz_dataOut_payload_0_3934);
    _zz_dataOut_payload_0_3944 <= _zz_dataOut_payload_0_3928;
    _zz_dataOut_payload_0_3945 <= _zz_dataOut_payload_0_3929;
    _zz_dataOut_payload_0_3946 <= _zz_dataOut_payload_0_3930;
    _zz_dataOut_payload_0_3947 <= _zz_dataOut_payload_0_3931;
    _zz_dataOut_payload_0_3948 <= _zz_dataOut_payload_0_3940;
    _zz_dataOut_payload_0_3949 <= _zz_dataOut_payload_0_3941;
    _zz_dataOut_payload_0_3950 <= _zz_dataOut_payload_0_3942;
    _zz_dataOut_payload_0_3951 <= _zz_dataOut_payload_0_3943;
    _zz_dataOut_payload_0_3952 <= _zz_dataOut_payload_0_3900;
    _zz_dataOut_payload_0_3953 <= _zz_dataOut_payload_0_3901;
    _zz_dataOut_payload_0_3954 <= _zz_dataOut_payload_0_3902;
    _zz_dataOut_payload_0_3955 <= _zz_dataOut_payload_0_3903;
    _zz_dataOut_payload_0_3956 <= _zz_dataOut_payload_0_3904;
    _zz_dataOut_payload_0_3957 <= _zz_dataOut_payload_0_3905;
    _zz_dataOut_payload_0_3958 <= _zz_dataOut_payload_0_3906;
    _zz_dataOut_payload_0_3959 <= _zz_dataOut_payload_0_3907;
    _zz_dataOut_payload_0_3960 <= _zz_dataOut_payload_0_3944;
    _zz_dataOut_payload_0_3961 <= _zz_dataOut_payload_0_3945;
    _zz_dataOut_payload_0_3962 <= _zz_dataOut_payload_0_3946;
    _zz_dataOut_payload_0_3963 <= _zz_dataOut_payload_0_3947;
    _zz_dataOut_payload_0_3964 <= _zz_dataOut_payload_0_3948;
    _zz_dataOut_payload_0_3965 <= _zz_dataOut_payload_0_3949;
    _zz_dataOut_payload_0_3966 <= _zz_dataOut_payload_0_3950;
    _zz_dataOut_payload_0_3967 <= _zz_dataOut_payload_0_3951;
    _zz_dataOut_payload_0_4012 <= (_zz_dataOut_payload_0_4010 ? _zz_dataOut_payload_0_4005 : _zz_dataOut_payload_0_4008);
    _zz_dataOut_payload_0_4013 <= (_zz_dataOut_payload_0_4010 ? _zz_dataOut_payload_0_4008 : _zz_dataOut_payload_0_4005);
    _zz_dataOut_payload_0_4014 <= (_zz_dataOut_payload_0_4011 ? _zz_dataOut_payload_0_4006 : _zz_dataOut_payload_0_4009);
    _zz_dataOut_payload_0_4015 <= (_zz_dataOut_payload_0_4011 ? _zz_dataOut_payload_0_4009 : _zz_dataOut_payload_0_4006);
    _zz_dataOut_payload_0_4024 <= (_zz_dataOut_payload_0_4022 ? _zz_dataOut_payload_0_4017 : _zz_dataOut_payload_0_4020);
    _zz_dataOut_payload_0_4025 <= (_zz_dataOut_payload_0_4022 ? _zz_dataOut_payload_0_4020 : _zz_dataOut_payload_0_4017);
    _zz_dataOut_payload_0_4026 <= (_zz_dataOut_payload_0_4023 ? _zz_dataOut_payload_0_4018 : _zz_dataOut_payload_0_4021);
    _zz_dataOut_payload_0_4027 <= (_zz_dataOut_payload_0_4023 ? _zz_dataOut_payload_0_4021 : _zz_dataOut_payload_0_4018);
    _zz_dataOut_payload_0_4028 <= _zz_dataOut_payload_0_4012;
    _zz_dataOut_payload_0_4029 <= _zz_dataOut_payload_0_4013;
    _zz_dataOut_payload_0_4030 <= _zz_dataOut_payload_0_4014;
    _zz_dataOut_payload_0_4031 <= _zz_dataOut_payload_0_4015;
    _zz_dataOut_payload_0_4032 <= _zz_dataOut_payload_0_4024;
    _zz_dataOut_payload_0_4033 <= _zz_dataOut_payload_0_4025;
    _zz_dataOut_payload_0_4034 <= _zz_dataOut_payload_0_4026;
    _zz_dataOut_payload_0_4035 <= _zz_dataOut_payload_0_4027;
    _zz_dataOut_payload_0_4056 <= (_zz_dataOut_payload_0_4054 ? _zz_dataOut_payload_0_4049 : _zz_dataOut_payload_0_4052);
    _zz_dataOut_payload_0_4057 <= (_zz_dataOut_payload_0_4054 ? _zz_dataOut_payload_0_4052 : _zz_dataOut_payload_0_4049);
    _zz_dataOut_payload_0_4058 <= (_zz_dataOut_payload_0_4055 ? _zz_dataOut_payload_0_4050 : _zz_dataOut_payload_0_4053);
    _zz_dataOut_payload_0_4059 <= (_zz_dataOut_payload_0_4055 ? _zz_dataOut_payload_0_4053 : _zz_dataOut_payload_0_4050);
    _zz_dataOut_payload_0_4068 <= (_zz_dataOut_payload_0_4066 ? _zz_dataOut_payload_0_4061 : _zz_dataOut_payload_0_4064);
    _zz_dataOut_payload_0_4069 <= (_zz_dataOut_payload_0_4066 ? _zz_dataOut_payload_0_4064 : _zz_dataOut_payload_0_4061);
    _zz_dataOut_payload_0_4070 <= (_zz_dataOut_payload_0_4067 ? _zz_dataOut_payload_0_4062 : _zz_dataOut_payload_0_4065);
    _zz_dataOut_payload_0_4071 <= (_zz_dataOut_payload_0_4067 ? _zz_dataOut_payload_0_4065 : _zz_dataOut_payload_0_4062);
    _zz_dataOut_payload_0_4072 <= _zz_dataOut_payload_0_4056;
    _zz_dataOut_payload_0_4073 <= _zz_dataOut_payload_0_4057;
    _zz_dataOut_payload_0_4074 <= _zz_dataOut_payload_0_4058;
    _zz_dataOut_payload_0_4075 <= _zz_dataOut_payload_0_4059;
    _zz_dataOut_payload_0_4076 <= _zz_dataOut_payload_0_4068;
    _zz_dataOut_payload_0_4077 <= _zz_dataOut_payload_0_4069;
    _zz_dataOut_payload_0_4078 <= _zz_dataOut_payload_0_4070;
    _zz_dataOut_payload_0_4079 <= _zz_dataOut_payload_0_4071;
    _zz_dataOut_payload_0_4080 <= _zz_dataOut_payload_0_4028;
    _zz_dataOut_payload_0_4081 <= _zz_dataOut_payload_0_4029;
    _zz_dataOut_payload_0_4082 <= _zz_dataOut_payload_0_4030;
    _zz_dataOut_payload_0_4083 <= _zz_dataOut_payload_0_4031;
    _zz_dataOut_payload_0_4084 <= _zz_dataOut_payload_0_4032;
    _zz_dataOut_payload_0_4085 <= _zz_dataOut_payload_0_4033;
    _zz_dataOut_payload_0_4086 <= _zz_dataOut_payload_0_4034;
    _zz_dataOut_payload_0_4087 <= _zz_dataOut_payload_0_4035;
    _zz_dataOut_payload_0_4088 <= _zz_dataOut_payload_0_4072;
    _zz_dataOut_payload_0_4089 <= _zz_dataOut_payload_0_4073;
    _zz_dataOut_payload_0_4090 <= _zz_dataOut_payload_0_4074;
    _zz_dataOut_payload_0_4091 <= _zz_dataOut_payload_0_4075;
    _zz_dataOut_payload_0_4092 <= _zz_dataOut_payload_0_4076;
    _zz_dataOut_payload_0_4093 <= _zz_dataOut_payload_0_4077;
    _zz_dataOut_payload_0_4094 <= _zz_dataOut_payload_0_4078;
    _zz_dataOut_payload_0_4095 <= _zz_dataOut_payload_0_4079;
    _zz_dataOut_payload_0_4140 <= (_zz_dataOut_payload_0_4138 ? _zz_dataOut_payload_0_4133 : _zz_dataOut_payload_0_4136);
    _zz_dataOut_payload_0_4141 <= (_zz_dataOut_payload_0_4138 ? _zz_dataOut_payload_0_4136 : _zz_dataOut_payload_0_4133);
    _zz_dataOut_payload_0_4142 <= (_zz_dataOut_payload_0_4139 ? _zz_dataOut_payload_0_4134 : _zz_dataOut_payload_0_4137);
    _zz_dataOut_payload_0_4143 <= (_zz_dataOut_payload_0_4139 ? _zz_dataOut_payload_0_4137 : _zz_dataOut_payload_0_4134);
    _zz_dataOut_payload_0_4152 <= (_zz_dataOut_payload_0_4150 ? _zz_dataOut_payload_0_4145 : _zz_dataOut_payload_0_4148);
    _zz_dataOut_payload_0_4153 <= (_zz_dataOut_payload_0_4150 ? _zz_dataOut_payload_0_4148 : _zz_dataOut_payload_0_4145);
    _zz_dataOut_payload_0_4154 <= (_zz_dataOut_payload_0_4151 ? _zz_dataOut_payload_0_4146 : _zz_dataOut_payload_0_4149);
    _zz_dataOut_payload_0_4155 <= (_zz_dataOut_payload_0_4151 ? _zz_dataOut_payload_0_4149 : _zz_dataOut_payload_0_4146);
    _zz_dataOut_payload_0_4156 <= _zz_dataOut_payload_0_4140;
    _zz_dataOut_payload_0_4157 <= _zz_dataOut_payload_0_4141;
    _zz_dataOut_payload_0_4158 <= _zz_dataOut_payload_0_4142;
    _zz_dataOut_payload_0_4159 <= _zz_dataOut_payload_0_4143;
    _zz_dataOut_payload_0_4160 <= _zz_dataOut_payload_0_4152;
    _zz_dataOut_payload_0_4161 <= _zz_dataOut_payload_0_4153;
    _zz_dataOut_payload_0_4162 <= _zz_dataOut_payload_0_4154;
    _zz_dataOut_payload_0_4163 <= _zz_dataOut_payload_0_4155;
    _zz_dataOut_payload_0_4184 <= (_zz_dataOut_payload_0_4182 ? _zz_dataOut_payload_0_4177 : _zz_dataOut_payload_0_4180);
    _zz_dataOut_payload_0_4185 <= (_zz_dataOut_payload_0_4182 ? _zz_dataOut_payload_0_4180 : _zz_dataOut_payload_0_4177);
    _zz_dataOut_payload_0_4186 <= (_zz_dataOut_payload_0_4183 ? _zz_dataOut_payload_0_4178 : _zz_dataOut_payload_0_4181);
    _zz_dataOut_payload_0_4187 <= (_zz_dataOut_payload_0_4183 ? _zz_dataOut_payload_0_4181 : _zz_dataOut_payload_0_4178);
    _zz_dataOut_payload_0_4196 <= (_zz_dataOut_payload_0_4194 ? _zz_dataOut_payload_0_4189 : _zz_dataOut_payload_0_4192);
    _zz_dataOut_payload_0_4197 <= (_zz_dataOut_payload_0_4194 ? _zz_dataOut_payload_0_4192 : _zz_dataOut_payload_0_4189);
    _zz_dataOut_payload_0_4198 <= (_zz_dataOut_payload_0_4195 ? _zz_dataOut_payload_0_4190 : _zz_dataOut_payload_0_4193);
    _zz_dataOut_payload_0_4199 <= (_zz_dataOut_payload_0_4195 ? _zz_dataOut_payload_0_4193 : _zz_dataOut_payload_0_4190);
    _zz_dataOut_payload_0_4200 <= _zz_dataOut_payload_0_4184;
    _zz_dataOut_payload_0_4201 <= _zz_dataOut_payload_0_4185;
    _zz_dataOut_payload_0_4202 <= _zz_dataOut_payload_0_4186;
    _zz_dataOut_payload_0_4203 <= _zz_dataOut_payload_0_4187;
    _zz_dataOut_payload_0_4204 <= _zz_dataOut_payload_0_4196;
    _zz_dataOut_payload_0_4205 <= _zz_dataOut_payload_0_4197;
    _zz_dataOut_payload_0_4206 <= _zz_dataOut_payload_0_4198;
    _zz_dataOut_payload_0_4207 <= _zz_dataOut_payload_0_4199;
    _zz_dataOut_payload_0_4208 <= _zz_dataOut_payload_0_4156;
    _zz_dataOut_payload_0_4209 <= _zz_dataOut_payload_0_4157;
    _zz_dataOut_payload_0_4210 <= _zz_dataOut_payload_0_4158;
    _zz_dataOut_payload_0_4211 <= _zz_dataOut_payload_0_4159;
    _zz_dataOut_payload_0_4212 <= _zz_dataOut_payload_0_4160;
    _zz_dataOut_payload_0_4213 <= _zz_dataOut_payload_0_4161;
    _zz_dataOut_payload_0_4214 <= _zz_dataOut_payload_0_4162;
    _zz_dataOut_payload_0_4215 <= _zz_dataOut_payload_0_4163;
    _zz_dataOut_payload_0_4216 <= _zz_dataOut_payload_0_4200;
    _zz_dataOut_payload_0_4217 <= _zz_dataOut_payload_0_4201;
    _zz_dataOut_payload_0_4218 <= _zz_dataOut_payload_0_4202;
    _zz_dataOut_payload_0_4219 <= _zz_dataOut_payload_0_4203;
    _zz_dataOut_payload_0_4220 <= _zz_dataOut_payload_0_4204;
    _zz_dataOut_payload_0_4221 <= _zz_dataOut_payload_0_4205;
    _zz_dataOut_payload_0_4222 <= _zz_dataOut_payload_0_4206;
    _zz_dataOut_payload_0_4223 <= _zz_dataOut_payload_0_4207;
    _zz_dataOut_payload_0_4268 <= (_zz_dataOut_payload_0_4266 ? _zz_dataOut_payload_0_4261 : _zz_dataOut_payload_0_4264);
    _zz_dataOut_payload_0_4269 <= (_zz_dataOut_payload_0_4266 ? _zz_dataOut_payload_0_4264 : _zz_dataOut_payload_0_4261);
    _zz_dataOut_payload_0_4270 <= (_zz_dataOut_payload_0_4267 ? _zz_dataOut_payload_0_4262 : _zz_dataOut_payload_0_4265);
    _zz_dataOut_payload_0_4271 <= (_zz_dataOut_payload_0_4267 ? _zz_dataOut_payload_0_4265 : _zz_dataOut_payload_0_4262);
    _zz_dataOut_payload_0_4280 <= (_zz_dataOut_payload_0_4278 ? _zz_dataOut_payload_0_4273 : _zz_dataOut_payload_0_4276);
    _zz_dataOut_payload_0_4281 <= (_zz_dataOut_payload_0_4278 ? _zz_dataOut_payload_0_4276 : _zz_dataOut_payload_0_4273);
    _zz_dataOut_payload_0_4282 <= (_zz_dataOut_payload_0_4279 ? _zz_dataOut_payload_0_4274 : _zz_dataOut_payload_0_4277);
    _zz_dataOut_payload_0_4283 <= (_zz_dataOut_payload_0_4279 ? _zz_dataOut_payload_0_4277 : _zz_dataOut_payload_0_4274);
    _zz_dataOut_payload_0_4284 <= _zz_dataOut_payload_0_4268;
    _zz_dataOut_payload_0_4285 <= _zz_dataOut_payload_0_4269;
    _zz_dataOut_payload_0_4286 <= _zz_dataOut_payload_0_4270;
    _zz_dataOut_payload_0_4287 <= _zz_dataOut_payload_0_4271;
    _zz_dataOut_payload_0_4288 <= _zz_dataOut_payload_0_4280;
    _zz_dataOut_payload_0_4289 <= _zz_dataOut_payload_0_4281;
    _zz_dataOut_payload_0_4290 <= _zz_dataOut_payload_0_4282;
    _zz_dataOut_payload_0_4291 <= _zz_dataOut_payload_0_4283;
    _zz_dataOut_payload_0_4312 <= (_zz_dataOut_payload_0_4310 ? _zz_dataOut_payload_0_4305 : _zz_dataOut_payload_0_4308);
    _zz_dataOut_payload_0_4313 <= (_zz_dataOut_payload_0_4310 ? _zz_dataOut_payload_0_4308 : _zz_dataOut_payload_0_4305);
    _zz_dataOut_payload_0_4314 <= (_zz_dataOut_payload_0_4311 ? _zz_dataOut_payload_0_4306 : _zz_dataOut_payload_0_4309);
    _zz_dataOut_payload_0_4315 <= (_zz_dataOut_payload_0_4311 ? _zz_dataOut_payload_0_4309 : _zz_dataOut_payload_0_4306);
    _zz_dataOut_payload_0_4324 <= (_zz_dataOut_payload_0_4322 ? _zz_dataOut_payload_0_4317 : _zz_dataOut_payload_0_4320);
    _zz_dataOut_payload_0_4325 <= (_zz_dataOut_payload_0_4322 ? _zz_dataOut_payload_0_4320 : _zz_dataOut_payload_0_4317);
    _zz_dataOut_payload_0_4326 <= (_zz_dataOut_payload_0_4323 ? _zz_dataOut_payload_0_4318 : _zz_dataOut_payload_0_4321);
    _zz_dataOut_payload_0_4327 <= (_zz_dataOut_payload_0_4323 ? _zz_dataOut_payload_0_4321 : _zz_dataOut_payload_0_4318);
    _zz_dataOut_payload_0_4328 <= _zz_dataOut_payload_0_4312;
    _zz_dataOut_payload_0_4329 <= _zz_dataOut_payload_0_4313;
    _zz_dataOut_payload_0_4330 <= _zz_dataOut_payload_0_4314;
    _zz_dataOut_payload_0_4331 <= _zz_dataOut_payload_0_4315;
    _zz_dataOut_payload_0_4332 <= _zz_dataOut_payload_0_4324;
    _zz_dataOut_payload_0_4333 <= _zz_dataOut_payload_0_4325;
    _zz_dataOut_payload_0_4334 <= _zz_dataOut_payload_0_4326;
    _zz_dataOut_payload_0_4335 <= _zz_dataOut_payload_0_4327;
    _zz_dataOut_payload_0_4336 <= _zz_dataOut_payload_0_4284;
    _zz_dataOut_payload_0_4337 <= _zz_dataOut_payload_0_4285;
    _zz_dataOut_payload_0_4338 <= _zz_dataOut_payload_0_4286;
    _zz_dataOut_payload_0_4339 <= _zz_dataOut_payload_0_4287;
    _zz_dataOut_payload_0_4340 <= _zz_dataOut_payload_0_4288;
    _zz_dataOut_payload_0_4341 <= _zz_dataOut_payload_0_4289;
    _zz_dataOut_payload_0_4342 <= _zz_dataOut_payload_0_4290;
    _zz_dataOut_payload_0_4343 <= _zz_dataOut_payload_0_4291;
    _zz_dataOut_payload_0_4344 <= _zz_dataOut_payload_0_4328;
    _zz_dataOut_payload_0_4345 <= _zz_dataOut_payload_0_4329;
    _zz_dataOut_payload_0_4346 <= _zz_dataOut_payload_0_4330;
    _zz_dataOut_payload_0_4347 <= _zz_dataOut_payload_0_4331;
    _zz_dataOut_payload_0_4348 <= _zz_dataOut_payload_0_4332;
    _zz_dataOut_payload_0_4349 <= _zz_dataOut_payload_0_4333;
    _zz_dataOut_payload_0_4350 <= _zz_dataOut_payload_0_4334;
    _zz_dataOut_payload_0_4351 <= _zz_dataOut_payload_0_4335;
    _zz_dataOut_payload_0_4396 <= (_zz_dataOut_payload_0_4394 ? _zz_dataOut_payload_0_4389 : _zz_dataOut_payload_0_4392);
    _zz_dataOut_payload_0_4397 <= (_zz_dataOut_payload_0_4394 ? _zz_dataOut_payload_0_4392 : _zz_dataOut_payload_0_4389);
    _zz_dataOut_payload_0_4398 <= (_zz_dataOut_payload_0_4395 ? _zz_dataOut_payload_0_4390 : _zz_dataOut_payload_0_4393);
    _zz_dataOut_payload_0_4399 <= (_zz_dataOut_payload_0_4395 ? _zz_dataOut_payload_0_4393 : _zz_dataOut_payload_0_4390);
    _zz_dataOut_payload_0_4408 <= (_zz_dataOut_payload_0_4406 ? _zz_dataOut_payload_0_4401 : _zz_dataOut_payload_0_4404);
    _zz_dataOut_payload_0_4409 <= (_zz_dataOut_payload_0_4406 ? _zz_dataOut_payload_0_4404 : _zz_dataOut_payload_0_4401);
    _zz_dataOut_payload_0_4410 <= (_zz_dataOut_payload_0_4407 ? _zz_dataOut_payload_0_4402 : _zz_dataOut_payload_0_4405);
    _zz_dataOut_payload_0_4411 <= (_zz_dataOut_payload_0_4407 ? _zz_dataOut_payload_0_4405 : _zz_dataOut_payload_0_4402);
    _zz_dataOut_payload_0_4412 <= _zz_dataOut_payload_0_4396;
    _zz_dataOut_payload_0_4413 <= _zz_dataOut_payload_0_4397;
    _zz_dataOut_payload_0_4414 <= _zz_dataOut_payload_0_4398;
    _zz_dataOut_payload_0_4415 <= _zz_dataOut_payload_0_4399;
    _zz_dataOut_payload_0_4416 <= _zz_dataOut_payload_0_4408;
    _zz_dataOut_payload_0_4417 <= _zz_dataOut_payload_0_4409;
    _zz_dataOut_payload_0_4418 <= _zz_dataOut_payload_0_4410;
    _zz_dataOut_payload_0_4419 <= _zz_dataOut_payload_0_4411;
    _zz_dataOut_payload_0_4440 <= (_zz_dataOut_payload_0_4438 ? _zz_dataOut_payload_0_4433 : _zz_dataOut_payload_0_4436);
    _zz_dataOut_payload_0_4441 <= (_zz_dataOut_payload_0_4438 ? _zz_dataOut_payload_0_4436 : _zz_dataOut_payload_0_4433);
    _zz_dataOut_payload_0_4442 <= (_zz_dataOut_payload_0_4439 ? _zz_dataOut_payload_0_4434 : _zz_dataOut_payload_0_4437);
    _zz_dataOut_payload_0_4443 <= (_zz_dataOut_payload_0_4439 ? _zz_dataOut_payload_0_4437 : _zz_dataOut_payload_0_4434);
    _zz_dataOut_payload_0_4452 <= (_zz_dataOut_payload_0_4450 ? _zz_dataOut_payload_0_4445 : _zz_dataOut_payload_0_4448);
    _zz_dataOut_payload_0_4453 <= (_zz_dataOut_payload_0_4450 ? _zz_dataOut_payload_0_4448 : _zz_dataOut_payload_0_4445);
    _zz_dataOut_payload_0_4454 <= (_zz_dataOut_payload_0_4451 ? _zz_dataOut_payload_0_4446 : _zz_dataOut_payload_0_4449);
    _zz_dataOut_payload_0_4455 <= (_zz_dataOut_payload_0_4451 ? _zz_dataOut_payload_0_4449 : _zz_dataOut_payload_0_4446);
    _zz_dataOut_payload_0_4456 <= _zz_dataOut_payload_0_4440;
    _zz_dataOut_payload_0_4457 <= _zz_dataOut_payload_0_4441;
    _zz_dataOut_payload_0_4458 <= _zz_dataOut_payload_0_4442;
    _zz_dataOut_payload_0_4459 <= _zz_dataOut_payload_0_4443;
    _zz_dataOut_payload_0_4460 <= _zz_dataOut_payload_0_4452;
    _zz_dataOut_payload_0_4461 <= _zz_dataOut_payload_0_4453;
    _zz_dataOut_payload_0_4462 <= _zz_dataOut_payload_0_4454;
    _zz_dataOut_payload_0_4463 <= _zz_dataOut_payload_0_4455;
    _zz_dataOut_payload_0_4464 <= _zz_dataOut_payload_0_4412;
    _zz_dataOut_payload_0_4465 <= _zz_dataOut_payload_0_4413;
    _zz_dataOut_payload_0_4466 <= _zz_dataOut_payload_0_4414;
    _zz_dataOut_payload_0_4467 <= _zz_dataOut_payload_0_4415;
    _zz_dataOut_payload_0_4468 <= _zz_dataOut_payload_0_4416;
    _zz_dataOut_payload_0_4469 <= _zz_dataOut_payload_0_4417;
    _zz_dataOut_payload_0_4470 <= _zz_dataOut_payload_0_4418;
    _zz_dataOut_payload_0_4471 <= _zz_dataOut_payload_0_4419;
    _zz_dataOut_payload_0_4472 <= _zz_dataOut_payload_0_4456;
    _zz_dataOut_payload_0_4473 <= _zz_dataOut_payload_0_4457;
    _zz_dataOut_payload_0_4474 <= _zz_dataOut_payload_0_4458;
    _zz_dataOut_payload_0_4475 <= _zz_dataOut_payload_0_4459;
    _zz_dataOut_payload_0_4476 <= _zz_dataOut_payload_0_4460;
    _zz_dataOut_payload_0_4477 <= _zz_dataOut_payload_0_4461;
    _zz_dataOut_payload_0_4478 <= _zz_dataOut_payload_0_4462;
    _zz_dataOut_payload_0_4479 <= _zz_dataOut_payload_0_4463;
    _zz_dataOut_payload_0_4524 <= (_zz_dataOut_payload_0_4522 ? _zz_dataOut_payload_0_4517 : _zz_dataOut_payload_0_4520);
    _zz_dataOut_payload_0_4525 <= (_zz_dataOut_payload_0_4522 ? _zz_dataOut_payload_0_4520 : _zz_dataOut_payload_0_4517);
    _zz_dataOut_payload_0_4526 <= (_zz_dataOut_payload_0_4523 ? _zz_dataOut_payload_0_4518 : _zz_dataOut_payload_0_4521);
    _zz_dataOut_payload_0_4527 <= (_zz_dataOut_payload_0_4523 ? _zz_dataOut_payload_0_4521 : _zz_dataOut_payload_0_4518);
    _zz_dataOut_payload_0_4536 <= (_zz_dataOut_payload_0_4534 ? _zz_dataOut_payload_0_4529 : _zz_dataOut_payload_0_4532);
    _zz_dataOut_payload_0_4537 <= (_zz_dataOut_payload_0_4534 ? _zz_dataOut_payload_0_4532 : _zz_dataOut_payload_0_4529);
    _zz_dataOut_payload_0_4538 <= (_zz_dataOut_payload_0_4535 ? _zz_dataOut_payload_0_4530 : _zz_dataOut_payload_0_4533);
    _zz_dataOut_payload_0_4539 <= (_zz_dataOut_payload_0_4535 ? _zz_dataOut_payload_0_4533 : _zz_dataOut_payload_0_4530);
    _zz_dataOut_payload_0_4540 <= _zz_dataOut_payload_0_4524;
    _zz_dataOut_payload_0_4541 <= _zz_dataOut_payload_0_4525;
    _zz_dataOut_payload_0_4542 <= _zz_dataOut_payload_0_4526;
    _zz_dataOut_payload_0_4543 <= _zz_dataOut_payload_0_4527;
    _zz_dataOut_payload_0_4544 <= _zz_dataOut_payload_0_4536;
    _zz_dataOut_payload_0_4545 <= _zz_dataOut_payload_0_4537;
    _zz_dataOut_payload_0_4546 <= _zz_dataOut_payload_0_4538;
    _zz_dataOut_payload_0_4547 <= _zz_dataOut_payload_0_4539;
    _zz_dataOut_payload_0_4568 <= (_zz_dataOut_payload_0_4566 ? _zz_dataOut_payload_0_4561 : _zz_dataOut_payload_0_4564);
    _zz_dataOut_payload_0_4569 <= (_zz_dataOut_payload_0_4566 ? _zz_dataOut_payload_0_4564 : _zz_dataOut_payload_0_4561);
    _zz_dataOut_payload_0_4570 <= (_zz_dataOut_payload_0_4567 ? _zz_dataOut_payload_0_4562 : _zz_dataOut_payload_0_4565);
    _zz_dataOut_payload_0_4571 <= (_zz_dataOut_payload_0_4567 ? _zz_dataOut_payload_0_4565 : _zz_dataOut_payload_0_4562);
    _zz_dataOut_payload_0_4580 <= (_zz_dataOut_payload_0_4578 ? _zz_dataOut_payload_0_4573 : _zz_dataOut_payload_0_4576);
    _zz_dataOut_payload_0_4581 <= (_zz_dataOut_payload_0_4578 ? _zz_dataOut_payload_0_4576 : _zz_dataOut_payload_0_4573);
    _zz_dataOut_payload_0_4582 <= (_zz_dataOut_payload_0_4579 ? _zz_dataOut_payload_0_4574 : _zz_dataOut_payload_0_4577);
    _zz_dataOut_payload_0_4583 <= (_zz_dataOut_payload_0_4579 ? _zz_dataOut_payload_0_4577 : _zz_dataOut_payload_0_4574);
    _zz_dataOut_payload_0_4584 <= _zz_dataOut_payload_0_4568;
    _zz_dataOut_payload_0_4585 <= _zz_dataOut_payload_0_4569;
    _zz_dataOut_payload_0_4586 <= _zz_dataOut_payload_0_4570;
    _zz_dataOut_payload_0_4587 <= _zz_dataOut_payload_0_4571;
    _zz_dataOut_payload_0_4588 <= _zz_dataOut_payload_0_4580;
    _zz_dataOut_payload_0_4589 <= _zz_dataOut_payload_0_4581;
    _zz_dataOut_payload_0_4590 <= _zz_dataOut_payload_0_4582;
    _zz_dataOut_payload_0_4591 <= _zz_dataOut_payload_0_4583;
    _zz_dataOut_payload_0_4592 <= _zz_dataOut_payload_0_4540;
    _zz_dataOut_payload_0_4593 <= _zz_dataOut_payload_0_4541;
    _zz_dataOut_payload_0_4594 <= _zz_dataOut_payload_0_4542;
    _zz_dataOut_payload_0_4595 <= _zz_dataOut_payload_0_4543;
    _zz_dataOut_payload_0_4596 <= _zz_dataOut_payload_0_4544;
    _zz_dataOut_payload_0_4597 <= _zz_dataOut_payload_0_4545;
    _zz_dataOut_payload_0_4598 <= _zz_dataOut_payload_0_4546;
    _zz_dataOut_payload_0_4599 <= _zz_dataOut_payload_0_4547;
    _zz_dataOut_payload_0_4600 <= _zz_dataOut_payload_0_4584;
    _zz_dataOut_payload_0_4601 <= _zz_dataOut_payload_0_4585;
    _zz_dataOut_payload_0_4602 <= _zz_dataOut_payload_0_4586;
    _zz_dataOut_payload_0_4603 <= _zz_dataOut_payload_0_4587;
    _zz_dataOut_payload_0_4604 <= _zz_dataOut_payload_0_4588;
    _zz_dataOut_payload_0_4605 <= _zz_dataOut_payload_0_4589;
    _zz_dataOut_payload_0_4606 <= _zz_dataOut_payload_0_4590;
    _zz_dataOut_payload_0_4607 <= _zz_dataOut_payload_0_4591;
    _zz_dataOut_payload_0_4652 <= (_zz_dataOut_payload_0_4650 ? _zz_dataOut_payload_0_4645 : _zz_dataOut_payload_0_4648);
    _zz_dataOut_payload_0_4653 <= (_zz_dataOut_payload_0_4650 ? _zz_dataOut_payload_0_4648 : _zz_dataOut_payload_0_4645);
    _zz_dataOut_payload_0_4654 <= (_zz_dataOut_payload_0_4651 ? _zz_dataOut_payload_0_4646 : _zz_dataOut_payload_0_4649);
    _zz_dataOut_payload_0_4655 <= (_zz_dataOut_payload_0_4651 ? _zz_dataOut_payload_0_4649 : _zz_dataOut_payload_0_4646);
    _zz_dataOut_payload_0_4664 <= (_zz_dataOut_payload_0_4662 ? _zz_dataOut_payload_0_4657 : _zz_dataOut_payload_0_4660);
    _zz_dataOut_payload_0_4665 <= (_zz_dataOut_payload_0_4662 ? _zz_dataOut_payload_0_4660 : _zz_dataOut_payload_0_4657);
    _zz_dataOut_payload_0_4666 <= (_zz_dataOut_payload_0_4663 ? _zz_dataOut_payload_0_4658 : _zz_dataOut_payload_0_4661);
    _zz_dataOut_payload_0_4667 <= (_zz_dataOut_payload_0_4663 ? _zz_dataOut_payload_0_4661 : _zz_dataOut_payload_0_4658);
    _zz_dataOut_payload_0_4668 <= _zz_dataOut_payload_0_4652;
    _zz_dataOut_payload_0_4669 <= _zz_dataOut_payload_0_4653;
    _zz_dataOut_payload_0_4670 <= _zz_dataOut_payload_0_4654;
    _zz_dataOut_payload_0_4671 <= _zz_dataOut_payload_0_4655;
    _zz_dataOut_payload_0_4672 <= _zz_dataOut_payload_0_4664;
    _zz_dataOut_payload_0_4673 <= _zz_dataOut_payload_0_4665;
    _zz_dataOut_payload_0_4674 <= _zz_dataOut_payload_0_4666;
    _zz_dataOut_payload_0_4675 <= _zz_dataOut_payload_0_4667;
    _zz_dataOut_payload_0_4696 <= (_zz_dataOut_payload_0_4694 ? _zz_dataOut_payload_0_4689 : _zz_dataOut_payload_0_4692);
    _zz_dataOut_payload_0_4697 <= (_zz_dataOut_payload_0_4694 ? _zz_dataOut_payload_0_4692 : _zz_dataOut_payload_0_4689);
    _zz_dataOut_payload_0_4698 <= (_zz_dataOut_payload_0_4695 ? _zz_dataOut_payload_0_4690 : _zz_dataOut_payload_0_4693);
    _zz_dataOut_payload_0_4699 <= (_zz_dataOut_payload_0_4695 ? _zz_dataOut_payload_0_4693 : _zz_dataOut_payload_0_4690);
    _zz_dataOut_payload_0_4708 <= (_zz_dataOut_payload_0_4706 ? _zz_dataOut_payload_0_4701 : _zz_dataOut_payload_0_4704);
    _zz_dataOut_payload_0_4709 <= (_zz_dataOut_payload_0_4706 ? _zz_dataOut_payload_0_4704 : _zz_dataOut_payload_0_4701);
    _zz_dataOut_payload_0_4710 <= (_zz_dataOut_payload_0_4707 ? _zz_dataOut_payload_0_4702 : _zz_dataOut_payload_0_4705);
    _zz_dataOut_payload_0_4711 <= (_zz_dataOut_payload_0_4707 ? _zz_dataOut_payload_0_4705 : _zz_dataOut_payload_0_4702);
    _zz_dataOut_payload_0_4712 <= _zz_dataOut_payload_0_4696;
    _zz_dataOut_payload_0_4713 <= _zz_dataOut_payload_0_4697;
    _zz_dataOut_payload_0_4714 <= _zz_dataOut_payload_0_4698;
    _zz_dataOut_payload_0_4715 <= _zz_dataOut_payload_0_4699;
    _zz_dataOut_payload_0_4716 <= _zz_dataOut_payload_0_4708;
    _zz_dataOut_payload_0_4717 <= _zz_dataOut_payload_0_4709;
    _zz_dataOut_payload_0_4718 <= _zz_dataOut_payload_0_4710;
    _zz_dataOut_payload_0_4719 <= _zz_dataOut_payload_0_4711;
    _zz_dataOut_payload_0_4720 <= _zz_dataOut_payload_0_4668;
    _zz_dataOut_payload_0_4721 <= _zz_dataOut_payload_0_4669;
    _zz_dataOut_payload_0_4722 <= _zz_dataOut_payload_0_4670;
    _zz_dataOut_payload_0_4723 <= _zz_dataOut_payload_0_4671;
    _zz_dataOut_payload_0_4724 <= _zz_dataOut_payload_0_4672;
    _zz_dataOut_payload_0_4725 <= _zz_dataOut_payload_0_4673;
    _zz_dataOut_payload_0_4726 <= _zz_dataOut_payload_0_4674;
    _zz_dataOut_payload_0_4727 <= _zz_dataOut_payload_0_4675;
    _zz_dataOut_payload_0_4728 <= _zz_dataOut_payload_0_4712;
    _zz_dataOut_payload_0_4729 <= _zz_dataOut_payload_0_4713;
    _zz_dataOut_payload_0_4730 <= _zz_dataOut_payload_0_4714;
    _zz_dataOut_payload_0_4731 <= _zz_dataOut_payload_0_4715;
    _zz_dataOut_payload_0_4732 <= _zz_dataOut_payload_0_4716;
    _zz_dataOut_payload_0_4733 <= _zz_dataOut_payload_0_4717;
    _zz_dataOut_payload_0_4734 <= _zz_dataOut_payload_0_4718;
    _zz_dataOut_payload_0_4735 <= _zz_dataOut_payload_0_4719;
    _zz_dataOut_payload_0_4780 <= (_zz_dataOut_payload_0_4778 ? _zz_dataOut_payload_0_4773 : _zz_dataOut_payload_0_4776);
    _zz_dataOut_payload_0_4781 <= (_zz_dataOut_payload_0_4778 ? _zz_dataOut_payload_0_4776 : _zz_dataOut_payload_0_4773);
    _zz_dataOut_payload_0_4782 <= (_zz_dataOut_payload_0_4779 ? _zz_dataOut_payload_0_4774 : _zz_dataOut_payload_0_4777);
    _zz_dataOut_payload_0_4783 <= (_zz_dataOut_payload_0_4779 ? _zz_dataOut_payload_0_4777 : _zz_dataOut_payload_0_4774);
    _zz_dataOut_payload_0_4792 <= (_zz_dataOut_payload_0_4790 ? _zz_dataOut_payload_0_4785 : _zz_dataOut_payload_0_4788);
    _zz_dataOut_payload_0_4793 <= (_zz_dataOut_payload_0_4790 ? _zz_dataOut_payload_0_4788 : _zz_dataOut_payload_0_4785);
    _zz_dataOut_payload_0_4794 <= (_zz_dataOut_payload_0_4791 ? _zz_dataOut_payload_0_4786 : _zz_dataOut_payload_0_4789);
    _zz_dataOut_payload_0_4795 <= (_zz_dataOut_payload_0_4791 ? _zz_dataOut_payload_0_4789 : _zz_dataOut_payload_0_4786);
    _zz_dataOut_payload_0_4796 <= _zz_dataOut_payload_0_4780;
    _zz_dataOut_payload_0_4797 <= _zz_dataOut_payload_0_4781;
    _zz_dataOut_payload_0_4798 <= _zz_dataOut_payload_0_4782;
    _zz_dataOut_payload_0_4799 <= _zz_dataOut_payload_0_4783;
    _zz_dataOut_payload_0_4800 <= _zz_dataOut_payload_0_4792;
    _zz_dataOut_payload_0_4801 <= _zz_dataOut_payload_0_4793;
    _zz_dataOut_payload_0_4802 <= _zz_dataOut_payload_0_4794;
    _zz_dataOut_payload_0_4803 <= _zz_dataOut_payload_0_4795;
    _zz_dataOut_payload_0_4824 <= (_zz_dataOut_payload_0_4822 ? _zz_dataOut_payload_0_4817 : _zz_dataOut_payload_0_4820);
    _zz_dataOut_payload_0_4825 <= (_zz_dataOut_payload_0_4822 ? _zz_dataOut_payload_0_4820 : _zz_dataOut_payload_0_4817);
    _zz_dataOut_payload_0_4826 <= (_zz_dataOut_payload_0_4823 ? _zz_dataOut_payload_0_4818 : _zz_dataOut_payload_0_4821);
    _zz_dataOut_payload_0_4827 <= (_zz_dataOut_payload_0_4823 ? _zz_dataOut_payload_0_4821 : _zz_dataOut_payload_0_4818);
    _zz_dataOut_payload_0_4836 <= (_zz_dataOut_payload_0_4834 ? _zz_dataOut_payload_0_4829 : _zz_dataOut_payload_0_4832);
    _zz_dataOut_payload_0_4837 <= (_zz_dataOut_payload_0_4834 ? _zz_dataOut_payload_0_4832 : _zz_dataOut_payload_0_4829);
    _zz_dataOut_payload_0_4838 <= (_zz_dataOut_payload_0_4835 ? _zz_dataOut_payload_0_4830 : _zz_dataOut_payload_0_4833);
    _zz_dataOut_payload_0_4839 <= (_zz_dataOut_payload_0_4835 ? _zz_dataOut_payload_0_4833 : _zz_dataOut_payload_0_4830);
    _zz_dataOut_payload_0_4840 <= _zz_dataOut_payload_0_4824;
    _zz_dataOut_payload_0_4841 <= _zz_dataOut_payload_0_4825;
    _zz_dataOut_payload_0_4842 <= _zz_dataOut_payload_0_4826;
    _zz_dataOut_payload_0_4843 <= _zz_dataOut_payload_0_4827;
    _zz_dataOut_payload_0_4844 <= _zz_dataOut_payload_0_4836;
    _zz_dataOut_payload_0_4845 <= _zz_dataOut_payload_0_4837;
    _zz_dataOut_payload_0_4846 <= _zz_dataOut_payload_0_4838;
    _zz_dataOut_payload_0_4847 <= _zz_dataOut_payload_0_4839;
    _zz_dataOut_payload_0_4848 <= _zz_dataOut_payload_0_4796;
    _zz_dataOut_payload_0_4849 <= _zz_dataOut_payload_0_4797;
    _zz_dataOut_payload_0_4850 <= _zz_dataOut_payload_0_4798;
    _zz_dataOut_payload_0_4851 <= _zz_dataOut_payload_0_4799;
    _zz_dataOut_payload_0_4852 <= _zz_dataOut_payload_0_4800;
    _zz_dataOut_payload_0_4853 <= _zz_dataOut_payload_0_4801;
    _zz_dataOut_payload_0_4854 <= _zz_dataOut_payload_0_4802;
    _zz_dataOut_payload_0_4855 <= _zz_dataOut_payload_0_4803;
    _zz_dataOut_payload_0_4856 <= _zz_dataOut_payload_0_4840;
    _zz_dataOut_payload_0_4857 <= _zz_dataOut_payload_0_4841;
    _zz_dataOut_payload_0_4858 <= _zz_dataOut_payload_0_4842;
    _zz_dataOut_payload_0_4859 <= _zz_dataOut_payload_0_4843;
    _zz_dataOut_payload_0_4860 <= _zz_dataOut_payload_0_4844;
    _zz_dataOut_payload_0_4861 <= _zz_dataOut_payload_0_4845;
    _zz_dataOut_payload_0_4862 <= _zz_dataOut_payload_0_4846;
    _zz_dataOut_payload_0_4863 <= _zz_dataOut_payload_0_4847;
    _zz_dataOut_payload_0_4908 <= (_zz_dataOut_payload_0_4906 ? _zz_dataOut_payload_0_4901 : _zz_dataOut_payload_0_4904);
    _zz_dataOut_payload_0_4909 <= (_zz_dataOut_payload_0_4906 ? _zz_dataOut_payload_0_4904 : _zz_dataOut_payload_0_4901);
    _zz_dataOut_payload_0_4910 <= (_zz_dataOut_payload_0_4907 ? _zz_dataOut_payload_0_4902 : _zz_dataOut_payload_0_4905);
    _zz_dataOut_payload_0_4911 <= (_zz_dataOut_payload_0_4907 ? _zz_dataOut_payload_0_4905 : _zz_dataOut_payload_0_4902);
    _zz_dataOut_payload_0_4920 <= (_zz_dataOut_payload_0_4918 ? _zz_dataOut_payload_0_4913 : _zz_dataOut_payload_0_4916);
    _zz_dataOut_payload_0_4921 <= (_zz_dataOut_payload_0_4918 ? _zz_dataOut_payload_0_4916 : _zz_dataOut_payload_0_4913);
    _zz_dataOut_payload_0_4922 <= (_zz_dataOut_payload_0_4919 ? _zz_dataOut_payload_0_4914 : _zz_dataOut_payload_0_4917);
    _zz_dataOut_payload_0_4923 <= (_zz_dataOut_payload_0_4919 ? _zz_dataOut_payload_0_4917 : _zz_dataOut_payload_0_4914);
    _zz_dataOut_payload_0_4924 <= _zz_dataOut_payload_0_4908;
    _zz_dataOut_payload_0_4925 <= _zz_dataOut_payload_0_4909;
    _zz_dataOut_payload_0_4926 <= _zz_dataOut_payload_0_4910;
    _zz_dataOut_payload_0_4927 <= _zz_dataOut_payload_0_4911;
    _zz_dataOut_payload_0_4928 <= _zz_dataOut_payload_0_4920;
    _zz_dataOut_payload_0_4929 <= _zz_dataOut_payload_0_4921;
    _zz_dataOut_payload_0_4930 <= _zz_dataOut_payload_0_4922;
    _zz_dataOut_payload_0_4931 <= _zz_dataOut_payload_0_4923;
    _zz_dataOut_payload_0_4952 <= (_zz_dataOut_payload_0_4950 ? _zz_dataOut_payload_0_4945 : _zz_dataOut_payload_0_4948);
    _zz_dataOut_payload_0_4953 <= (_zz_dataOut_payload_0_4950 ? _zz_dataOut_payload_0_4948 : _zz_dataOut_payload_0_4945);
    _zz_dataOut_payload_0_4954 <= (_zz_dataOut_payload_0_4951 ? _zz_dataOut_payload_0_4946 : _zz_dataOut_payload_0_4949);
    _zz_dataOut_payload_0_4955 <= (_zz_dataOut_payload_0_4951 ? _zz_dataOut_payload_0_4949 : _zz_dataOut_payload_0_4946);
    _zz_dataOut_payload_0_4964 <= (_zz_dataOut_payload_0_4962 ? _zz_dataOut_payload_0_4957 : _zz_dataOut_payload_0_4960);
    _zz_dataOut_payload_0_4965 <= (_zz_dataOut_payload_0_4962 ? _zz_dataOut_payload_0_4960 : _zz_dataOut_payload_0_4957);
    _zz_dataOut_payload_0_4966 <= (_zz_dataOut_payload_0_4963 ? _zz_dataOut_payload_0_4958 : _zz_dataOut_payload_0_4961);
    _zz_dataOut_payload_0_4967 <= (_zz_dataOut_payload_0_4963 ? _zz_dataOut_payload_0_4961 : _zz_dataOut_payload_0_4958);
    _zz_dataOut_payload_0_4968 <= _zz_dataOut_payload_0_4952;
    _zz_dataOut_payload_0_4969 <= _zz_dataOut_payload_0_4953;
    _zz_dataOut_payload_0_4970 <= _zz_dataOut_payload_0_4954;
    _zz_dataOut_payload_0_4971 <= _zz_dataOut_payload_0_4955;
    _zz_dataOut_payload_0_4972 <= _zz_dataOut_payload_0_4964;
    _zz_dataOut_payload_0_4973 <= _zz_dataOut_payload_0_4965;
    _zz_dataOut_payload_0_4974 <= _zz_dataOut_payload_0_4966;
    _zz_dataOut_payload_0_4975 <= _zz_dataOut_payload_0_4967;
    _zz_dataOut_payload_0_4976 <= _zz_dataOut_payload_0_4924;
    _zz_dataOut_payload_0_4977 <= _zz_dataOut_payload_0_4925;
    _zz_dataOut_payload_0_4978 <= _zz_dataOut_payload_0_4926;
    _zz_dataOut_payload_0_4979 <= _zz_dataOut_payload_0_4927;
    _zz_dataOut_payload_0_4980 <= _zz_dataOut_payload_0_4928;
    _zz_dataOut_payload_0_4981 <= _zz_dataOut_payload_0_4929;
    _zz_dataOut_payload_0_4982 <= _zz_dataOut_payload_0_4930;
    _zz_dataOut_payload_0_4983 <= _zz_dataOut_payload_0_4931;
    _zz_dataOut_payload_0_4984 <= _zz_dataOut_payload_0_4968;
    _zz_dataOut_payload_0_4985 <= _zz_dataOut_payload_0_4969;
    _zz_dataOut_payload_0_4986 <= _zz_dataOut_payload_0_4970;
    _zz_dataOut_payload_0_4987 <= _zz_dataOut_payload_0_4971;
    _zz_dataOut_payload_0_4988 <= _zz_dataOut_payload_0_4972;
    _zz_dataOut_payload_0_4989 <= _zz_dataOut_payload_0_4973;
    _zz_dataOut_payload_0_4990 <= _zz_dataOut_payload_0_4974;
    _zz_dataOut_payload_0_4991 <= _zz_dataOut_payload_0_4975;
    _zz_dataOut_payload_0_5036 <= (_zz_dataOut_payload_0_5034 ? _zz_dataOut_payload_0_5029 : _zz_dataOut_payload_0_5032);
    _zz_dataOut_payload_0_5037 <= (_zz_dataOut_payload_0_5034 ? _zz_dataOut_payload_0_5032 : _zz_dataOut_payload_0_5029);
    _zz_dataOut_payload_0_5038 <= (_zz_dataOut_payload_0_5035 ? _zz_dataOut_payload_0_5030 : _zz_dataOut_payload_0_5033);
    _zz_dataOut_payload_0_5039 <= (_zz_dataOut_payload_0_5035 ? _zz_dataOut_payload_0_5033 : _zz_dataOut_payload_0_5030);
    _zz_dataOut_payload_0_5048 <= (_zz_dataOut_payload_0_5046 ? _zz_dataOut_payload_0_5041 : _zz_dataOut_payload_0_5044);
    _zz_dataOut_payload_0_5049 <= (_zz_dataOut_payload_0_5046 ? _zz_dataOut_payload_0_5044 : _zz_dataOut_payload_0_5041);
    _zz_dataOut_payload_0_5050 <= (_zz_dataOut_payload_0_5047 ? _zz_dataOut_payload_0_5042 : _zz_dataOut_payload_0_5045);
    _zz_dataOut_payload_0_5051 <= (_zz_dataOut_payload_0_5047 ? _zz_dataOut_payload_0_5045 : _zz_dataOut_payload_0_5042);
    _zz_dataOut_payload_0_5052 <= _zz_dataOut_payload_0_5036;
    _zz_dataOut_payload_0_5053 <= _zz_dataOut_payload_0_5037;
    _zz_dataOut_payload_0_5054 <= _zz_dataOut_payload_0_5038;
    _zz_dataOut_payload_0_5055 <= _zz_dataOut_payload_0_5039;
    _zz_dataOut_payload_0_5056 <= _zz_dataOut_payload_0_5048;
    _zz_dataOut_payload_0_5057 <= _zz_dataOut_payload_0_5049;
    _zz_dataOut_payload_0_5058 <= _zz_dataOut_payload_0_5050;
    _zz_dataOut_payload_0_5059 <= _zz_dataOut_payload_0_5051;
    _zz_dataOut_payload_0_5080 <= (_zz_dataOut_payload_0_5078 ? _zz_dataOut_payload_0_5073 : _zz_dataOut_payload_0_5076);
    _zz_dataOut_payload_0_5081 <= (_zz_dataOut_payload_0_5078 ? _zz_dataOut_payload_0_5076 : _zz_dataOut_payload_0_5073);
    _zz_dataOut_payload_0_5082 <= (_zz_dataOut_payload_0_5079 ? _zz_dataOut_payload_0_5074 : _zz_dataOut_payload_0_5077);
    _zz_dataOut_payload_0_5083 <= (_zz_dataOut_payload_0_5079 ? _zz_dataOut_payload_0_5077 : _zz_dataOut_payload_0_5074);
    _zz_dataOut_payload_0_5092 <= (_zz_dataOut_payload_0_5090 ? _zz_dataOut_payload_0_5085 : _zz_dataOut_payload_0_5088);
    _zz_dataOut_payload_0_5093 <= (_zz_dataOut_payload_0_5090 ? _zz_dataOut_payload_0_5088 : _zz_dataOut_payload_0_5085);
    _zz_dataOut_payload_0_5094 <= (_zz_dataOut_payload_0_5091 ? _zz_dataOut_payload_0_5086 : _zz_dataOut_payload_0_5089);
    _zz_dataOut_payload_0_5095 <= (_zz_dataOut_payload_0_5091 ? _zz_dataOut_payload_0_5089 : _zz_dataOut_payload_0_5086);
    _zz_dataOut_payload_0_5096 <= _zz_dataOut_payload_0_5080;
    _zz_dataOut_payload_0_5097 <= _zz_dataOut_payload_0_5081;
    _zz_dataOut_payload_0_5098 <= _zz_dataOut_payload_0_5082;
    _zz_dataOut_payload_0_5099 <= _zz_dataOut_payload_0_5083;
    _zz_dataOut_payload_0_5100 <= _zz_dataOut_payload_0_5092;
    _zz_dataOut_payload_0_5101 <= _zz_dataOut_payload_0_5093;
    _zz_dataOut_payload_0_5102 <= _zz_dataOut_payload_0_5094;
    _zz_dataOut_payload_0_5103 <= _zz_dataOut_payload_0_5095;
    _zz_dataOut_payload_0_5104 <= _zz_dataOut_payload_0_5052;
    _zz_dataOut_payload_0_5105 <= _zz_dataOut_payload_0_5053;
    _zz_dataOut_payload_0_5106 <= _zz_dataOut_payload_0_5054;
    _zz_dataOut_payload_0_5107 <= _zz_dataOut_payload_0_5055;
    _zz_dataOut_payload_0_5108 <= _zz_dataOut_payload_0_5056;
    _zz_dataOut_payload_0_5109 <= _zz_dataOut_payload_0_5057;
    _zz_dataOut_payload_0_5110 <= _zz_dataOut_payload_0_5058;
    _zz_dataOut_payload_0_5111 <= _zz_dataOut_payload_0_5059;
    _zz_dataOut_payload_0_5112 <= _zz_dataOut_payload_0_5096;
    _zz_dataOut_payload_0_5113 <= _zz_dataOut_payload_0_5097;
    _zz_dataOut_payload_0_5114 <= _zz_dataOut_payload_0_5098;
    _zz_dataOut_payload_0_5115 <= _zz_dataOut_payload_0_5099;
    _zz_dataOut_payload_0_5116 <= _zz_dataOut_payload_0_5100;
    _zz_dataOut_payload_0_5117 <= _zz_dataOut_payload_0_5101;
    _zz_dataOut_payload_0_5118 <= _zz_dataOut_payload_0_5102;
    _zz_dataOut_payload_0_5119 <= _zz_dataOut_payload_0_5103;
    _zz_dataOut_payload_0_5120 <= _zz_dataOut_payload_0_3184;
    _zz_dataOut_payload_0_5121 <= _zz_dataOut_payload_0_3185;
    _zz_dataOut_payload_0_5122 <= _zz_dataOut_payload_0_3186;
    _zz_dataOut_payload_0_5123 <= _zz_dataOut_payload_0_3187;
    _zz_dataOut_payload_0_5124 <= _zz_dataOut_payload_0_3188;
    _zz_dataOut_payload_0_5125 <= _zz_dataOut_payload_0_3189;
    _zz_dataOut_payload_0_5126 <= _zz_dataOut_payload_0_3190;
    _zz_dataOut_payload_0_5127 <= _zz_dataOut_payload_0_3191;
    _zz_dataOut_payload_0_5128 <= _zz_dataOut_payload_0_3192;
    _zz_dataOut_payload_0_5129 <= _zz_dataOut_payload_0_3193;
    _zz_dataOut_payload_0_5130 <= _zz_dataOut_payload_0_3194;
    _zz_dataOut_payload_0_5131 <= _zz_dataOut_payload_0_3195;
    _zz_dataOut_payload_0_5132 <= _zz_dataOut_payload_0_3196;
    _zz_dataOut_payload_0_5133 <= _zz_dataOut_payload_0_3197;
    _zz_dataOut_payload_0_5134 <= _zz_dataOut_payload_0_3198;
    _zz_dataOut_payload_0_5135 <= _zz_dataOut_payload_0_3199;
    _zz_dataOut_payload_0_5136 <= _zz_dataOut_payload_0_3312;
    _zz_dataOut_payload_0_5137 <= _zz_dataOut_payload_0_3313;
    _zz_dataOut_payload_0_5138 <= _zz_dataOut_payload_0_3314;
    _zz_dataOut_payload_0_5139 <= _zz_dataOut_payload_0_3315;
    _zz_dataOut_payload_0_5140 <= _zz_dataOut_payload_0_3316;
    _zz_dataOut_payload_0_5141 <= _zz_dataOut_payload_0_3317;
    _zz_dataOut_payload_0_5142 <= _zz_dataOut_payload_0_3318;
    _zz_dataOut_payload_0_5143 <= _zz_dataOut_payload_0_3319;
    _zz_dataOut_payload_0_5144 <= _zz_dataOut_payload_0_3320;
    _zz_dataOut_payload_0_5145 <= _zz_dataOut_payload_0_3321;
    _zz_dataOut_payload_0_5146 <= _zz_dataOut_payload_0_3322;
    _zz_dataOut_payload_0_5147 <= _zz_dataOut_payload_0_3323;
    _zz_dataOut_payload_0_5148 <= _zz_dataOut_payload_0_3324;
    _zz_dataOut_payload_0_5149 <= _zz_dataOut_payload_0_3325;
    _zz_dataOut_payload_0_5150 <= _zz_dataOut_payload_0_3326;
    _zz_dataOut_payload_0_5151 <= _zz_dataOut_payload_0_3327;
    _zz_dataOut_payload_0_5152 <= _zz_dataOut_payload_0_3440;
    _zz_dataOut_payload_0_5153 <= _zz_dataOut_payload_0_3441;
    _zz_dataOut_payload_0_5154 <= _zz_dataOut_payload_0_3442;
    _zz_dataOut_payload_0_5155 <= _zz_dataOut_payload_0_3443;
    _zz_dataOut_payload_0_5156 <= _zz_dataOut_payload_0_3444;
    _zz_dataOut_payload_0_5157 <= _zz_dataOut_payload_0_3445;
    _zz_dataOut_payload_0_5158 <= _zz_dataOut_payload_0_3446;
    _zz_dataOut_payload_0_5159 <= _zz_dataOut_payload_0_3447;
    _zz_dataOut_payload_0_5160 <= _zz_dataOut_payload_0_3448;
    _zz_dataOut_payload_0_5161 <= _zz_dataOut_payload_0_3449;
    _zz_dataOut_payload_0_5162 <= _zz_dataOut_payload_0_3450;
    _zz_dataOut_payload_0_5163 <= _zz_dataOut_payload_0_3451;
    _zz_dataOut_payload_0_5164 <= _zz_dataOut_payload_0_3452;
    _zz_dataOut_payload_0_5165 <= _zz_dataOut_payload_0_3453;
    _zz_dataOut_payload_0_5166 <= _zz_dataOut_payload_0_3454;
    _zz_dataOut_payload_0_5167 <= _zz_dataOut_payload_0_3455;
    _zz_dataOut_payload_0_5168 <= _zz_dataOut_payload_0_3568;
    _zz_dataOut_payload_0_5169 <= _zz_dataOut_payload_0_3569;
    _zz_dataOut_payload_0_5170 <= _zz_dataOut_payload_0_3570;
    _zz_dataOut_payload_0_5171 <= _zz_dataOut_payload_0_3571;
    _zz_dataOut_payload_0_5172 <= _zz_dataOut_payload_0_3572;
    _zz_dataOut_payload_0_5173 <= _zz_dataOut_payload_0_3573;
    _zz_dataOut_payload_0_5174 <= _zz_dataOut_payload_0_3574;
    _zz_dataOut_payload_0_5175 <= _zz_dataOut_payload_0_3575;
    _zz_dataOut_payload_0_5176 <= _zz_dataOut_payload_0_3576;
    _zz_dataOut_payload_0_5177 <= _zz_dataOut_payload_0_3577;
    _zz_dataOut_payload_0_5178 <= _zz_dataOut_payload_0_3578;
    _zz_dataOut_payload_0_5179 <= _zz_dataOut_payload_0_3579;
    _zz_dataOut_payload_0_5180 <= _zz_dataOut_payload_0_3580;
    _zz_dataOut_payload_0_5181 <= _zz_dataOut_payload_0_3581;
    _zz_dataOut_payload_0_5182 <= _zz_dataOut_payload_0_3582;
    _zz_dataOut_payload_0_5183 <= _zz_dataOut_payload_0_3583;
    _zz_dataOut_payload_0_5184 <= _zz_dataOut_payload_0_3696;
    _zz_dataOut_payload_0_5185 <= _zz_dataOut_payload_0_3697;
    _zz_dataOut_payload_0_5186 <= _zz_dataOut_payload_0_3698;
    _zz_dataOut_payload_0_5187 <= _zz_dataOut_payload_0_3699;
    _zz_dataOut_payload_0_5188 <= _zz_dataOut_payload_0_3700;
    _zz_dataOut_payload_0_5189 <= _zz_dataOut_payload_0_3701;
    _zz_dataOut_payload_0_5190 <= _zz_dataOut_payload_0_3702;
    _zz_dataOut_payload_0_5191 <= _zz_dataOut_payload_0_3703;
    _zz_dataOut_payload_0_5192 <= _zz_dataOut_payload_0_3704;
    _zz_dataOut_payload_0_5193 <= _zz_dataOut_payload_0_3705;
    _zz_dataOut_payload_0_5194 <= _zz_dataOut_payload_0_3706;
    _zz_dataOut_payload_0_5195 <= _zz_dataOut_payload_0_3707;
    _zz_dataOut_payload_0_5196 <= _zz_dataOut_payload_0_3708;
    _zz_dataOut_payload_0_5197 <= _zz_dataOut_payload_0_3709;
    _zz_dataOut_payload_0_5198 <= _zz_dataOut_payload_0_3710;
    _zz_dataOut_payload_0_5199 <= _zz_dataOut_payload_0_3711;
    _zz_dataOut_payload_0_5200 <= _zz_dataOut_payload_0_3824;
    _zz_dataOut_payload_0_5201 <= _zz_dataOut_payload_0_3825;
    _zz_dataOut_payload_0_5202 <= _zz_dataOut_payload_0_3826;
    _zz_dataOut_payload_0_5203 <= _zz_dataOut_payload_0_3827;
    _zz_dataOut_payload_0_5204 <= _zz_dataOut_payload_0_3828;
    _zz_dataOut_payload_0_5205 <= _zz_dataOut_payload_0_3829;
    _zz_dataOut_payload_0_5206 <= _zz_dataOut_payload_0_3830;
    _zz_dataOut_payload_0_5207 <= _zz_dataOut_payload_0_3831;
    _zz_dataOut_payload_0_5208 <= _zz_dataOut_payload_0_3832;
    _zz_dataOut_payload_0_5209 <= _zz_dataOut_payload_0_3833;
    _zz_dataOut_payload_0_5210 <= _zz_dataOut_payload_0_3834;
    _zz_dataOut_payload_0_5211 <= _zz_dataOut_payload_0_3835;
    _zz_dataOut_payload_0_5212 <= _zz_dataOut_payload_0_3836;
    _zz_dataOut_payload_0_5213 <= _zz_dataOut_payload_0_3837;
    _zz_dataOut_payload_0_5214 <= _zz_dataOut_payload_0_3838;
    _zz_dataOut_payload_0_5215 <= _zz_dataOut_payload_0_3839;
    _zz_dataOut_payload_0_5216 <= _zz_dataOut_payload_0_3952;
    _zz_dataOut_payload_0_5217 <= _zz_dataOut_payload_0_3953;
    _zz_dataOut_payload_0_5218 <= _zz_dataOut_payload_0_3954;
    _zz_dataOut_payload_0_5219 <= _zz_dataOut_payload_0_3955;
    _zz_dataOut_payload_0_5220 <= _zz_dataOut_payload_0_3956;
    _zz_dataOut_payload_0_5221 <= _zz_dataOut_payload_0_3957;
    _zz_dataOut_payload_0_5222 <= _zz_dataOut_payload_0_3958;
    _zz_dataOut_payload_0_5223 <= _zz_dataOut_payload_0_3959;
    _zz_dataOut_payload_0_5224 <= _zz_dataOut_payload_0_3960;
    _zz_dataOut_payload_0_5225 <= _zz_dataOut_payload_0_3961;
    _zz_dataOut_payload_0_5226 <= _zz_dataOut_payload_0_3962;
    _zz_dataOut_payload_0_5227 <= _zz_dataOut_payload_0_3963;
    _zz_dataOut_payload_0_5228 <= _zz_dataOut_payload_0_3964;
    _zz_dataOut_payload_0_5229 <= _zz_dataOut_payload_0_3965;
    _zz_dataOut_payload_0_5230 <= _zz_dataOut_payload_0_3966;
    _zz_dataOut_payload_0_5231 <= _zz_dataOut_payload_0_3967;
    _zz_dataOut_payload_0_5232 <= _zz_dataOut_payload_0_4080;
    _zz_dataOut_payload_0_5233 <= _zz_dataOut_payload_0_4081;
    _zz_dataOut_payload_0_5234 <= _zz_dataOut_payload_0_4082;
    _zz_dataOut_payload_0_5235 <= _zz_dataOut_payload_0_4083;
    _zz_dataOut_payload_0_5236 <= _zz_dataOut_payload_0_4084;
    _zz_dataOut_payload_0_5237 <= _zz_dataOut_payload_0_4085;
    _zz_dataOut_payload_0_5238 <= _zz_dataOut_payload_0_4086;
    _zz_dataOut_payload_0_5239 <= _zz_dataOut_payload_0_4087;
    _zz_dataOut_payload_0_5240 <= _zz_dataOut_payload_0_4088;
    _zz_dataOut_payload_0_5241 <= _zz_dataOut_payload_0_4089;
    _zz_dataOut_payload_0_5242 <= _zz_dataOut_payload_0_4090;
    _zz_dataOut_payload_0_5243 <= _zz_dataOut_payload_0_4091;
    _zz_dataOut_payload_0_5244 <= _zz_dataOut_payload_0_4092;
    _zz_dataOut_payload_0_5245 <= _zz_dataOut_payload_0_4093;
    _zz_dataOut_payload_0_5246 <= _zz_dataOut_payload_0_4094;
    _zz_dataOut_payload_0_5247 <= _zz_dataOut_payload_0_4095;
    _zz_dataOut_payload_0_5248 <= _zz_dataOut_payload_0_4208;
    _zz_dataOut_payload_0_5249 <= _zz_dataOut_payload_0_4209;
    _zz_dataOut_payload_0_5250 <= _zz_dataOut_payload_0_4210;
    _zz_dataOut_payload_0_5251 <= _zz_dataOut_payload_0_4211;
    _zz_dataOut_payload_0_5252 <= _zz_dataOut_payload_0_4212;
    _zz_dataOut_payload_0_5253 <= _zz_dataOut_payload_0_4213;
    _zz_dataOut_payload_0_5254 <= _zz_dataOut_payload_0_4214;
    _zz_dataOut_payload_0_5255 <= _zz_dataOut_payload_0_4215;
    _zz_dataOut_payload_0_5256 <= _zz_dataOut_payload_0_4216;
    _zz_dataOut_payload_0_5257 <= _zz_dataOut_payload_0_4217;
    _zz_dataOut_payload_0_5258 <= _zz_dataOut_payload_0_4218;
    _zz_dataOut_payload_0_5259 <= _zz_dataOut_payload_0_4219;
    _zz_dataOut_payload_0_5260 <= _zz_dataOut_payload_0_4220;
    _zz_dataOut_payload_0_5261 <= _zz_dataOut_payload_0_4221;
    _zz_dataOut_payload_0_5262 <= _zz_dataOut_payload_0_4222;
    _zz_dataOut_payload_0_5263 <= _zz_dataOut_payload_0_4223;
    _zz_dataOut_payload_0_5264 <= _zz_dataOut_payload_0_4336;
    _zz_dataOut_payload_0_5265 <= _zz_dataOut_payload_0_4337;
    _zz_dataOut_payload_0_5266 <= _zz_dataOut_payload_0_4338;
    _zz_dataOut_payload_0_5267 <= _zz_dataOut_payload_0_4339;
    _zz_dataOut_payload_0_5268 <= _zz_dataOut_payload_0_4340;
    _zz_dataOut_payload_0_5269 <= _zz_dataOut_payload_0_4341;
    _zz_dataOut_payload_0_5270 <= _zz_dataOut_payload_0_4342;
    _zz_dataOut_payload_0_5271 <= _zz_dataOut_payload_0_4343;
    _zz_dataOut_payload_0_5272 <= _zz_dataOut_payload_0_4344;
    _zz_dataOut_payload_0_5273 <= _zz_dataOut_payload_0_4345;
    _zz_dataOut_payload_0_5274 <= _zz_dataOut_payload_0_4346;
    _zz_dataOut_payload_0_5275 <= _zz_dataOut_payload_0_4347;
    _zz_dataOut_payload_0_5276 <= _zz_dataOut_payload_0_4348;
    _zz_dataOut_payload_0_5277 <= _zz_dataOut_payload_0_4349;
    _zz_dataOut_payload_0_5278 <= _zz_dataOut_payload_0_4350;
    _zz_dataOut_payload_0_5279 <= _zz_dataOut_payload_0_4351;
    _zz_dataOut_payload_0_5280 <= _zz_dataOut_payload_0_4464;
    _zz_dataOut_payload_0_5281 <= _zz_dataOut_payload_0_4465;
    _zz_dataOut_payload_0_5282 <= _zz_dataOut_payload_0_4466;
    _zz_dataOut_payload_0_5283 <= _zz_dataOut_payload_0_4467;
    _zz_dataOut_payload_0_5284 <= _zz_dataOut_payload_0_4468;
    _zz_dataOut_payload_0_5285 <= _zz_dataOut_payload_0_4469;
    _zz_dataOut_payload_0_5286 <= _zz_dataOut_payload_0_4470;
    _zz_dataOut_payload_0_5287 <= _zz_dataOut_payload_0_4471;
    _zz_dataOut_payload_0_5288 <= _zz_dataOut_payload_0_4472;
    _zz_dataOut_payload_0_5289 <= _zz_dataOut_payload_0_4473;
    _zz_dataOut_payload_0_5290 <= _zz_dataOut_payload_0_4474;
    _zz_dataOut_payload_0_5291 <= _zz_dataOut_payload_0_4475;
    _zz_dataOut_payload_0_5292 <= _zz_dataOut_payload_0_4476;
    _zz_dataOut_payload_0_5293 <= _zz_dataOut_payload_0_4477;
    _zz_dataOut_payload_0_5294 <= _zz_dataOut_payload_0_4478;
    _zz_dataOut_payload_0_5295 <= _zz_dataOut_payload_0_4479;
    _zz_dataOut_payload_0_5296 <= _zz_dataOut_payload_0_4592;
    _zz_dataOut_payload_0_5297 <= _zz_dataOut_payload_0_4593;
    _zz_dataOut_payload_0_5298 <= _zz_dataOut_payload_0_4594;
    _zz_dataOut_payload_0_5299 <= _zz_dataOut_payload_0_4595;
    _zz_dataOut_payload_0_5300 <= _zz_dataOut_payload_0_4596;
    _zz_dataOut_payload_0_5301 <= _zz_dataOut_payload_0_4597;
    _zz_dataOut_payload_0_5302 <= _zz_dataOut_payload_0_4598;
    _zz_dataOut_payload_0_5303 <= _zz_dataOut_payload_0_4599;
    _zz_dataOut_payload_0_5304 <= _zz_dataOut_payload_0_4600;
    _zz_dataOut_payload_0_5305 <= _zz_dataOut_payload_0_4601;
    _zz_dataOut_payload_0_5306 <= _zz_dataOut_payload_0_4602;
    _zz_dataOut_payload_0_5307 <= _zz_dataOut_payload_0_4603;
    _zz_dataOut_payload_0_5308 <= _zz_dataOut_payload_0_4604;
    _zz_dataOut_payload_0_5309 <= _zz_dataOut_payload_0_4605;
    _zz_dataOut_payload_0_5310 <= _zz_dataOut_payload_0_4606;
    _zz_dataOut_payload_0_5311 <= _zz_dataOut_payload_0_4607;
    _zz_dataOut_payload_0_5312 <= _zz_dataOut_payload_0_4720;
    _zz_dataOut_payload_0_5313 <= _zz_dataOut_payload_0_4721;
    _zz_dataOut_payload_0_5314 <= _zz_dataOut_payload_0_4722;
    _zz_dataOut_payload_0_5315 <= _zz_dataOut_payload_0_4723;
    _zz_dataOut_payload_0_5316 <= _zz_dataOut_payload_0_4724;
    _zz_dataOut_payload_0_5317 <= _zz_dataOut_payload_0_4725;
    _zz_dataOut_payload_0_5318 <= _zz_dataOut_payload_0_4726;
    _zz_dataOut_payload_0_5319 <= _zz_dataOut_payload_0_4727;
    _zz_dataOut_payload_0_5320 <= _zz_dataOut_payload_0_4728;
    _zz_dataOut_payload_0_5321 <= _zz_dataOut_payload_0_4729;
    _zz_dataOut_payload_0_5322 <= _zz_dataOut_payload_0_4730;
    _zz_dataOut_payload_0_5323 <= _zz_dataOut_payload_0_4731;
    _zz_dataOut_payload_0_5324 <= _zz_dataOut_payload_0_4732;
    _zz_dataOut_payload_0_5325 <= _zz_dataOut_payload_0_4733;
    _zz_dataOut_payload_0_5326 <= _zz_dataOut_payload_0_4734;
    _zz_dataOut_payload_0_5327 <= _zz_dataOut_payload_0_4735;
    _zz_dataOut_payload_0_5328 <= _zz_dataOut_payload_0_4848;
    _zz_dataOut_payload_0_5329 <= _zz_dataOut_payload_0_4849;
    _zz_dataOut_payload_0_5330 <= _zz_dataOut_payload_0_4850;
    _zz_dataOut_payload_0_5331 <= _zz_dataOut_payload_0_4851;
    _zz_dataOut_payload_0_5332 <= _zz_dataOut_payload_0_4852;
    _zz_dataOut_payload_0_5333 <= _zz_dataOut_payload_0_4853;
    _zz_dataOut_payload_0_5334 <= _zz_dataOut_payload_0_4854;
    _zz_dataOut_payload_0_5335 <= _zz_dataOut_payload_0_4855;
    _zz_dataOut_payload_0_5336 <= _zz_dataOut_payload_0_4856;
    _zz_dataOut_payload_0_5337 <= _zz_dataOut_payload_0_4857;
    _zz_dataOut_payload_0_5338 <= _zz_dataOut_payload_0_4858;
    _zz_dataOut_payload_0_5339 <= _zz_dataOut_payload_0_4859;
    _zz_dataOut_payload_0_5340 <= _zz_dataOut_payload_0_4860;
    _zz_dataOut_payload_0_5341 <= _zz_dataOut_payload_0_4861;
    _zz_dataOut_payload_0_5342 <= _zz_dataOut_payload_0_4862;
    _zz_dataOut_payload_0_5343 <= _zz_dataOut_payload_0_4863;
    _zz_dataOut_payload_0_5344 <= _zz_dataOut_payload_0_4976;
    _zz_dataOut_payload_0_5345 <= _zz_dataOut_payload_0_4977;
    _zz_dataOut_payload_0_5346 <= _zz_dataOut_payload_0_4978;
    _zz_dataOut_payload_0_5347 <= _zz_dataOut_payload_0_4979;
    _zz_dataOut_payload_0_5348 <= _zz_dataOut_payload_0_4980;
    _zz_dataOut_payload_0_5349 <= _zz_dataOut_payload_0_4981;
    _zz_dataOut_payload_0_5350 <= _zz_dataOut_payload_0_4982;
    _zz_dataOut_payload_0_5351 <= _zz_dataOut_payload_0_4983;
    _zz_dataOut_payload_0_5352 <= _zz_dataOut_payload_0_4984;
    _zz_dataOut_payload_0_5353 <= _zz_dataOut_payload_0_4985;
    _zz_dataOut_payload_0_5354 <= _zz_dataOut_payload_0_4986;
    _zz_dataOut_payload_0_5355 <= _zz_dataOut_payload_0_4987;
    _zz_dataOut_payload_0_5356 <= _zz_dataOut_payload_0_4988;
    _zz_dataOut_payload_0_5357 <= _zz_dataOut_payload_0_4989;
    _zz_dataOut_payload_0_5358 <= _zz_dataOut_payload_0_4990;
    _zz_dataOut_payload_0_5359 <= _zz_dataOut_payload_0_4991;
    _zz_dataOut_payload_0_5360 <= _zz_dataOut_payload_0_5104;
    _zz_dataOut_payload_0_5361 <= _zz_dataOut_payload_0_5105;
    _zz_dataOut_payload_0_5362 <= _zz_dataOut_payload_0_5106;
    _zz_dataOut_payload_0_5363 <= _zz_dataOut_payload_0_5107;
    _zz_dataOut_payload_0_5364 <= _zz_dataOut_payload_0_5108;
    _zz_dataOut_payload_0_5365 <= _zz_dataOut_payload_0_5109;
    _zz_dataOut_payload_0_5366 <= _zz_dataOut_payload_0_5110;
    _zz_dataOut_payload_0_5367 <= _zz_dataOut_payload_0_5111;
    _zz_dataOut_payload_0_5368 <= _zz_dataOut_payload_0_5112;
    _zz_dataOut_payload_0_5369 <= _zz_dataOut_payload_0_5113;
    _zz_dataOut_payload_0_5370 <= _zz_dataOut_payload_0_5114;
    _zz_dataOut_payload_0_5371 <= _zz_dataOut_payload_0_5115;
    _zz_dataOut_payload_0_5372 <= _zz_dataOut_payload_0_5116;
    _zz_dataOut_payload_0_5373 <= _zz_dataOut_payload_0_5117;
    _zz_dataOut_payload_0_5374 <= _zz_dataOut_payload_0_5118;
    _zz_dataOut_payload_0_5375 <= _zz_dataOut_payload_0_5119;
    _zz_dataOut_payload_0_5468 <= (_zz_dataOut_payload_0_5466 ? _zz_dataOut_payload_0_5461 : _zz_dataOut_payload_0_5464);
    _zz_dataOut_payload_0_5469 <= (_zz_dataOut_payload_0_5466 ? _zz_dataOut_payload_0_5464 : _zz_dataOut_payload_0_5461);
    _zz_dataOut_payload_0_5470 <= (_zz_dataOut_payload_0_5467 ? _zz_dataOut_payload_0_5462 : _zz_dataOut_payload_0_5465);
    _zz_dataOut_payload_0_5471 <= (_zz_dataOut_payload_0_5467 ? _zz_dataOut_payload_0_5465 : _zz_dataOut_payload_0_5462);
    _zz_dataOut_payload_0_5480 <= (_zz_dataOut_payload_0_5478 ? _zz_dataOut_payload_0_5473 : _zz_dataOut_payload_0_5476);
    _zz_dataOut_payload_0_5481 <= (_zz_dataOut_payload_0_5478 ? _zz_dataOut_payload_0_5476 : _zz_dataOut_payload_0_5473);
    _zz_dataOut_payload_0_5482 <= (_zz_dataOut_payload_0_5479 ? _zz_dataOut_payload_0_5474 : _zz_dataOut_payload_0_5477);
    _zz_dataOut_payload_0_5483 <= (_zz_dataOut_payload_0_5479 ? _zz_dataOut_payload_0_5477 : _zz_dataOut_payload_0_5474);
    _zz_dataOut_payload_0_5484 <= _zz_dataOut_payload_0_5468;
    _zz_dataOut_payload_0_5485 <= _zz_dataOut_payload_0_5469;
    _zz_dataOut_payload_0_5486 <= _zz_dataOut_payload_0_5470;
    _zz_dataOut_payload_0_5487 <= _zz_dataOut_payload_0_5471;
    _zz_dataOut_payload_0_5488 <= _zz_dataOut_payload_0_5480;
    _zz_dataOut_payload_0_5489 <= _zz_dataOut_payload_0_5481;
    _zz_dataOut_payload_0_5490 <= _zz_dataOut_payload_0_5482;
    _zz_dataOut_payload_0_5491 <= _zz_dataOut_payload_0_5483;
    _zz_dataOut_payload_0_5512 <= (_zz_dataOut_payload_0_5510 ? _zz_dataOut_payload_0_5505 : _zz_dataOut_payload_0_5508);
    _zz_dataOut_payload_0_5513 <= (_zz_dataOut_payload_0_5510 ? _zz_dataOut_payload_0_5508 : _zz_dataOut_payload_0_5505);
    _zz_dataOut_payload_0_5514 <= (_zz_dataOut_payload_0_5511 ? _zz_dataOut_payload_0_5506 : _zz_dataOut_payload_0_5509);
    _zz_dataOut_payload_0_5515 <= (_zz_dataOut_payload_0_5511 ? _zz_dataOut_payload_0_5509 : _zz_dataOut_payload_0_5506);
    _zz_dataOut_payload_0_5524 <= (_zz_dataOut_payload_0_5522 ? _zz_dataOut_payload_0_5517 : _zz_dataOut_payload_0_5520);
    _zz_dataOut_payload_0_5525 <= (_zz_dataOut_payload_0_5522 ? _zz_dataOut_payload_0_5520 : _zz_dataOut_payload_0_5517);
    _zz_dataOut_payload_0_5526 <= (_zz_dataOut_payload_0_5523 ? _zz_dataOut_payload_0_5518 : _zz_dataOut_payload_0_5521);
    _zz_dataOut_payload_0_5527 <= (_zz_dataOut_payload_0_5523 ? _zz_dataOut_payload_0_5521 : _zz_dataOut_payload_0_5518);
    _zz_dataOut_payload_0_5528 <= _zz_dataOut_payload_0_5512;
    _zz_dataOut_payload_0_5529 <= _zz_dataOut_payload_0_5513;
    _zz_dataOut_payload_0_5530 <= _zz_dataOut_payload_0_5514;
    _zz_dataOut_payload_0_5531 <= _zz_dataOut_payload_0_5515;
    _zz_dataOut_payload_0_5532 <= _zz_dataOut_payload_0_5524;
    _zz_dataOut_payload_0_5533 <= _zz_dataOut_payload_0_5525;
    _zz_dataOut_payload_0_5534 <= _zz_dataOut_payload_0_5526;
    _zz_dataOut_payload_0_5535 <= _zz_dataOut_payload_0_5527;
    _zz_dataOut_payload_0_5536 <= _zz_dataOut_payload_0_5484;
    _zz_dataOut_payload_0_5537 <= _zz_dataOut_payload_0_5485;
    _zz_dataOut_payload_0_5538 <= _zz_dataOut_payload_0_5486;
    _zz_dataOut_payload_0_5539 <= _zz_dataOut_payload_0_5487;
    _zz_dataOut_payload_0_5540 <= _zz_dataOut_payload_0_5488;
    _zz_dataOut_payload_0_5541 <= _zz_dataOut_payload_0_5489;
    _zz_dataOut_payload_0_5542 <= _zz_dataOut_payload_0_5490;
    _zz_dataOut_payload_0_5543 <= _zz_dataOut_payload_0_5491;
    _zz_dataOut_payload_0_5544 <= _zz_dataOut_payload_0_5528;
    _zz_dataOut_payload_0_5545 <= _zz_dataOut_payload_0_5529;
    _zz_dataOut_payload_0_5546 <= _zz_dataOut_payload_0_5530;
    _zz_dataOut_payload_0_5547 <= _zz_dataOut_payload_0_5531;
    _zz_dataOut_payload_0_5548 <= _zz_dataOut_payload_0_5532;
    _zz_dataOut_payload_0_5549 <= _zz_dataOut_payload_0_5533;
    _zz_dataOut_payload_0_5550 <= _zz_dataOut_payload_0_5534;
    _zz_dataOut_payload_0_5551 <= _zz_dataOut_payload_0_5535;
    _zz_dataOut_payload_0_5596 <= (_zz_dataOut_payload_0_5594 ? _zz_dataOut_payload_0_5589 : _zz_dataOut_payload_0_5592);
    _zz_dataOut_payload_0_5597 <= (_zz_dataOut_payload_0_5594 ? _zz_dataOut_payload_0_5592 : _zz_dataOut_payload_0_5589);
    _zz_dataOut_payload_0_5598 <= (_zz_dataOut_payload_0_5595 ? _zz_dataOut_payload_0_5590 : _zz_dataOut_payload_0_5593);
    _zz_dataOut_payload_0_5599 <= (_zz_dataOut_payload_0_5595 ? _zz_dataOut_payload_0_5593 : _zz_dataOut_payload_0_5590);
    _zz_dataOut_payload_0_5608 <= (_zz_dataOut_payload_0_5606 ? _zz_dataOut_payload_0_5601 : _zz_dataOut_payload_0_5604);
    _zz_dataOut_payload_0_5609 <= (_zz_dataOut_payload_0_5606 ? _zz_dataOut_payload_0_5604 : _zz_dataOut_payload_0_5601);
    _zz_dataOut_payload_0_5610 <= (_zz_dataOut_payload_0_5607 ? _zz_dataOut_payload_0_5602 : _zz_dataOut_payload_0_5605);
    _zz_dataOut_payload_0_5611 <= (_zz_dataOut_payload_0_5607 ? _zz_dataOut_payload_0_5605 : _zz_dataOut_payload_0_5602);
    _zz_dataOut_payload_0_5612 <= _zz_dataOut_payload_0_5596;
    _zz_dataOut_payload_0_5613 <= _zz_dataOut_payload_0_5597;
    _zz_dataOut_payload_0_5614 <= _zz_dataOut_payload_0_5598;
    _zz_dataOut_payload_0_5615 <= _zz_dataOut_payload_0_5599;
    _zz_dataOut_payload_0_5616 <= _zz_dataOut_payload_0_5608;
    _zz_dataOut_payload_0_5617 <= _zz_dataOut_payload_0_5609;
    _zz_dataOut_payload_0_5618 <= _zz_dataOut_payload_0_5610;
    _zz_dataOut_payload_0_5619 <= _zz_dataOut_payload_0_5611;
    _zz_dataOut_payload_0_5640 <= (_zz_dataOut_payload_0_5638 ? _zz_dataOut_payload_0_5633 : _zz_dataOut_payload_0_5636);
    _zz_dataOut_payload_0_5641 <= (_zz_dataOut_payload_0_5638 ? _zz_dataOut_payload_0_5636 : _zz_dataOut_payload_0_5633);
    _zz_dataOut_payload_0_5642 <= (_zz_dataOut_payload_0_5639 ? _zz_dataOut_payload_0_5634 : _zz_dataOut_payload_0_5637);
    _zz_dataOut_payload_0_5643 <= (_zz_dataOut_payload_0_5639 ? _zz_dataOut_payload_0_5637 : _zz_dataOut_payload_0_5634);
    _zz_dataOut_payload_0_5652 <= (_zz_dataOut_payload_0_5650 ? _zz_dataOut_payload_0_5645 : _zz_dataOut_payload_0_5648);
    _zz_dataOut_payload_0_5653 <= (_zz_dataOut_payload_0_5650 ? _zz_dataOut_payload_0_5648 : _zz_dataOut_payload_0_5645);
    _zz_dataOut_payload_0_5654 <= (_zz_dataOut_payload_0_5651 ? _zz_dataOut_payload_0_5646 : _zz_dataOut_payload_0_5649);
    _zz_dataOut_payload_0_5655 <= (_zz_dataOut_payload_0_5651 ? _zz_dataOut_payload_0_5649 : _zz_dataOut_payload_0_5646);
    _zz_dataOut_payload_0_5656 <= _zz_dataOut_payload_0_5640;
    _zz_dataOut_payload_0_5657 <= _zz_dataOut_payload_0_5641;
    _zz_dataOut_payload_0_5658 <= _zz_dataOut_payload_0_5642;
    _zz_dataOut_payload_0_5659 <= _zz_dataOut_payload_0_5643;
    _zz_dataOut_payload_0_5660 <= _zz_dataOut_payload_0_5652;
    _zz_dataOut_payload_0_5661 <= _zz_dataOut_payload_0_5653;
    _zz_dataOut_payload_0_5662 <= _zz_dataOut_payload_0_5654;
    _zz_dataOut_payload_0_5663 <= _zz_dataOut_payload_0_5655;
    _zz_dataOut_payload_0_5664 <= _zz_dataOut_payload_0_5612;
    _zz_dataOut_payload_0_5665 <= _zz_dataOut_payload_0_5613;
    _zz_dataOut_payload_0_5666 <= _zz_dataOut_payload_0_5614;
    _zz_dataOut_payload_0_5667 <= _zz_dataOut_payload_0_5615;
    _zz_dataOut_payload_0_5668 <= _zz_dataOut_payload_0_5616;
    _zz_dataOut_payload_0_5669 <= _zz_dataOut_payload_0_5617;
    _zz_dataOut_payload_0_5670 <= _zz_dataOut_payload_0_5618;
    _zz_dataOut_payload_0_5671 <= _zz_dataOut_payload_0_5619;
    _zz_dataOut_payload_0_5672 <= _zz_dataOut_payload_0_5656;
    _zz_dataOut_payload_0_5673 <= _zz_dataOut_payload_0_5657;
    _zz_dataOut_payload_0_5674 <= _zz_dataOut_payload_0_5658;
    _zz_dataOut_payload_0_5675 <= _zz_dataOut_payload_0_5659;
    _zz_dataOut_payload_0_5676 <= _zz_dataOut_payload_0_5660;
    _zz_dataOut_payload_0_5677 <= _zz_dataOut_payload_0_5661;
    _zz_dataOut_payload_0_5678 <= _zz_dataOut_payload_0_5662;
    _zz_dataOut_payload_0_5679 <= _zz_dataOut_payload_0_5663;
    _zz_dataOut_payload_0_5680 <= _zz_dataOut_payload_0_5536;
    _zz_dataOut_payload_0_5681 <= _zz_dataOut_payload_0_5537;
    _zz_dataOut_payload_0_5682 <= _zz_dataOut_payload_0_5538;
    _zz_dataOut_payload_0_5683 <= _zz_dataOut_payload_0_5539;
    _zz_dataOut_payload_0_5684 <= _zz_dataOut_payload_0_5540;
    _zz_dataOut_payload_0_5685 <= _zz_dataOut_payload_0_5541;
    _zz_dataOut_payload_0_5686 <= _zz_dataOut_payload_0_5542;
    _zz_dataOut_payload_0_5687 <= _zz_dataOut_payload_0_5543;
    _zz_dataOut_payload_0_5688 <= _zz_dataOut_payload_0_5544;
    _zz_dataOut_payload_0_5689 <= _zz_dataOut_payload_0_5545;
    _zz_dataOut_payload_0_5690 <= _zz_dataOut_payload_0_5546;
    _zz_dataOut_payload_0_5691 <= _zz_dataOut_payload_0_5547;
    _zz_dataOut_payload_0_5692 <= _zz_dataOut_payload_0_5548;
    _zz_dataOut_payload_0_5693 <= _zz_dataOut_payload_0_5549;
    _zz_dataOut_payload_0_5694 <= _zz_dataOut_payload_0_5550;
    _zz_dataOut_payload_0_5695 <= _zz_dataOut_payload_0_5551;
    _zz_dataOut_payload_0_5696 <= _zz_dataOut_payload_0_5664;
    _zz_dataOut_payload_0_5697 <= _zz_dataOut_payload_0_5665;
    _zz_dataOut_payload_0_5698 <= _zz_dataOut_payload_0_5666;
    _zz_dataOut_payload_0_5699 <= _zz_dataOut_payload_0_5667;
    _zz_dataOut_payload_0_5700 <= _zz_dataOut_payload_0_5668;
    _zz_dataOut_payload_0_5701 <= _zz_dataOut_payload_0_5669;
    _zz_dataOut_payload_0_5702 <= _zz_dataOut_payload_0_5670;
    _zz_dataOut_payload_0_5703 <= _zz_dataOut_payload_0_5671;
    _zz_dataOut_payload_0_5704 <= _zz_dataOut_payload_0_5672;
    _zz_dataOut_payload_0_5705 <= _zz_dataOut_payload_0_5673;
    _zz_dataOut_payload_0_5706 <= _zz_dataOut_payload_0_5674;
    _zz_dataOut_payload_0_5707 <= _zz_dataOut_payload_0_5675;
    _zz_dataOut_payload_0_5708 <= _zz_dataOut_payload_0_5676;
    _zz_dataOut_payload_0_5709 <= _zz_dataOut_payload_0_5677;
    _zz_dataOut_payload_0_5710 <= _zz_dataOut_payload_0_5678;
    _zz_dataOut_payload_0_5711 <= _zz_dataOut_payload_0_5679;
    _zz_dataOut_payload_0_5804 <= (_zz_dataOut_payload_0_5802 ? _zz_dataOut_payload_0_5797 : _zz_dataOut_payload_0_5800);
    _zz_dataOut_payload_0_5805 <= (_zz_dataOut_payload_0_5802 ? _zz_dataOut_payload_0_5800 : _zz_dataOut_payload_0_5797);
    _zz_dataOut_payload_0_5806 <= (_zz_dataOut_payload_0_5803 ? _zz_dataOut_payload_0_5798 : _zz_dataOut_payload_0_5801);
    _zz_dataOut_payload_0_5807 <= (_zz_dataOut_payload_0_5803 ? _zz_dataOut_payload_0_5801 : _zz_dataOut_payload_0_5798);
    _zz_dataOut_payload_0_5816 <= (_zz_dataOut_payload_0_5814 ? _zz_dataOut_payload_0_5809 : _zz_dataOut_payload_0_5812);
    _zz_dataOut_payload_0_5817 <= (_zz_dataOut_payload_0_5814 ? _zz_dataOut_payload_0_5812 : _zz_dataOut_payload_0_5809);
    _zz_dataOut_payload_0_5818 <= (_zz_dataOut_payload_0_5815 ? _zz_dataOut_payload_0_5810 : _zz_dataOut_payload_0_5813);
    _zz_dataOut_payload_0_5819 <= (_zz_dataOut_payload_0_5815 ? _zz_dataOut_payload_0_5813 : _zz_dataOut_payload_0_5810);
    _zz_dataOut_payload_0_5820 <= _zz_dataOut_payload_0_5804;
    _zz_dataOut_payload_0_5821 <= _zz_dataOut_payload_0_5805;
    _zz_dataOut_payload_0_5822 <= _zz_dataOut_payload_0_5806;
    _zz_dataOut_payload_0_5823 <= _zz_dataOut_payload_0_5807;
    _zz_dataOut_payload_0_5824 <= _zz_dataOut_payload_0_5816;
    _zz_dataOut_payload_0_5825 <= _zz_dataOut_payload_0_5817;
    _zz_dataOut_payload_0_5826 <= _zz_dataOut_payload_0_5818;
    _zz_dataOut_payload_0_5827 <= _zz_dataOut_payload_0_5819;
    _zz_dataOut_payload_0_5848 <= (_zz_dataOut_payload_0_5846 ? _zz_dataOut_payload_0_5841 : _zz_dataOut_payload_0_5844);
    _zz_dataOut_payload_0_5849 <= (_zz_dataOut_payload_0_5846 ? _zz_dataOut_payload_0_5844 : _zz_dataOut_payload_0_5841);
    _zz_dataOut_payload_0_5850 <= (_zz_dataOut_payload_0_5847 ? _zz_dataOut_payload_0_5842 : _zz_dataOut_payload_0_5845);
    _zz_dataOut_payload_0_5851 <= (_zz_dataOut_payload_0_5847 ? _zz_dataOut_payload_0_5845 : _zz_dataOut_payload_0_5842);
    _zz_dataOut_payload_0_5860 <= (_zz_dataOut_payload_0_5858 ? _zz_dataOut_payload_0_5853 : _zz_dataOut_payload_0_5856);
    _zz_dataOut_payload_0_5861 <= (_zz_dataOut_payload_0_5858 ? _zz_dataOut_payload_0_5856 : _zz_dataOut_payload_0_5853);
    _zz_dataOut_payload_0_5862 <= (_zz_dataOut_payload_0_5859 ? _zz_dataOut_payload_0_5854 : _zz_dataOut_payload_0_5857);
    _zz_dataOut_payload_0_5863 <= (_zz_dataOut_payload_0_5859 ? _zz_dataOut_payload_0_5857 : _zz_dataOut_payload_0_5854);
    _zz_dataOut_payload_0_5864 <= _zz_dataOut_payload_0_5848;
    _zz_dataOut_payload_0_5865 <= _zz_dataOut_payload_0_5849;
    _zz_dataOut_payload_0_5866 <= _zz_dataOut_payload_0_5850;
    _zz_dataOut_payload_0_5867 <= _zz_dataOut_payload_0_5851;
    _zz_dataOut_payload_0_5868 <= _zz_dataOut_payload_0_5860;
    _zz_dataOut_payload_0_5869 <= _zz_dataOut_payload_0_5861;
    _zz_dataOut_payload_0_5870 <= _zz_dataOut_payload_0_5862;
    _zz_dataOut_payload_0_5871 <= _zz_dataOut_payload_0_5863;
    _zz_dataOut_payload_0_5872 <= _zz_dataOut_payload_0_5820;
    _zz_dataOut_payload_0_5873 <= _zz_dataOut_payload_0_5821;
    _zz_dataOut_payload_0_5874 <= _zz_dataOut_payload_0_5822;
    _zz_dataOut_payload_0_5875 <= _zz_dataOut_payload_0_5823;
    _zz_dataOut_payload_0_5876 <= _zz_dataOut_payload_0_5824;
    _zz_dataOut_payload_0_5877 <= _zz_dataOut_payload_0_5825;
    _zz_dataOut_payload_0_5878 <= _zz_dataOut_payload_0_5826;
    _zz_dataOut_payload_0_5879 <= _zz_dataOut_payload_0_5827;
    _zz_dataOut_payload_0_5880 <= _zz_dataOut_payload_0_5864;
    _zz_dataOut_payload_0_5881 <= _zz_dataOut_payload_0_5865;
    _zz_dataOut_payload_0_5882 <= _zz_dataOut_payload_0_5866;
    _zz_dataOut_payload_0_5883 <= _zz_dataOut_payload_0_5867;
    _zz_dataOut_payload_0_5884 <= _zz_dataOut_payload_0_5868;
    _zz_dataOut_payload_0_5885 <= _zz_dataOut_payload_0_5869;
    _zz_dataOut_payload_0_5886 <= _zz_dataOut_payload_0_5870;
    _zz_dataOut_payload_0_5887 <= _zz_dataOut_payload_0_5871;
    _zz_dataOut_payload_0_5932 <= (_zz_dataOut_payload_0_5930 ? _zz_dataOut_payload_0_5925 : _zz_dataOut_payload_0_5928);
    _zz_dataOut_payload_0_5933 <= (_zz_dataOut_payload_0_5930 ? _zz_dataOut_payload_0_5928 : _zz_dataOut_payload_0_5925);
    _zz_dataOut_payload_0_5934 <= (_zz_dataOut_payload_0_5931 ? _zz_dataOut_payload_0_5926 : _zz_dataOut_payload_0_5929);
    _zz_dataOut_payload_0_5935 <= (_zz_dataOut_payload_0_5931 ? _zz_dataOut_payload_0_5929 : _zz_dataOut_payload_0_5926);
    _zz_dataOut_payload_0_5944 <= (_zz_dataOut_payload_0_5942 ? _zz_dataOut_payload_0_5937 : _zz_dataOut_payload_0_5940);
    _zz_dataOut_payload_0_5945 <= (_zz_dataOut_payload_0_5942 ? _zz_dataOut_payload_0_5940 : _zz_dataOut_payload_0_5937);
    _zz_dataOut_payload_0_5946 <= (_zz_dataOut_payload_0_5943 ? _zz_dataOut_payload_0_5938 : _zz_dataOut_payload_0_5941);
    _zz_dataOut_payload_0_5947 <= (_zz_dataOut_payload_0_5943 ? _zz_dataOut_payload_0_5941 : _zz_dataOut_payload_0_5938);
    _zz_dataOut_payload_0_5948 <= _zz_dataOut_payload_0_5932;
    _zz_dataOut_payload_0_5949 <= _zz_dataOut_payload_0_5933;
    _zz_dataOut_payload_0_5950 <= _zz_dataOut_payload_0_5934;
    _zz_dataOut_payload_0_5951 <= _zz_dataOut_payload_0_5935;
    _zz_dataOut_payload_0_5952 <= _zz_dataOut_payload_0_5944;
    _zz_dataOut_payload_0_5953 <= _zz_dataOut_payload_0_5945;
    _zz_dataOut_payload_0_5954 <= _zz_dataOut_payload_0_5946;
    _zz_dataOut_payload_0_5955 <= _zz_dataOut_payload_0_5947;
    _zz_dataOut_payload_0_5976 <= (_zz_dataOut_payload_0_5974 ? _zz_dataOut_payload_0_5969 : _zz_dataOut_payload_0_5972);
    _zz_dataOut_payload_0_5977 <= (_zz_dataOut_payload_0_5974 ? _zz_dataOut_payload_0_5972 : _zz_dataOut_payload_0_5969);
    _zz_dataOut_payload_0_5978 <= (_zz_dataOut_payload_0_5975 ? _zz_dataOut_payload_0_5970 : _zz_dataOut_payload_0_5973);
    _zz_dataOut_payload_0_5979 <= (_zz_dataOut_payload_0_5975 ? _zz_dataOut_payload_0_5973 : _zz_dataOut_payload_0_5970);
    _zz_dataOut_payload_0_5988 <= (_zz_dataOut_payload_0_5986 ? _zz_dataOut_payload_0_5981 : _zz_dataOut_payload_0_5984);
    _zz_dataOut_payload_0_5989 <= (_zz_dataOut_payload_0_5986 ? _zz_dataOut_payload_0_5984 : _zz_dataOut_payload_0_5981);
    _zz_dataOut_payload_0_5990 <= (_zz_dataOut_payload_0_5987 ? _zz_dataOut_payload_0_5982 : _zz_dataOut_payload_0_5985);
    _zz_dataOut_payload_0_5991 <= (_zz_dataOut_payload_0_5987 ? _zz_dataOut_payload_0_5985 : _zz_dataOut_payload_0_5982);
    _zz_dataOut_payload_0_5992 <= _zz_dataOut_payload_0_5976;
    _zz_dataOut_payload_0_5993 <= _zz_dataOut_payload_0_5977;
    _zz_dataOut_payload_0_5994 <= _zz_dataOut_payload_0_5978;
    _zz_dataOut_payload_0_5995 <= _zz_dataOut_payload_0_5979;
    _zz_dataOut_payload_0_5996 <= _zz_dataOut_payload_0_5988;
    _zz_dataOut_payload_0_5997 <= _zz_dataOut_payload_0_5989;
    _zz_dataOut_payload_0_5998 <= _zz_dataOut_payload_0_5990;
    _zz_dataOut_payload_0_5999 <= _zz_dataOut_payload_0_5991;
    _zz_dataOut_payload_0_6000 <= _zz_dataOut_payload_0_5948;
    _zz_dataOut_payload_0_6001 <= _zz_dataOut_payload_0_5949;
    _zz_dataOut_payload_0_6002 <= _zz_dataOut_payload_0_5950;
    _zz_dataOut_payload_0_6003 <= _zz_dataOut_payload_0_5951;
    _zz_dataOut_payload_0_6004 <= _zz_dataOut_payload_0_5952;
    _zz_dataOut_payload_0_6005 <= _zz_dataOut_payload_0_5953;
    _zz_dataOut_payload_0_6006 <= _zz_dataOut_payload_0_5954;
    _zz_dataOut_payload_0_6007 <= _zz_dataOut_payload_0_5955;
    _zz_dataOut_payload_0_6008 <= _zz_dataOut_payload_0_5992;
    _zz_dataOut_payload_0_6009 <= _zz_dataOut_payload_0_5993;
    _zz_dataOut_payload_0_6010 <= _zz_dataOut_payload_0_5994;
    _zz_dataOut_payload_0_6011 <= _zz_dataOut_payload_0_5995;
    _zz_dataOut_payload_0_6012 <= _zz_dataOut_payload_0_5996;
    _zz_dataOut_payload_0_6013 <= _zz_dataOut_payload_0_5997;
    _zz_dataOut_payload_0_6014 <= _zz_dataOut_payload_0_5998;
    _zz_dataOut_payload_0_6015 <= _zz_dataOut_payload_0_5999;
    _zz_dataOut_payload_0_6016 <= _zz_dataOut_payload_0_5872;
    _zz_dataOut_payload_0_6017 <= _zz_dataOut_payload_0_5873;
    _zz_dataOut_payload_0_6018 <= _zz_dataOut_payload_0_5874;
    _zz_dataOut_payload_0_6019 <= _zz_dataOut_payload_0_5875;
    _zz_dataOut_payload_0_6020 <= _zz_dataOut_payload_0_5876;
    _zz_dataOut_payload_0_6021 <= _zz_dataOut_payload_0_5877;
    _zz_dataOut_payload_0_6022 <= _zz_dataOut_payload_0_5878;
    _zz_dataOut_payload_0_6023 <= _zz_dataOut_payload_0_5879;
    _zz_dataOut_payload_0_6024 <= _zz_dataOut_payload_0_5880;
    _zz_dataOut_payload_0_6025 <= _zz_dataOut_payload_0_5881;
    _zz_dataOut_payload_0_6026 <= _zz_dataOut_payload_0_5882;
    _zz_dataOut_payload_0_6027 <= _zz_dataOut_payload_0_5883;
    _zz_dataOut_payload_0_6028 <= _zz_dataOut_payload_0_5884;
    _zz_dataOut_payload_0_6029 <= _zz_dataOut_payload_0_5885;
    _zz_dataOut_payload_0_6030 <= _zz_dataOut_payload_0_5886;
    _zz_dataOut_payload_0_6031 <= _zz_dataOut_payload_0_5887;
    _zz_dataOut_payload_0_6032 <= _zz_dataOut_payload_0_6000;
    _zz_dataOut_payload_0_6033 <= _zz_dataOut_payload_0_6001;
    _zz_dataOut_payload_0_6034 <= _zz_dataOut_payload_0_6002;
    _zz_dataOut_payload_0_6035 <= _zz_dataOut_payload_0_6003;
    _zz_dataOut_payload_0_6036 <= _zz_dataOut_payload_0_6004;
    _zz_dataOut_payload_0_6037 <= _zz_dataOut_payload_0_6005;
    _zz_dataOut_payload_0_6038 <= _zz_dataOut_payload_0_6006;
    _zz_dataOut_payload_0_6039 <= _zz_dataOut_payload_0_6007;
    _zz_dataOut_payload_0_6040 <= _zz_dataOut_payload_0_6008;
    _zz_dataOut_payload_0_6041 <= _zz_dataOut_payload_0_6009;
    _zz_dataOut_payload_0_6042 <= _zz_dataOut_payload_0_6010;
    _zz_dataOut_payload_0_6043 <= _zz_dataOut_payload_0_6011;
    _zz_dataOut_payload_0_6044 <= _zz_dataOut_payload_0_6012;
    _zz_dataOut_payload_0_6045 <= _zz_dataOut_payload_0_6013;
    _zz_dataOut_payload_0_6046 <= _zz_dataOut_payload_0_6014;
    _zz_dataOut_payload_0_6047 <= _zz_dataOut_payload_0_6015;
    _zz_dataOut_payload_0_6140 <= (_zz_dataOut_payload_0_6138 ? _zz_dataOut_payload_0_6133 : _zz_dataOut_payload_0_6136);
    _zz_dataOut_payload_0_6141 <= (_zz_dataOut_payload_0_6138 ? _zz_dataOut_payload_0_6136 : _zz_dataOut_payload_0_6133);
    _zz_dataOut_payload_0_6142 <= (_zz_dataOut_payload_0_6139 ? _zz_dataOut_payload_0_6134 : _zz_dataOut_payload_0_6137);
    _zz_dataOut_payload_0_6143 <= (_zz_dataOut_payload_0_6139 ? _zz_dataOut_payload_0_6137 : _zz_dataOut_payload_0_6134);
    _zz_dataOut_payload_0_6152 <= (_zz_dataOut_payload_0_6150 ? _zz_dataOut_payload_0_6145 : _zz_dataOut_payload_0_6148);
    _zz_dataOut_payload_0_6153 <= (_zz_dataOut_payload_0_6150 ? _zz_dataOut_payload_0_6148 : _zz_dataOut_payload_0_6145);
    _zz_dataOut_payload_0_6154 <= (_zz_dataOut_payload_0_6151 ? _zz_dataOut_payload_0_6146 : _zz_dataOut_payload_0_6149);
    _zz_dataOut_payload_0_6155 <= (_zz_dataOut_payload_0_6151 ? _zz_dataOut_payload_0_6149 : _zz_dataOut_payload_0_6146);
    _zz_dataOut_payload_0_6156 <= _zz_dataOut_payload_0_6140;
    _zz_dataOut_payload_0_6157 <= _zz_dataOut_payload_0_6141;
    _zz_dataOut_payload_0_6158 <= _zz_dataOut_payload_0_6142;
    _zz_dataOut_payload_0_6159 <= _zz_dataOut_payload_0_6143;
    _zz_dataOut_payload_0_6160 <= _zz_dataOut_payload_0_6152;
    _zz_dataOut_payload_0_6161 <= _zz_dataOut_payload_0_6153;
    _zz_dataOut_payload_0_6162 <= _zz_dataOut_payload_0_6154;
    _zz_dataOut_payload_0_6163 <= _zz_dataOut_payload_0_6155;
    _zz_dataOut_payload_0_6184 <= (_zz_dataOut_payload_0_6182 ? _zz_dataOut_payload_0_6177 : _zz_dataOut_payload_0_6180);
    _zz_dataOut_payload_0_6185 <= (_zz_dataOut_payload_0_6182 ? _zz_dataOut_payload_0_6180 : _zz_dataOut_payload_0_6177);
    _zz_dataOut_payload_0_6186 <= (_zz_dataOut_payload_0_6183 ? _zz_dataOut_payload_0_6178 : _zz_dataOut_payload_0_6181);
    _zz_dataOut_payload_0_6187 <= (_zz_dataOut_payload_0_6183 ? _zz_dataOut_payload_0_6181 : _zz_dataOut_payload_0_6178);
    _zz_dataOut_payload_0_6196 <= (_zz_dataOut_payload_0_6194 ? _zz_dataOut_payload_0_6189 : _zz_dataOut_payload_0_6192);
    _zz_dataOut_payload_0_6197 <= (_zz_dataOut_payload_0_6194 ? _zz_dataOut_payload_0_6192 : _zz_dataOut_payload_0_6189);
    _zz_dataOut_payload_0_6198 <= (_zz_dataOut_payload_0_6195 ? _zz_dataOut_payload_0_6190 : _zz_dataOut_payload_0_6193);
    _zz_dataOut_payload_0_6199 <= (_zz_dataOut_payload_0_6195 ? _zz_dataOut_payload_0_6193 : _zz_dataOut_payload_0_6190);
    _zz_dataOut_payload_0_6200 <= _zz_dataOut_payload_0_6184;
    _zz_dataOut_payload_0_6201 <= _zz_dataOut_payload_0_6185;
    _zz_dataOut_payload_0_6202 <= _zz_dataOut_payload_0_6186;
    _zz_dataOut_payload_0_6203 <= _zz_dataOut_payload_0_6187;
    _zz_dataOut_payload_0_6204 <= _zz_dataOut_payload_0_6196;
    _zz_dataOut_payload_0_6205 <= _zz_dataOut_payload_0_6197;
    _zz_dataOut_payload_0_6206 <= _zz_dataOut_payload_0_6198;
    _zz_dataOut_payload_0_6207 <= _zz_dataOut_payload_0_6199;
    _zz_dataOut_payload_0_6208 <= _zz_dataOut_payload_0_6156;
    _zz_dataOut_payload_0_6209 <= _zz_dataOut_payload_0_6157;
    _zz_dataOut_payload_0_6210 <= _zz_dataOut_payload_0_6158;
    _zz_dataOut_payload_0_6211 <= _zz_dataOut_payload_0_6159;
    _zz_dataOut_payload_0_6212 <= _zz_dataOut_payload_0_6160;
    _zz_dataOut_payload_0_6213 <= _zz_dataOut_payload_0_6161;
    _zz_dataOut_payload_0_6214 <= _zz_dataOut_payload_0_6162;
    _zz_dataOut_payload_0_6215 <= _zz_dataOut_payload_0_6163;
    _zz_dataOut_payload_0_6216 <= _zz_dataOut_payload_0_6200;
    _zz_dataOut_payload_0_6217 <= _zz_dataOut_payload_0_6201;
    _zz_dataOut_payload_0_6218 <= _zz_dataOut_payload_0_6202;
    _zz_dataOut_payload_0_6219 <= _zz_dataOut_payload_0_6203;
    _zz_dataOut_payload_0_6220 <= _zz_dataOut_payload_0_6204;
    _zz_dataOut_payload_0_6221 <= _zz_dataOut_payload_0_6205;
    _zz_dataOut_payload_0_6222 <= _zz_dataOut_payload_0_6206;
    _zz_dataOut_payload_0_6223 <= _zz_dataOut_payload_0_6207;
    _zz_dataOut_payload_0_6268 <= (_zz_dataOut_payload_0_6266 ? _zz_dataOut_payload_0_6261 : _zz_dataOut_payload_0_6264);
    _zz_dataOut_payload_0_6269 <= (_zz_dataOut_payload_0_6266 ? _zz_dataOut_payload_0_6264 : _zz_dataOut_payload_0_6261);
    _zz_dataOut_payload_0_6270 <= (_zz_dataOut_payload_0_6267 ? _zz_dataOut_payload_0_6262 : _zz_dataOut_payload_0_6265);
    _zz_dataOut_payload_0_6271 <= (_zz_dataOut_payload_0_6267 ? _zz_dataOut_payload_0_6265 : _zz_dataOut_payload_0_6262);
    _zz_dataOut_payload_0_6280 <= (_zz_dataOut_payload_0_6278 ? _zz_dataOut_payload_0_6273 : _zz_dataOut_payload_0_6276);
    _zz_dataOut_payload_0_6281 <= (_zz_dataOut_payload_0_6278 ? _zz_dataOut_payload_0_6276 : _zz_dataOut_payload_0_6273);
    _zz_dataOut_payload_0_6282 <= (_zz_dataOut_payload_0_6279 ? _zz_dataOut_payload_0_6274 : _zz_dataOut_payload_0_6277);
    _zz_dataOut_payload_0_6283 <= (_zz_dataOut_payload_0_6279 ? _zz_dataOut_payload_0_6277 : _zz_dataOut_payload_0_6274);
    _zz_dataOut_payload_0_6284 <= _zz_dataOut_payload_0_6268;
    _zz_dataOut_payload_0_6285 <= _zz_dataOut_payload_0_6269;
    _zz_dataOut_payload_0_6286 <= _zz_dataOut_payload_0_6270;
    _zz_dataOut_payload_0_6287 <= _zz_dataOut_payload_0_6271;
    _zz_dataOut_payload_0_6288 <= _zz_dataOut_payload_0_6280;
    _zz_dataOut_payload_0_6289 <= _zz_dataOut_payload_0_6281;
    _zz_dataOut_payload_0_6290 <= _zz_dataOut_payload_0_6282;
    _zz_dataOut_payload_0_6291 <= _zz_dataOut_payload_0_6283;
    _zz_dataOut_payload_0_6312 <= (_zz_dataOut_payload_0_6310 ? _zz_dataOut_payload_0_6305 : _zz_dataOut_payload_0_6308);
    _zz_dataOut_payload_0_6313 <= (_zz_dataOut_payload_0_6310 ? _zz_dataOut_payload_0_6308 : _zz_dataOut_payload_0_6305);
    _zz_dataOut_payload_0_6314 <= (_zz_dataOut_payload_0_6311 ? _zz_dataOut_payload_0_6306 : _zz_dataOut_payload_0_6309);
    _zz_dataOut_payload_0_6315 <= (_zz_dataOut_payload_0_6311 ? _zz_dataOut_payload_0_6309 : _zz_dataOut_payload_0_6306);
    _zz_dataOut_payload_0_6324 <= (_zz_dataOut_payload_0_6322 ? _zz_dataOut_payload_0_6317 : _zz_dataOut_payload_0_6320);
    _zz_dataOut_payload_0_6325 <= (_zz_dataOut_payload_0_6322 ? _zz_dataOut_payload_0_6320 : _zz_dataOut_payload_0_6317);
    _zz_dataOut_payload_0_6326 <= (_zz_dataOut_payload_0_6323 ? _zz_dataOut_payload_0_6318 : _zz_dataOut_payload_0_6321);
    _zz_dataOut_payload_0_6327 <= (_zz_dataOut_payload_0_6323 ? _zz_dataOut_payload_0_6321 : _zz_dataOut_payload_0_6318);
    _zz_dataOut_payload_0_6328 <= _zz_dataOut_payload_0_6312;
    _zz_dataOut_payload_0_6329 <= _zz_dataOut_payload_0_6313;
    _zz_dataOut_payload_0_6330 <= _zz_dataOut_payload_0_6314;
    _zz_dataOut_payload_0_6331 <= _zz_dataOut_payload_0_6315;
    _zz_dataOut_payload_0_6332 <= _zz_dataOut_payload_0_6324;
    _zz_dataOut_payload_0_6333 <= _zz_dataOut_payload_0_6325;
    _zz_dataOut_payload_0_6334 <= _zz_dataOut_payload_0_6326;
    _zz_dataOut_payload_0_6335 <= _zz_dataOut_payload_0_6327;
    _zz_dataOut_payload_0_6336 <= _zz_dataOut_payload_0_6284;
    _zz_dataOut_payload_0_6337 <= _zz_dataOut_payload_0_6285;
    _zz_dataOut_payload_0_6338 <= _zz_dataOut_payload_0_6286;
    _zz_dataOut_payload_0_6339 <= _zz_dataOut_payload_0_6287;
    _zz_dataOut_payload_0_6340 <= _zz_dataOut_payload_0_6288;
    _zz_dataOut_payload_0_6341 <= _zz_dataOut_payload_0_6289;
    _zz_dataOut_payload_0_6342 <= _zz_dataOut_payload_0_6290;
    _zz_dataOut_payload_0_6343 <= _zz_dataOut_payload_0_6291;
    _zz_dataOut_payload_0_6344 <= _zz_dataOut_payload_0_6328;
    _zz_dataOut_payload_0_6345 <= _zz_dataOut_payload_0_6329;
    _zz_dataOut_payload_0_6346 <= _zz_dataOut_payload_0_6330;
    _zz_dataOut_payload_0_6347 <= _zz_dataOut_payload_0_6331;
    _zz_dataOut_payload_0_6348 <= _zz_dataOut_payload_0_6332;
    _zz_dataOut_payload_0_6349 <= _zz_dataOut_payload_0_6333;
    _zz_dataOut_payload_0_6350 <= _zz_dataOut_payload_0_6334;
    _zz_dataOut_payload_0_6351 <= _zz_dataOut_payload_0_6335;
    _zz_dataOut_payload_0_6352 <= _zz_dataOut_payload_0_6208;
    _zz_dataOut_payload_0_6353 <= _zz_dataOut_payload_0_6209;
    _zz_dataOut_payload_0_6354 <= _zz_dataOut_payload_0_6210;
    _zz_dataOut_payload_0_6355 <= _zz_dataOut_payload_0_6211;
    _zz_dataOut_payload_0_6356 <= _zz_dataOut_payload_0_6212;
    _zz_dataOut_payload_0_6357 <= _zz_dataOut_payload_0_6213;
    _zz_dataOut_payload_0_6358 <= _zz_dataOut_payload_0_6214;
    _zz_dataOut_payload_0_6359 <= _zz_dataOut_payload_0_6215;
    _zz_dataOut_payload_0_6360 <= _zz_dataOut_payload_0_6216;
    _zz_dataOut_payload_0_6361 <= _zz_dataOut_payload_0_6217;
    _zz_dataOut_payload_0_6362 <= _zz_dataOut_payload_0_6218;
    _zz_dataOut_payload_0_6363 <= _zz_dataOut_payload_0_6219;
    _zz_dataOut_payload_0_6364 <= _zz_dataOut_payload_0_6220;
    _zz_dataOut_payload_0_6365 <= _zz_dataOut_payload_0_6221;
    _zz_dataOut_payload_0_6366 <= _zz_dataOut_payload_0_6222;
    _zz_dataOut_payload_0_6367 <= _zz_dataOut_payload_0_6223;
    _zz_dataOut_payload_0_6368 <= _zz_dataOut_payload_0_6336;
    _zz_dataOut_payload_0_6369 <= _zz_dataOut_payload_0_6337;
    _zz_dataOut_payload_0_6370 <= _zz_dataOut_payload_0_6338;
    _zz_dataOut_payload_0_6371 <= _zz_dataOut_payload_0_6339;
    _zz_dataOut_payload_0_6372 <= _zz_dataOut_payload_0_6340;
    _zz_dataOut_payload_0_6373 <= _zz_dataOut_payload_0_6341;
    _zz_dataOut_payload_0_6374 <= _zz_dataOut_payload_0_6342;
    _zz_dataOut_payload_0_6375 <= _zz_dataOut_payload_0_6343;
    _zz_dataOut_payload_0_6376 <= _zz_dataOut_payload_0_6344;
    _zz_dataOut_payload_0_6377 <= _zz_dataOut_payload_0_6345;
    _zz_dataOut_payload_0_6378 <= _zz_dataOut_payload_0_6346;
    _zz_dataOut_payload_0_6379 <= _zz_dataOut_payload_0_6347;
    _zz_dataOut_payload_0_6380 <= _zz_dataOut_payload_0_6348;
    _zz_dataOut_payload_0_6381 <= _zz_dataOut_payload_0_6349;
    _zz_dataOut_payload_0_6382 <= _zz_dataOut_payload_0_6350;
    _zz_dataOut_payload_0_6383 <= _zz_dataOut_payload_0_6351;
    _zz_dataOut_payload_0_6476 <= (_zz_dataOut_payload_0_6474 ? _zz_dataOut_payload_0_6469 : _zz_dataOut_payload_0_6472);
    _zz_dataOut_payload_0_6477 <= (_zz_dataOut_payload_0_6474 ? _zz_dataOut_payload_0_6472 : _zz_dataOut_payload_0_6469);
    _zz_dataOut_payload_0_6478 <= (_zz_dataOut_payload_0_6475 ? _zz_dataOut_payload_0_6470 : _zz_dataOut_payload_0_6473);
    _zz_dataOut_payload_0_6479 <= (_zz_dataOut_payload_0_6475 ? _zz_dataOut_payload_0_6473 : _zz_dataOut_payload_0_6470);
    _zz_dataOut_payload_0_6488 <= (_zz_dataOut_payload_0_6486 ? _zz_dataOut_payload_0_6481 : _zz_dataOut_payload_0_6484);
    _zz_dataOut_payload_0_6489 <= (_zz_dataOut_payload_0_6486 ? _zz_dataOut_payload_0_6484 : _zz_dataOut_payload_0_6481);
    _zz_dataOut_payload_0_6490 <= (_zz_dataOut_payload_0_6487 ? _zz_dataOut_payload_0_6482 : _zz_dataOut_payload_0_6485);
    _zz_dataOut_payload_0_6491 <= (_zz_dataOut_payload_0_6487 ? _zz_dataOut_payload_0_6485 : _zz_dataOut_payload_0_6482);
    _zz_dataOut_payload_0_6492 <= _zz_dataOut_payload_0_6476;
    _zz_dataOut_payload_0_6493 <= _zz_dataOut_payload_0_6477;
    _zz_dataOut_payload_0_6494 <= _zz_dataOut_payload_0_6478;
    _zz_dataOut_payload_0_6495 <= _zz_dataOut_payload_0_6479;
    _zz_dataOut_payload_0_6496 <= _zz_dataOut_payload_0_6488;
    _zz_dataOut_payload_0_6497 <= _zz_dataOut_payload_0_6489;
    _zz_dataOut_payload_0_6498 <= _zz_dataOut_payload_0_6490;
    _zz_dataOut_payload_0_6499 <= _zz_dataOut_payload_0_6491;
    _zz_dataOut_payload_0_6520 <= (_zz_dataOut_payload_0_6518 ? _zz_dataOut_payload_0_6513 : _zz_dataOut_payload_0_6516);
    _zz_dataOut_payload_0_6521 <= (_zz_dataOut_payload_0_6518 ? _zz_dataOut_payload_0_6516 : _zz_dataOut_payload_0_6513);
    _zz_dataOut_payload_0_6522 <= (_zz_dataOut_payload_0_6519 ? _zz_dataOut_payload_0_6514 : _zz_dataOut_payload_0_6517);
    _zz_dataOut_payload_0_6523 <= (_zz_dataOut_payload_0_6519 ? _zz_dataOut_payload_0_6517 : _zz_dataOut_payload_0_6514);
    _zz_dataOut_payload_0_6532 <= (_zz_dataOut_payload_0_6530 ? _zz_dataOut_payload_0_6525 : _zz_dataOut_payload_0_6528);
    _zz_dataOut_payload_0_6533 <= (_zz_dataOut_payload_0_6530 ? _zz_dataOut_payload_0_6528 : _zz_dataOut_payload_0_6525);
    _zz_dataOut_payload_0_6534 <= (_zz_dataOut_payload_0_6531 ? _zz_dataOut_payload_0_6526 : _zz_dataOut_payload_0_6529);
    _zz_dataOut_payload_0_6535 <= (_zz_dataOut_payload_0_6531 ? _zz_dataOut_payload_0_6529 : _zz_dataOut_payload_0_6526);
    _zz_dataOut_payload_0_6536 <= _zz_dataOut_payload_0_6520;
    _zz_dataOut_payload_0_6537 <= _zz_dataOut_payload_0_6521;
    _zz_dataOut_payload_0_6538 <= _zz_dataOut_payload_0_6522;
    _zz_dataOut_payload_0_6539 <= _zz_dataOut_payload_0_6523;
    _zz_dataOut_payload_0_6540 <= _zz_dataOut_payload_0_6532;
    _zz_dataOut_payload_0_6541 <= _zz_dataOut_payload_0_6533;
    _zz_dataOut_payload_0_6542 <= _zz_dataOut_payload_0_6534;
    _zz_dataOut_payload_0_6543 <= _zz_dataOut_payload_0_6535;
    _zz_dataOut_payload_0_6544 <= _zz_dataOut_payload_0_6492;
    _zz_dataOut_payload_0_6545 <= _zz_dataOut_payload_0_6493;
    _zz_dataOut_payload_0_6546 <= _zz_dataOut_payload_0_6494;
    _zz_dataOut_payload_0_6547 <= _zz_dataOut_payload_0_6495;
    _zz_dataOut_payload_0_6548 <= _zz_dataOut_payload_0_6496;
    _zz_dataOut_payload_0_6549 <= _zz_dataOut_payload_0_6497;
    _zz_dataOut_payload_0_6550 <= _zz_dataOut_payload_0_6498;
    _zz_dataOut_payload_0_6551 <= _zz_dataOut_payload_0_6499;
    _zz_dataOut_payload_0_6552 <= _zz_dataOut_payload_0_6536;
    _zz_dataOut_payload_0_6553 <= _zz_dataOut_payload_0_6537;
    _zz_dataOut_payload_0_6554 <= _zz_dataOut_payload_0_6538;
    _zz_dataOut_payload_0_6555 <= _zz_dataOut_payload_0_6539;
    _zz_dataOut_payload_0_6556 <= _zz_dataOut_payload_0_6540;
    _zz_dataOut_payload_0_6557 <= _zz_dataOut_payload_0_6541;
    _zz_dataOut_payload_0_6558 <= _zz_dataOut_payload_0_6542;
    _zz_dataOut_payload_0_6559 <= _zz_dataOut_payload_0_6543;
    _zz_dataOut_payload_0_6604 <= (_zz_dataOut_payload_0_6602 ? _zz_dataOut_payload_0_6597 : _zz_dataOut_payload_0_6600);
    _zz_dataOut_payload_0_6605 <= (_zz_dataOut_payload_0_6602 ? _zz_dataOut_payload_0_6600 : _zz_dataOut_payload_0_6597);
    _zz_dataOut_payload_0_6606 <= (_zz_dataOut_payload_0_6603 ? _zz_dataOut_payload_0_6598 : _zz_dataOut_payload_0_6601);
    _zz_dataOut_payload_0_6607 <= (_zz_dataOut_payload_0_6603 ? _zz_dataOut_payload_0_6601 : _zz_dataOut_payload_0_6598);
    _zz_dataOut_payload_0_6616 <= (_zz_dataOut_payload_0_6614 ? _zz_dataOut_payload_0_6609 : _zz_dataOut_payload_0_6612);
    _zz_dataOut_payload_0_6617 <= (_zz_dataOut_payload_0_6614 ? _zz_dataOut_payload_0_6612 : _zz_dataOut_payload_0_6609);
    _zz_dataOut_payload_0_6618 <= (_zz_dataOut_payload_0_6615 ? _zz_dataOut_payload_0_6610 : _zz_dataOut_payload_0_6613);
    _zz_dataOut_payload_0_6619 <= (_zz_dataOut_payload_0_6615 ? _zz_dataOut_payload_0_6613 : _zz_dataOut_payload_0_6610);
    _zz_dataOut_payload_0_6620 <= _zz_dataOut_payload_0_6604;
    _zz_dataOut_payload_0_6621 <= _zz_dataOut_payload_0_6605;
    _zz_dataOut_payload_0_6622 <= _zz_dataOut_payload_0_6606;
    _zz_dataOut_payload_0_6623 <= _zz_dataOut_payload_0_6607;
    _zz_dataOut_payload_0_6624 <= _zz_dataOut_payload_0_6616;
    _zz_dataOut_payload_0_6625 <= _zz_dataOut_payload_0_6617;
    _zz_dataOut_payload_0_6626 <= _zz_dataOut_payload_0_6618;
    _zz_dataOut_payload_0_6627 <= _zz_dataOut_payload_0_6619;
    _zz_dataOut_payload_0_6648 <= (_zz_dataOut_payload_0_6646 ? _zz_dataOut_payload_0_6641 : _zz_dataOut_payload_0_6644);
    _zz_dataOut_payload_0_6649 <= (_zz_dataOut_payload_0_6646 ? _zz_dataOut_payload_0_6644 : _zz_dataOut_payload_0_6641);
    _zz_dataOut_payload_0_6650 <= (_zz_dataOut_payload_0_6647 ? _zz_dataOut_payload_0_6642 : _zz_dataOut_payload_0_6645);
    _zz_dataOut_payload_0_6651 <= (_zz_dataOut_payload_0_6647 ? _zz_dataOut_payload_0_6645 : _zz_dataOut_payload_0_6642);
    _zz_dataOut_payload_0_6660 <= (_zz_dataOut_payload_0_6658 ? _zz_dataOut_payload_0_6653 : _zz_dataOut_payload_0_6656);
    _zz_dataOut_payload_0_6661 <= (_zz_dataOut_payload_0_6658 ? _zz_dataOut_payload_0_6656 : _zz_dataOut_payload_0_6653);
    _zz_dataOut_payload_0_6662 <= (_zz_dataOut_payload_0_6659 ? _zz_dataOut_payload_0_6654 : _zz_dataOut_payload_0_6657);
    _zz_dataOut_payload_0_6663 <= (_zz_dataOut_payload_0_6659 ? _zz_dataOut_payload_0_6657 : _zz_dataOut_payload_0_6654);
    _zz_dataOut_payload_0_6664 <= _zz_dataOut_payload_0_6648;
    _zz_dataOut_payload_0_6665 <= _zz_dataOut_payload_0_6649;
    _zz_dataOut_payload_0_6666 <= _zz_dataOut_payload_0_6650;
    _zz_dataOut_payload_0_6667 <= _zz_dataOut_payload_0_6651;
    _zz_dataOut_payload_0_6668 <= _zz_dataOut_payload_0_6660;
    _zz_dataOut_payload_0_6669 <= _zz_dataOut_payload_0_6661;
    _zz_dataOut_payload_0_6670 <= _zz_dataOut_payload_0_6662;
    _zz_dataOut_payload_0_6671 <= _zz_dataOut_payload_0_6663;
    _zz_dataOut_payload_0_6672 <= _zz_dataOut_payload_0_6620;
    _zz_dataOut_payload_0_6673 <= _zz_dataOut_payload_0_6621;
    _zz_dataOut_payload_0_6674 <= _zz_dataOut_payload_0_6622;
    _zz_dataOut_payload_0_6675 <= _zz_dataOut_payload_0_6623;
    _zz_dataOut_payload_0_6676 <= _zz_dataOut_payload_0_6624;
    _zz_dataOut_payload_0_6677 <= _zz_dataOut_payload_0_6625;
    _zz_dataOut_payload_0_6678 <= _zz_dataOut_payload_0_6626;
    _zz_dataOut_payload_0_6679 <= _zz_dataOut_payload_0_6627;
    _zz_dataOut_payload_0_6680 <= _zz_dataOut_payload_0_6664;
    _zz_dataOut_payload_0_6681 <= _zz_dataOut_payload_0_6665;
    _zz_dataOut_payload_0_6682 <= _zz_dataOut_payload_0_6666;
    _zz_dataOut_payload_0_6683 <= _zz_dataOut_payload_0_6667;
    _zz_dataOut_payload_0_6684 <= _zz_dataOut_payload_0_6668;
    _zz_dataOut_payload_0_6685 <= _zz_dataOut_payload_0_6669;
    _zz_dataOut_payload_0_6686 <= _zz_dataOut_payload_0_6670;
    _zz_dataOut_payload_0_6687 <= _zz_dataOut_payload_0_6671;
    _zz_dataOut_payload_0_6688 <= _zz_dataOut_payload_0_6544;
    _zz_dataOut_payload_0_6689 <= _zz_dataOut_payload_0_6545;
    _zz_dataOut_payload_0_6690 <= _zz_dataOut_payload_0_6546;
    _zz_dataOut_payload_0_6691 <= _zz_dataOut_payload_0_6547;
    _zz_dataOut_payload_0_6692 <= _zz_dataOut_payload_0_6548;
    _zz_dataOut_payload_0_6693 <= _zz_dataOut_payload_0_6549;
    _zz_dataOut_payload_0_6694 <= _zz_dataOut_payload_0_6550;
    _zz_dataOut_payload_0_6695 <= _zz_dataOut_payload_0_6551;
    _zz_dataOut_payload_0_6696 <= _zz_dataOut_payload_0_6552;
    _zz_dataOut_payload_0_6697 <= _zz_dataOut_payload_0_6553;
    _zz_dataOut_payload_0_6698 <= _zz_dataOut_payload_0_6554;
    _zz_dataOut_payload_0_6699 <= _zz_dataOut_payload_0_6555;
    _zz_dataOut_payload_0_6700 <= _zz_dataOut_payload_0_6556;
    _zz_dataOut_payload_0_6701 <= _zz_dataOut_payload_0_6557;
    _zz_dataOut_payload_0_6702 <= _zz_dataOut_payload_0_6558;
    _zz_dataOut_payload_0_6703 <= _zz_dataOut_payload_0_6559;
    _zz_dataOut_payload_0_6704 <= _zz_dataOut_payload_0_6672;
    _zz_dataOut_payload_0_6705 <= _zz_dataOut_payload_0_6673;
    _zz_dataOut_payload_0_6706 <= _zz_dataOut_payload_0_6674;
    _zz_dataOut_payload_0_6707 <= _zz_dataOut_payload_0_6675;
    _zz_dataOut_payload_0_6708 <= _zz_dataOut_payload_0_6676;
    _zz_dataOut_payload_0_6709 <= _zz_dataOut_payload_0_6677;
    _zz_dataOut_payload_0_6710 <= _zz_dataOut_payload_0_6678;
    _zz_dataOut_payload_0_6711 <= _zz_dataOut_payload_0_6679;
    _zz_dataOut_payload_0_6712 <= _zz_dataOut_payload_0_6680;
    _zz_dataOut_payload_0_6713 <= _zz_dataOut_payload_0_6681;
    _zz_dataOut_payload_0_6714 <= _zz_dataOut_payload_0_6682;
    _zz_dataOut_payload_0_6715 <= _zz_dataOut_payload_0_6683;
    _zz_dataOut_payload_0_6716 <= _zz_dataOut_payload_0_6684;
    _zz_dataOut_payload_0_6717 <= _zz_dataOut_payload_0_6685;
    _zz_dataOut_payload_0_6718 <= _zz_dataOut_payload_0_6686;
    _zz_dataOut_payload_0_6719 <= _zz_dataOut_payload_0_6687;
    _zz_dataOut_payload_0_6812 <= (_zz_dataOut_payload_0_6810 ? _zz_dataOut_payload_0_6805 : _zz_dataOut_payload_0_6808);
    _zz_dataOut_payload_0_6813 <= (_zz_dataOut_payload_0_6810 ? _zz_dataOut_payload_0_6808 : _zz_dataOut_payload_0_6805);
    _zz_dataOut_payload_0_6814 <= (_zz_dataOut_payload_0_6811 ? _zz_dataOut_payload_0_6806 : _zz_dataOut_payload_0_6809);
    _zz_dataOut_payload_0_6815 <= (_zz_dataOut_payload_0_6811 ? _zz_dataOut_payload_0_6809 : _zz_dataOut_payload_0_6806);
    _zz_dataOut_payload_0_6824 <= (_zz_dataOut_payload_0_6822 ? _zz_dataOut_payload_0_6817 : _zz_dataOut_payload_0_6820);
    _zz_dataOut_payload_0_6825 <= (_zz_dataOut_payload_0_6822 ? _zz_dataOut_payload_0_6820 : _zz_dataOut_payload_0_6817);
    _zz_dataOut_payload_0_6826 <= (_zz_dataOut_payload_0_6823 ? _zz_dataOut_payload_0_6818 : _zz_dataOut_payload_0_6821);
    _zz_dataOut_payload_0_6827 <= (_zz_dataOut_payload_0_6823 ? _zz_dataOut_payload_0_6821 : _zz_dataOut_payload_0_6818);
    _zz_dataOut_payload_0_6828 <= _zz_dataOut_payload_0_6812;
    _zz_dataOut_payload_0_6829 <= _zz_dataOut_payload_0_6813;
    _zz_dataOut_payload_0_6830 <= _zz_dataOut_payload_0_6814;
    _zz_dataOut_payload_0_6831 <= _zz_dataOut_payload_0_6815;
    _zz_dataOut_payload_0_6832 <= _zz_dataOut_payload_0_6824;
    _zz_dataOut_payload_0_6833 <= _zz_dataOut_payload_0_6825;
    _zz_dataOut_payload_0_6834 <= _zz_dataOut_payload_0_6826;
    _zz_dataOut_payload_0_6835 <= _zz_dataOut_payload_0_6827;
    _zz_dataOut_payload_0_6856 <= (_zz_dataOut_payload_0_6854 ? _zz_dataOut_payload_0_6849 : _zz_dataOut_payload_0_6852);
    _zz_dataOut_payload_0_6857 <= (_zz_dataOut_payload_0_6854 ? _zz_dataOut_payload_0_6852 : _zz_dataOut_payload_0_6849);
    _zz_dataOut_payload_0_6858 <= (_zz_dataOut_payload_0_6855 ? _zz_dataOut_payload_0_6850 : _zz_dataOut_payload_0_6853);
    _zz_dataOut_payload_0_6859 <= (_zz_dataOut_payload_0_6855 ? _zz_dataOut_payload_0_6853 : _zz_dataOut_payload_0_6850);
    _zz_dataOut_payload_0_6868 <= (_zz_dataOut_payload_0_6866 ? _zz_dataOut_payload_0_6861 : _zz_dataOut_payload_0_6864);
    _zz_dataOut_payload_0_6869 <= (_zz_dataOut_payload_0_6866 ? _zz_dataOut_payload_0_6864 : _zz_dataOut_payload_0_6861);
    _zz_dataOut_payload_0_6870 <= (_zz_dataOut_payload_0_6867 ? _zz_dataOut_payload_0_6862 : _zz_dataOut_payload_0_6865);
    _zz_dataOut_payload_0_6871 <= (_zz_dataOut_payload_0_6867 ? _zz_dataOut_payload_0_6865 : _zz_dataOut_payload_0_6862);
    _zz_dataOut_payload_0_6872 <= _zz_dataOut_payload_0_6856;
    _zz_dataOut_payload_0_6873 <= _zz_dataOut_payload_0_6857;
    _zz_dataOut_payload_0_6874 <= _zz_dataOut_payload_0_6858;
    _zz_dataOut_payload_0_6875 <= _zz_dataOut_payload_0_6859;
    _zz_dataOut_payload_0_6876 <= _zz_dataOut_payload_0_6868;
    _zz_dataOut_payload_0_6877 <= _zz_dataOut_payload_0_6869;
    _zz_dataOut_payload_0_6878 <= _zz_dataOut_payload_0_6870;
    _zz_dataOut_payload_0_6879 <= _zz_dataOut_payload_0_6871;
    _zz_dataOut_payload_0_6880 <= _zz_dataOut_payload_0_6828;
    _zz_dataOut_payload_0_6881 <= _zz_dataOut_payload_0_6829;
    _zz_dataOut_payload_0_6882 <= _zz_dataOut_payload_0_6830;
    _zz_dataOut_payload_0_6883 <= _zz_dataOut_payload_0_6831;
    _zz_dataOut_payload_0_6884 <= _zz_dataOut_payload_0_6832;
    _zz_dataOut_payload_0_6885 <= _zz_dataOut_payload_0_6833;
    _zz_dataOut_payload_0_6886 <= _zz_dataOut_payload_0_6834;
    _zz_dataOut_payload_0_6887 <= _zz_dataOut_payload_0_6835;
    _zz_dataOut_payload_0_6888 <= _zz_dataOut_payload_0_6872;
    _zz_dataOut_payload_0_6889 <= _zz_dataOut_payload_0_6873;
    _zz_dataOut_payload_0_6890 <= _zz_dataOut_payload_0_6874;
    _zz_dataOut_payload_0_6891 <= _zz_dataOut_payload_0_6875;
    _zz_dataOut_payload_0_6892 <= _zz_dataOut_payload_0_6876;
    _zz_dataOut_payload_0_6893 <= _zz_dataOut_payload_0_6877;
    _zz_dataOut_payload_0_6894 <= _zz_dataOut_payload_0_6878;
    _zz_dataOut_payload_0_6895 <= _zz_dataOut_payload_0_6879;
    _zz_dataOut_payload_0_6940 <= (_zz_dataOut_payload_0_6938 ? _zz_dataOut_payload_0_6933 : _zz_dataOut_payload_0_6936);
    _zz_dataOut_payload_0_6941 <= (_zz_dataOut_payload_0_6938 ? _zz_dataOut_payload_0_6936 : _zz_dataOut_payload_0_6933);
    _zz_dataOut_payload_0_6942 <= (_zz_dataOut_payload_0_6939 ? _zz_dataOut_payload_0_6934 : _zz_dataOut_payload_0_6937);
    _zz_dataOut_payload_0_6943 <= (_zz_dataOut_payload_0_6939 ? _zz_dataOut_payload_0_6937 : _zz_dataOut_payload_0_6934);
    _zz_dataOut_payload_0_6952 <= (_zz_dataOut_payload_0_6950 ? _zz_dataOut_payload_0_6945 : _zz_dataOut_payload_0_6948);
    _zz_dataOut_payload_0_6953 <= (_zz_dataOut_payload_0_6950 ? _zz_dataOut_payload_0_6948 : _zz_dataOut_payload_0_6945);
    _zz_dataOut_payload_0_6954 <= (_zz_dataOut_payload_0_6951 ? _zz_dataOut_payload_0_6946 : _zz_dataOut_payload_0_6949);
    _zz_dataOut_payload_0_6955 <= (_zz_dataOut_payload_0_6951 ? _zz_dataOut_payload_0_6949 : _zz_dataOut_payload_0_6946);
    _zz_dataOut_payload_0_6956 <= _zz_dataOut_payload_0_6940;
    _zz_dataOut_payload_0_6957 <= _zz_dataOut_payload_0_6941;
    _zz_dataOut_payload_0_6958 <= _zz_dataOut_payload_0_6942;
    _zz_dataOut_payload_0_6959 <= _zz_dataOut_payload_0_6943;
    _zz_dataOut_payload_0_6960 <= _zz_dataOut_payload_0_6952;
    _zz_dataOut_payload_0_6961 <= _zz_dataOut_payload_0_6953;
    _zz_dataOut_payload_0_6962 <= _zz_dataOut_payload_0_6954;
    _zz_dataOut_payload_0_6963 <= _zz_dataOut_payload_0_6955;
    _zz_dataOut_payload_0_6984 <= (_zz_dataOut_payload_0_6982 ? _zz_dataOut_payload_0_6977 : _zz_dataOut_payload_0_6980);
    _zz_dataOut_payload_0_6985 <= (_zz_dataOut_payload_0_6982 ? _zz_dataOut_payload_0_6980 : _zz_dataOut_payload_0_6977);
    _zz_dataOut_payload_0_6986 <= (_zz_dataOut_payload_0_6983 ? _zz_dataOut_payload_0_6978 : _zz_dataOut_payload_0_6981);
    _zz_dataOut_payload_0_6987 <= (_zz_dataOut_payload_0_6983 ? _zz_dataOut_payload_0_6981 : _zz_dataOut_payload_0_6978);
    _zz_dataOut_payload_0_6996 <= (_zz_dataOut_payload_0_6994 ? _zz_dataOut_payload_0_6989 : _zz_dataOut_payload_0_6992);
    _zz_dataOut_payload_0_6997 <= (_zz_dataOut_payload_0_6994 ? _zz_dataOut_payload_0_6992 : _zz_dataOut_payload_0_6989);
    _zz_dataOut_payload_0_6998 <= (_zz_dataOut_payload_0_6995 ? _zz_dataOut_payload_0_6990 : _zz_dataOut_payload_0_6993);
    _zz_dataOut_payload_0_6999 <= (_zz_dataOut_payload_0_6995 ? _zz_dataOut_payload_0_6993 : _zz_dataOut_payload_0_6990);
    _zz_dataOut_payload_0_7000 <= _zz_dataOut_payload_0_6984;
    _zz_dataOut_payload_0_7001 <= _zz_dataOut_payload_0_6985;
    _zz_dataOut_payload_0_7002 <= _zz_dataOut_payload_0_6986;
    _zz_dataOut_payload_0_7003 <= _zz_dataOut_payload_0_6987;
    _zz_dataOut_payload_0_7004 <= _zz_dataOut_payload_0_6996;
    _zz_dataOut_payload_0_7005 <= _zz_dataOut_payload_0_6997;
    _zz_dataOut_payload_0_7006 <= _zz_dataOut_payload_0_6998;
    _zz_dataOut_payload_0_7007 <= _zz_dataOut_payload_0_6999;
    _zz_dataOut_payload_0_7008 <= _zz_dataOut_payload_0_6956;
    _zz_dataOut_payload_0_7009 <= _zz_dataOut_payload_0_6957;
    _zz_dataOut_payload_0_7010 <= _zz_dataOut_payload_0_6958;
    _zz_dataOut_payload_0_7011 <= _zz_dataOut_payload_0_6959;
    _zz_dataOut_payload_0_7012 <= _zz_dataOut_payload_0_6960;
    _zz_dataOut_payload_0_7013 <= _zz_dataOut_payload_0_6961;
    _zz_dataOut_payload_0_7014 <= _zz_dataOut_payload_0_6962;
    _zz_dataOut_payload_0_7015 <= _zz_dataOut_payload_0_6963;
    _zz_dataOut_payload_0_7016 <= _zz_dataOut_payload_0_7000;
    _zz_dataOut_payload_0_7017 <= _zz_dataOut_payload_0_7001;
    _zz_dataOut_payload_0_7018 <= _zz_dataOut_payload_0_7002;
    _zz_dataOut_payload_0_7019 <= _zz_dataOut_payload_0_7003;
    _zz_dataOut_payload_0_7020 <= _zz_dataOut_payload_0_7004;
    _zz_dataOut_payload_0_7021 <= _zz_dataOut_payload_0_7005;
    _zz_dataOut_payload_0_7022 <= _zz_dataOut_payload_0_7006;
    _zz_dataOut_payload_0_7023 <= _zz_dataOut_payload_0_7007;
    _zz_dataOut_payload_0_7024 <= _zz_dataOut_payload_0_6880;
    _zz_dataOut_payload_0_7025 <= _zz_dataOut_payload_0_6881;
    _zz_dataOut_payload_0_7026 <= _zz_dataOut_payload_0_6882;
    _zz_dataOut_payload_0_7027 <= _zz_dataOut_payload_0_6883;
    _zz_dataOut_payload_0_7028 <= _zz_dataOut_payload_0_6884;
    _zz_dataOut_payload_0_7029 <= _zz_dataOut_payload_0_6885;
    _zz_dataOut_payload_0_7030 <= _zz_dataOut_payload_0_6886;
    _zz_dataOut_payload_0_7031 <= _zz_dataOut_payload_0_6887;
    _zz_dataOut_payload_0_7032 <= _zz_dataOut_payload_0_6888;
    _zz_dataOut_payload_0_7033 <= _zz_dataOut_payload_0_6889;
    _zz_dataOut_payload_0_7034 <= _zz_dataOut_payload_0_6890;
    _zz_dataOut_payload_0_7035 <= _zz_dataOut_payload_0_6891;
    _zz_dataOut_payload_0_7036 <= _zz_dataOut_payload_0_6892;
    _zz_dataOut_payload_0_7037 <= _zz_dataOut_payload_0_6893;
    _zz_dataOut_payload_0_7038 <= _zz_dataOut_payload_0_6894;
    _zz_dataOut_payload_0_7039 <= _zz_dataOut_payload_0_6895;
    _zz_dataOut_payload_0_7040 <= _zz_dataOut_payload_0_7008;
    _zz_dataOut_payload_0_7041 <= _zz_dataOut_payload_0_7009;
    _zz_dataOut_payload_0_7042 <= _zz_dataOut_payload_0_7010;
    _zz_dataOut_payload_0_7043 <= _zz_dataOut_payload_0_7011;
    _zz_dataOut_payload_0_7044 <= _zz_dataOut_payload_0_7012;
    _zz_dataOut_payload_0_7045 <= _zz_dataOut_payload_0_7013;
    _zz_dataOut_payload_0_7046 <= _zz_dataOut_payload_0_7014;
    _zz_dataOut_payload_0_7047 <= _zz_dataOut_payload_0_7015;
    _zz_dataOut_payload_0_7048 <= _zz_dataOut_payload_0_7016;
    _zz_dataOut_payload_0_7049 <= _zz_dataOut_payload_0_7017;
    _zz_dataOut_payload_0_7050 <= _zz_dataOut_payload_0_7018;
    _zz_dataOut_payload_0_7051 <= _zz_dataOut_payload_0_7019;
    _zz_dataOut_payload_0_7052 <= _zz_dataOut_payload_0_7020;
    _zz_dataOut_payload_0_7053 <= _zz_dataOut_payload_0_7021;
    _zz_dataOut_payload_0_7054 <= _zz_dataOut_payload_0_7022;
    _zz_dataOut_payload_0_7055 <= _zz_dataOut_payload_0_7023;
    _zz_dataOut_payload_0_7148 <= (_zz_dataOut_payload_0_7146 ? _zz_dataOut_payload_0_7141 : _zz_dataOut_payload_0_7144);
    _zz_dataOut_payload_0_7149 <= (_zz_dataOut_payload_0_7146 ? _zz_dataOut_payload_0_7144 : _zz_dataOut_payload_0_7141);
    _zz_dataOut_payload_0_7150 <= (_zz_dataOut_payload_0_7147 ? _zz_dataOut_payload_0_7142 : _zz_dataOut_payload_0_7145);
    _zz_dataOut_payload_0_7151 <= (_zz_dataOut_payload_0_7147 ? _zz_dataOut_payload_0_7145 : _zz_dataOut_payload_0_7142);
    _zz_dataOut_payload_0_7160 <= (_zz_dataOut_payload_0_7158 ? _zz_dataOut_payload_0_7153 : _zz_dataOut_payload_0_7156);
    _zz_dataOut_payload_0_7161 <= (_zz_dataOut_payload_0_7158 ? _zz_dataOut_payload_0_7156 : _zz_dataOut_payload_0_7153);
    _zz_dataOut_payload_0_7162 <= (_zz_dataOut_payload_0_7159 ? _zz_dataOut_payload_0_7154 : _zz_dataOut_payload_0_7157);
    _zz_dataOut_payload_0_7163 <= (_zz_dataOut_payload_0_7159 ? _zz_dataOut_payload_0_7157 : _zz_dataOut_payload_0_7154);
    _zz_dataOut_payload_0_7164 <= _zz_dataOut_payload_0_7148;
    _zz_dataOut_payload_0_7165 <= _zz_dataOut_payload_0_7149;
    _zz_dataOut_payload_0_7166 <= _zz_dataOut_payload_0_7150;
    _zz_dataOut_payload_0_7167 <= _zz_dataOut_payload_0_7151;
    _zz_dataOut_payload_0_7168 <= _zz_dataOut_payload_0_7160;
    _zz_dataOut_payload_0_7169 <= _zz_dataOut_payload_0_7161;
    _zz_dataOut_payload_0_7170 <= _zz_dataOut_payload_0_7162;
    _zz_dataOut_payload_0_7171 <= _zz_dataOut_payload_0_7163;
    _zz_dataOut_payload_0_7192 <= (_zz_dataOut_payload_0_7190 ? _zz_dataOut_payload_0_7185 : _zz_dataOut_payload_0_7188);
    _zz_dataOut_payload_0_7193 <= (_zz_dataOut_payload_0_7190 ? _zz_dataOut_payload_0_7188 : _zz_dataOut_payload_0_7185);
    _zz_dataOut_payload_0_7194 <= (_zz_dataOut_payload_0_7191 ? _zz_dataOut_payload_0_7186 : _zz_dataOut_payload_0_7189);
    _zz_dataOut_payload_0_7195 <= (_zz_dataOut_payload_0_7191 ? _zz_dataOut_payload_0_7189 : _zz_dataOut_payload_0_7186);
    _zz_dataOut_payload_0_7204 <= (_zz_dataOut_payload_0_7202 ? _zz_dataOut_payload_0_7197 : _zz_dataOut_payload_0_7200);
    _zz_dataOut_payload_0_7205 <= (_zz_dataOut_payload_0_7202 ? _zz_dataOut_payload_0_7200 : _zz_dataOut_payload_0_7197);
    _zz_dataOut_payload_0_7206 <= (_zz_dataOut_payload_0_7203 ? _zz_dataOut_payload_0_7198 : _zz_dataOut_payload_0_7201);
    _zz_dataOut_payload_0_7207 <= (_zz_dataOut_payload_0_7203 ? _zz_dataOut_payload_0_7201 : _zz_dataOut_payload_0_7198);
    _zz_dataOut_payload_0_7208 <= _zz_dataOut_payload_0_7192;
    _zz_dataOut_payload_0_7209 <= _zz_dataOut_payload_0_7193;
    _zz_dataOut_payload_0_7210 <= _zz_dataOut_payload_0_7194;
    _zz_dataOut_payload_0_7211 <= _zz_dataOut_payload_0_7195;
    _zz_dataOut_payload_0_7212 <= _zz_dataOut_payload_0_7204;
    _zz_dataOut_payload_0_7213 <= _zz_dataOut_payload_0_7205;
    _zz_dataOut_payload_0_7214 <= _zz_dataOut_payload_0_7206;
    _zz_dataOut_payload_0_7215 <= _zz_dataOut_payload_0_7207;
    _zz_dataOut_payload_0_7216 <= _zz_dataOut_payload_0_7164;
    _zz_dataOut_payload_0_7217 <= _zz_dataOut_payload_0_7165;
    _zz_dataOut_payload_0_7218 <= _zz_dataOut_payload_0_7166;
    _zz_dataOut_payload_0_7219 <= _zz_dataOut_payload_0_7167;
    _zz_dataOut_payload_0_7220 <= _zz_dataOut_payload_0_7168;
    _zz_dataOut_payload_0_7221 <= _zz_dataOut_payload_0_7169;
    _zz_dataOut_payload_0_7222 <= _zz_dataOut_payload_0_7170;
    _zz_dataOut_payload_0_7223 <= _zz_dataOut_payload_0_7171;
    _zz_dataOut_payload_0_7224 <= _zz_dataOut_payload_0_7208;
    _zz_dataOut_payload_0_7225 <= _zz_dataOut_payload_0_7209;
    _zz_dataOut_payload_0_7226 <= _zz_dataOut_payload_0_7210;
    _zz_dataOut_payload_0_7227 <= _zz_dataOut_payload_0_7211;
    _zz_dataOut_payload_0_7228 <= _zz_dataOut_payload_0_7212;
    _zz_dataOut_payload_0_7229 <= _zz_dataOut_payload_0_7213;
    _zz_dataOut_payload_0_7230 <= _zz_dataOut_payload_0_7214;
    _zz_dataOut_payload_0_7231 <= _zz_dataOut_payload_0_7215;
    _zz_dataOut_payload_0_7276 <= (_zz_dataOut_payload_0_7274 ? _zz_dataOut_payload_0_7269 : _zz_dataOut_payload_0_7272);
    _zz_dataOut_payload_0_7277 <= (_zz_dataOut_payload_0_7274 ? _zz_dataOut_payload_0_7272 : _zz_dataOut_payload_0_7269);
    _zz_dataOut_payload_0_7278 <= (_zz_dataOut_payload_0_7275 ? _zz_dataOut_payload_0_7270 : _zz_dataOut_payload_0_7273);
    _zz_dataOut_payload_0_7279 <= (_zz_dataOut_payload_0_7275 ? _zz_dataOut_payload_0_7273 : _zz_dataOut_payload_0_7270);
    _zz_dataOut_payload_0_7288 <= (_zz_dataOut_payload_0_7286 ? _zz_dataOut_payload_0_7281 : _zz_dataOut_payload_0_7284);
    _zz_dataOut_payload_0_7289 <= (_zz_dataOut_payload_0_7286 ? _zz_dataOut_payload_0_7284 : _zz_dataOut_payload_0_7281);
    _zz_dataOut_payload_0_7290 <= (_zz_dataOut_payload_0_7287 ? _zz_dataOut_payload_0_7282 : _zz_dataOut_payload_0_7285);
    _zz_dataOut_payload_0_7291 <= (_zz_dataOut_payload_0_7287 ? _zz_dataOut_payload_0_7285 : _zz_dataOut_payload_0_7282);
    _zz_dataOut_payload_0_7292 <= _zz_dataOut_payload_0_7276;
    _zz_dataOut_payload_0_7293 <= _zz_dataOut_payload_0_7277;
    _zz_dataOut_payload_0_7294 <= _zz_dataOut_payload_0_7278;
    _zz_dataOut_payload_0_7295 <= _zz_dataOut_payload_0_7279;
    _zz_dataOut_payload_0_7296 <= _zz_dataOut_payload_0_7288;
    _zz_dataOut_payload_0_7297 <= _zz_dataOut_payload_0_7289;
    _zz_dataOut_payload_0_7298 <= _zz_dataOut_payload_0_7290;
    _zz_dataOut_payload_0_7299 <= _zz_dataOut_payload_0_7291;
    _zz_dataOut_payload_0_7320 <= (_zz_dataOut_payload_0_7318 ? _zz_dataOut_payload_0_7313 : _zz_dataOut_payload_0_7316);
    _zz_dataOut_payload_0_7321 <= (_zz_dataOut_payload_0_7318 ? _zz_dataOut_payload_0_7316 : _zz_dataOut_payload_0_7313);
    _zz_dataOut_payload_0_7322 <= (_zz_dataOut_payload_0_7319 ? _zz_dataOut_payload_0_7314 : _zz_dataOut_payload_0_7317);
    _zz_dataOut_payload_0_7323 <= (_zz_dataOut_payload_0_7319 ? _zz_dataOut_payload_0_7317 : _zz_dataOut_payload_0_7314);
    _zz_dataOut_payload_0_7332 <= (_zz_dataOut_payload_0_7330 ? _zz_dataOut_payload_0_7325 : _zz_dataOut_payload_0_7328);
    _zz_dataOut_payload_0_7333 <= (_zz_dataOut_payload_0_7330 ? _zz_dataOut_payload_0_7328 : _zz_dataOut_payload_0_7325);
    _zz_dataOut_payload_0_7334 <= (_zz_dataOut_payload_0_7331 ? _zz_dataOut_payload_0_7326 : _zz_dataOut_payload_0_7329);
    _zz_dataOut_payload_0_7335 <= (_zz_dataOut_payload_0_7331 ? _zz_dataOut_payload_0_7329 : _zz_dataOut_payload_0_7326);
    _zz_dataOut_payload_0_7336 <= _zz_dataOut_payload_0_7320;
    _zz_dataOut_payload_0_7337 <= _zz_dataOut_payload_0_7321;
    _zz_dataOut_payload_0_7338 <= _zz_dataOut_payload_0_7322;
    _zz_dataOut_payload_0_7339 <= _zz_dataOut_payload_0_7323;
    _zz_dataOut_payload_0_7340 <= _zz_dataOut_payload_0_7332;
    _zz_dataOut_payload_0_7341 <= _zz_dataOut_payload_0_7333;
    _zz_dataOut_payload_0_7342 <= _zz_dataOut_payload_0_7334;
    _zz_dataOut_payload_0_7343 <= _zz_dataOut_payload_0_7335;
    _zz_dataOut_payload_0_7344 <= _zz_dataOut_payload_0_7292;
    _zz_dataOut_payload_0_7345 <= _zz_dataOut_payload_0_7293;
    _zz_dataOut_payload_0_7346 <= _zz_dataOut_payload_0_7294;
    _zz_dataOut_payload_0_7347 <= _zz_dataOut_payload_0_7295;
    _zz_dataOut_payload_0_7348 <= _zz_dataOut_payload_0_7296;
    _zz_dataOut_payload_0_7349 <= _zz_dataOut_payload_0_7297;
    _zz_dataOut_payload_0_7350 <= _zz_dataOut_payload_0_7298;
    _zz_dataOut_payload_0_7351 <= _zz_dataOut_payload_0_7299;
    _zz_dataOut_payload_0_7352 <= _zz_dataOut_payload_0_7336;
    _zz_dataOut_payload_0_7353 <= _zz_dataOut_payload_0_7337;
    _zz_dataOut_payload_0_7354 <= _zz_dataOut_payload_0_7338;
    _zz_dataOut_payload_0_7355 <= _zz_dataOut_payload_0_7339;
    _zz_dataOut_payload_0_7356 <= _zz_dataOut_payload_0_7340;
    _zz_dataOut_payload_0_7357 <= _zz_dataOut_payload_0_7341;
    _zz_dataOut_payload_0_7358 <= _zz_dataOut_payload_0_7342;
    _zz_dataOut_payload_0_7359 <= _zz_dataOut_payload_0_7343;
    _zz_dataOut_payload_0_7360 <= _zz_dataOut_payload_0_7216;
    _zz_dataOut_payload_0_7361 <= _zz_dataOut_payload_0_7217;
    _zz_dataOut_payload_0_7362 <= _zz_dataOut_payload_0_7218;
    _zz_dataOut_payload_0_7363 <= _zz_dataOut_payload_0_7219;
    _zz_dataOut_payload_0_7364 <= _zz_dataOut_payload_0_7220;
    _zz_dataOut_payload_0_7365 <= _zz_dataOut_payload_0_7221;
    _zz_dataOut_payload_0_7366 <= _zz_dataOut_payload_0_7222;
    _zz_dataOut_payload_0_7367 <= _zz_dataOut_payload_0_7223;
    _zz_dataOut_payload_0_7368 <= _zz_dataOut_payload_0_7224;
    _zz_dataOut_payload_0_7369 <= _zz_dataOut_payload_0_7225;
    _zz_dataOut_payload_0_7370 <= _zz_dataOut_payload_0_7226;
    _zz_dataOut_payload_0_7371 <= _zz_dataOut_payload_0_7227;
    _zz_dataOut_payload_0_7372 <= _zz_dataOut_payload_0_7228;
    _zz_dataOut_payload_0_7373 <= _zz_dataOut_payload_0_7229;
    _zz_dataOut_payload_0_7374 <= _zz_dataOut_payload_0_7230;
    _zz_dataOut_payload_0_7375 <= _zz_dataOut_payload_0_7231;
    _zz_dataOut_payload_0_7376 <= _zz_dataOut_payload_0_7344;
    _zz_dataOut_payload_0_7377 <= _zz_dataOut_payload_0_7345;
    _zz_dataOut_payload_0_7378 <= _zz_dataOut_payload_0_7346;
    _zz_dataOut_payload_0_7379 <= _zz_dataOut_payload_0_7347;
    _zz_dataOut_payload_0_7380 <= _zz_dataOut_payload_0_7348;
    _zz_dataOut_payload_0_7381 <= _zz_dataOut_payload_0_7349;
    _zz_dataOut_payload_0_7382 <= _zz_dataOut_payload_0_7350;
    _zz_dataOut_payload_0_7383 <= _zz_dataOut_payload_0_7351;
    _zz_dataOut_payload_0_7384 <= _zz_dataOut_payload_0_7352;
    _zz_dataOut_payload_0_7385 <= _zz_dataOut_payload_0_7353;
    _zz_dataOut_payload_0_7386 <= _zz_dataOut_payload_0_7354;
    _zz_dataOut_payload_0_7387 <= _zz_dataOut_payload_0_7355;
    _zz_dataOut_payload_0_7388 <= _zz_dataOut_payload_0_7356;
    _zz_dataOut_payload_0_7389 <= _zz_dataOut_payload_0_7357;
    _zz_dataOut_payload_0_7390 <= _zz_dataOut_payload_0_7358;
    _zz_dataOut_payload_0_7391 <= _zz_dataOut_payload_0_7359;
    _zz_dataOut_payload_0_7484 <= (_zz_dataOut_payload_0_7482 ? _zz_dataOut_payload_0_7477 : _zz_dataOut_payload_0_7480);
    _zz_dataOut_payload_0_7485 <= (_zz_dataOut_payload_0_7482 ? _zz_dataOut_payload_0_7480 : _zz_dataOut_payload_0_7477);
    _zz_dataOut_payload_0_7486 <= (_zz_dataOut_payload_0_7483 ? _zz_dataOut_payload_0_7478 : _zz_dataOut_payload_0_7481);
    _zz_dataOut_payload_0_7487 <= (_zz_dataOut_payload_0_7483 ? _zz_dataOut_payload_0_7481 : _zz_dataOut_payload_0_7478);
    _zz_dataOut_payload_0_7496 <= (_zz_dataOut_payload_0_7494 ? _zz_dataOut_payload_0_7489 : _zz_dataOut_payload_0_7492);
    _zz_dataOut_payload_0_7497 <= (_zz_dataOut_payload_0_7494 ? _zz_dataOut_payload_0_7492 : _zz_dataOut_payload_0_7489);
    _zz_dataOut_payload_0_7498 <= (_zz_dataOut_payload_0_7495 ? _zz_dataOut_payload_0_7490 : _zz_dataOut_payload_0_7493);
    _zz_dataOut_payload_0_7499 <= (_zz_dataOut_payload_0_7495 ? _zz_dataOut_payload_0_7493 : _zz_dataOut_payload_0_7490);
    _zz_dataOut_payload_0_7500 <= _zz_dataOut_payload_0_7484;
    _zz_dataOut_payload_0_7501 <= _zz_dataOut_payload_0_7485;
    _zz_dataOut_payload_0_7502 <= _zz_dataOut_payload_0_7486;
    _zz_dataOut_payload_0_7503 <= _zz_dataOut_payload_0_7487;
    _zz_dataOut_payload_0_7504 <= _zz_dataOut_payload_0_7496;
    _zz_dataOut_payload_0_7505 <= _zz_dataOut_payload_0_7497;
    _zz_dataOut_payload_0_7506 <= _zz_dataOut_payload_0_7498;
    _zz_dataOut_payload_0_7507 <= _zz_dataOut_payload_0_7499;
    _zz_dataOut_payload_0_7528 <= (_zz_dataOut_payload_0_7526 ? _zz_dataOut_payload_0_7521 : _zz_dataOut_payload_0_7524);
    _zz_dataOut_payload_0_7529 <= (_zz_dataOut_payload_0_7526 ? _zz_dataOut_payload_0_7524 : _zz_dataOut_payload_0_7521);
    _zz_dataOut_payload_0_7530 <= (_zz_dataOut_payload_0_7527 ? _zz_dataOut_payload_0_7522 : _zz_dataOut_payload_0_7525);
    _zz_dataOut_payload_0_7531 <= (_zz_dataOut_payload_0_7527 ? _zz_dataOut_payload_0_7525 : _zz_dataOut_payload_0_7522);
    _zz_dataOut_payload_0_7540 <= (_zz_dataOut_payload_0_7538 ? _zz_dataOut_payload_0_7533 : _zz_dataOut_payload_0_7536);
    _zz_dataOut_payload_0_7541 <= (_zz_dataOut_payload_0_7538 ? _zz_dataOut_payload_0_7536 : _zz_dataOut_payload_0_7533);
    _zz_dataOut_payload_0_7542 <= (_zz_dataOut_payload_0_7539 ? _zz_dataOut_payload_0_7534 : _zz_dataOut_payload_0_7537);
    _zz_dataOut_payload_0_7543 <= (_zz_dataOut_payload_0_7539 ? _zz_dataOut_payload_0_7537 : _zz_dataOut_payload_0_7534);
    _zz_dataOut_payload_0_7544 <= _zz_dataOut_payload_0_7528;
    _zz_dataOut_payload_0_7545 <= _zz_dataOut_payload_0_7529;
    _zz_dataOut_payload_0_7546 <= _zz_dataOut_payload_0_7530;
    _zz_dataOut_payload_0_7547 <= _zz_dataOut_payload_0_7531;
    _zz_dataOut_payload_0_7548 <= _zz_dataOut_payload_0_7540;
    _zz_dataOut_payload_0_7549 <= _zz_dataOut_payload_0_7541;
    _zz_dataOut_payload_0_7550 <= _zz_dataOut_payload_0_7542;
    _zz_dataOut_payload_0_7551 <= _zz_dataOut_payload_0_7543;
    _zz_dataOut_payload_0_7552 <= _zz_dataOut_payload_0_7500;
    _zz_dataOut_payload_0_7553 <= _zz_dataOut_payload_0_7501;
    _zz_dataOut_payload_0_7554 <= _zz_dataOut_payload_0_7502;
    _zz_dataOut_payload_0_7555 <= _zz_dataOut_payload_0_7503;
    _zz_dataOut_payload_0_7556 <= _zz_dataOut_payload_0_7504;
    _zz_dataOut_payload_0_7557 <= _zz_dataOut_payload_0_7505;
    _zz_dataOut_payload_0_7558 <= _zz_dataOut_payload_0_7506;
    _zz_dataOut_payload_0_7559 <= _zz_dataOut_payload_0_7507;
    _zz_dataOut_payload_0_7560 <= _zz_dataOut_payload_0_7544;
    _zz_dataOut_payload_0_7561 <= _zz_dataOut_payload_0_7545;
    _zz_dataOut_payload_0_7562 <= _zz_dataOut_payload_0_7546;
    _zz_dataOut_payload_0_7563 <= _zz_dataOut_payload_0_7547;
    _zz_dataOut_payload_0_7564 <= _zz_dataOut_payload_0_7548;
    _zz_dataOut_payload_0_7565 <= _zz_dataOut_payload_0_7549;
    _zz_dataOut_payload_0_7566 <= _zz_dataOut_payload_0_7550;
    _zz_dataOut_payload_0_7567 <= _zz_dataOut_payload_0_7551;
    _zz_dataOut_payload_0_7612 <= (_zz_dataOut_payload_0_7610 ? _zz_dataOut_payload_0_7605 : _zz_dataOut_payload_0_7608);
    _zz_dataOut_payload_0_7613 <= (_zz_dataOut_payload_0_7610 ? _zz_dataOut_payload_0_7608 : _zz_dataOut_payload_0_7605);
    _zz_dataOut_payload_0_7614 <= (_zz_dataOut_payload_0_7611 ? _zz_dataOut_payload_0_7606 : _zz_dataOut_payload_0_7609);
    _zz_dataOut_payload_0_7615 <= (_zz_dataOut_payload_0_7611 ? _zz_dataOut_payload_0_7609 : _zz_dataOut_payload_0_7606);
    _zz_dataOut_payload_0_7624 <= (_zz_dataOut_payload_0_7622 ? _zz_dataOut_payload_0_7617 : _zz_dataOut_payload_0_7620);
    _zz_dataOut_payload_0_7625 <= (_zz_dataOut_payload_0_7622 ? _zz_dataOut_payload_0_7620 : _zz_dataOut_payload_0_7617);
    _zz_dataOut_payload_0_7626 <= (_zz_dataOut_payload_0_7623 ? _zz_dataOut_payload_0_7618 : _zz_dataOut_payload_0_7621);
    _zz_dataOut_payload_0_7627 <= (_zz_dataOut_payload_0_7623 ? _zz_dataOut_payload_0_7621 : _zz_dataOut_payload_0_7618);
    _zz_dataOut_payload_0_7628 <= _zz_dataOut_payload_0_7612;
    _zz_dataOut_payload_0_7629 <= _zz_dataOut_payload_0_7613;
    _zz_dataOut_payload_0_7630 <= _zz_dataOut_payload_0_7614;
    _zz_dataOut_payload_0_7631 <= _zz_dataOut_payload_0_7615;
    _zz_dataOut_payload_0_7632 <= _zz_dataOut_payload_0_7624;
    _zz_dataOut_payload_0_7633 <= _zz_dataOut_payload_0_7625;
    _zz_dataOut_payload_0_7634 <= _zz_dataOut_payload_0_7626;
    _zz_dataOut_payload_0_7635 <= _zz_dataOut_payload_0_7627;
    _zz_dataOut_payload_0_7656 <= (_zz_dataOut_payload_0_7654 ? _zz_dataOut_payload_0_7649 : _zz_dataOut_payload_0_7652);
    _zz_dataOut_payload_0_7657 <= (_zz_dataOut_payload_0_7654 ? _zz_dataOut_payload_0_7652 : _zz_dataOut_payload_0_7649);
    _zz_dataOut_payload_0_7658 <= (_zz_dataOut_payload_0_7655 ? _zz_dataOut_payload_0_7650 : _zz_dataOut_payload_0_7653);
    _zz_dataOut_payload_0_7659 <= (_zz_dataOut_payload_0_7655 ? _zz_dataOut_payload_0_7653 : _zz_dataOut_payload_0_7650);
    _zz_dataOut_payload_0_7668 <= (_zz_dataOut_payload_0_7666 ? _zz_dataOut_payload_0_7661 : _zz_dataOut_payload_0_7664);
    _zz_dataOut_payload_0_7669 <= (_zz_dataOut_payload_0_7666 ? _zz_dataOut_payload_0_7664 : _zz_dataOut_payload_0_7661);
    _zz_dataOut_payload_0_7670 <= (_zz_dataOut_payload_0_7667 ? _zz_dataOut_payload_0_7662 : _zz_dataOut_payload_0_7665);
    _zz_dataOut_payload_0_7671 <= (_zz_dataOut_payload_0_7667 ? _zz_dataOut_payload_0_7665 : _zz_dataOut_payload_0_7662);
    _zz_dataOut_payload_0_7672 <= _zz_dataOut_payload_0_7656;
    _zz_dataOut_payload_0_7673 <= _zz_dataOut_payload_0_7657;
    _zz_dataOut_payload_0_7674 <= _zz_dataOut_payload_0_7658;
    _zz_dataOut_payload_0_7675 <= _zz_dataOut_payload_0_7659;
    _zz_dataOut_payload_0_7676 <= _zz_dataOut_payload_0_7668;
    _zz_dataOut_payload_0_7677 <= _zz_dataOut_payload_0_7669;
    _zz_dataOut_payload_0_7678 <= _zz_dataOut_payload_0_7670;
    _zz_dataOut_payload_0_7679 <= _zz_dataOut_payload_0_7671;
    _zz_dataOut_payload_0_7680 <= _zz_dataOut_payload_0_7628;
    _zz_dataOut_payload_0_7681 <= _zz_dataOut_payload_0_7629;
    _zz_dataOut_payload_0_7682 <= _zz_dataOut_payload_0_7630;
    _zz_dataOut_payload_0_7683 <= _zz_dataOut_payload_0_7631;
    _zz_dataOut_payload_0_7684 <= _zz_dataOut_payload_0_7632;
    _zz_dataOut_payload_0_7685 <= _zz_dataOut_payload_0_7633;
    _zz_dataOut_payload_0_7686 <= _zz_dataOut_payload_0_7634;
    _zz_dataOut_payload_0_7687 <= _zz_dataOut_payload_0_7635;
    _zz_dataOut_payload_0_7688 <= _zz_dataOut_payload_0_7672;
    _zz_dataOut_payload_0_7689 <= _zz_dataOut_payload_0_7673;
    _zz_dataOut_payload_0_7690 <= _zz_dataOut_payload_0_7674;
    _zz_dataOut_payload_0_7691 <= _zz_dataOut_payload_0_7675;
    _zz_dataOut_payload_0_7692 <= _zz_dataOut_payload_0_7676;
    _zz_dataOut_payload_0_7693 <= _zz_dataOut_payload_0_7677;
    _zz_dataOut_payload_0_7694 <= _zz_dataOut_payload_0_7678;
    _zz_dataOut_payload_0_7695 <= _zz_dataOut_payload_0_7679;
    _zz_dataOut_payload_0_7696 <= _zz_dataOut_payload_0_7552;
    _zz_dataOut_payload_0_7697 <= _zz_dataOut_payload_0_7553;
    _zz_dataOut_payload_0_7698 <= _zz_dataOut_payload_0_7554;
    _zz_dataOut_payload_0_7699 <= _zz_dataOut_payload_0_7555;
    _zz_dataOut_payload_0_7700 <= _zz_dataOut_payload_0_7556;
    _zz_dataOut_payload_0_7701 <= _zz_dataOut_payload_0_7557;
    _zz_dataOut_payload_0_7702 <= _zz_dataOut_payload_0_7558;
    _zz_dataOut_payload_0_7703 <= _zz_dataOut_payload_0_7559;
    _zz_dataOut_payload_0_7704 <= _zz_dataOut_payload_0_7560;
    _zz_dataOut_payload_0_7705 <= _zz_dataOut_payload_0_7561;
    _zz_dataOut_payload_0_7706 <= _zz_dataOut_payload_0_7562;
    _zz_dataOut_payload_0_7707 <= _zz_dataOut_payload_0_7563;
    _zz_dataOut_payload_0_7708 <= _zz_dataOut_payload_0_7564;
    _zz_dataOut_payload_0_7709 <= _zz_dataOut_payload_0_7565;
    _zz_dataOut_payload_0_7710 <= _zz_dataOut_payload_0_7566;
    _zz_dataOut_payload_0_7711 <= _zz_dataOut_payload_0_7567;
    _zz_dataOut_payload_0_7712 <= _zz_dataOut_payload_0_7680;
    _zz_dataOut_payload_0_7713 <= _zz_dataOut_payload_0_7681;
    _zz_dataOut_payload_0_7714 <= _zz_dataOut_payload_0_7682;
    _zz_dataOut_payload_0_7715 <= _zz_dataOut_payload_0_7683;
    _zz_dataOut_payload_0_7716 <= _zz_dataOut_payload_0_7684;
    _zz_dataOut_payload_0_7717 <= _zz_dataOut_payload_0_7685;
    _zz_dataOut_payload_0_7718 <= _zz_dataOut_payload_0_7686;
    _zz_dataOut_payload_0_7719 <= _zz_dataOut_payload_0_7687;
    _zz_dataOut_payload_0_7720 <= _zz_dataOut_payload_0_7688;
    _zz_dataOut_payload_0_7721 <= _zz_dataOut_payload_0_7689;
    _zz_dataOut_payload_0_7722 <= _zz_dataOut_payload_0_7690;
    _zz_dataOut_payload_0_7723 <= _zz_dataOut_payload_0_7691;
    _zz_dataOut_payload_0_7724 <= _zz_dataOut_payload_0_7692;
    _zz_dataOut_payload_0_7725 <= _zz_dataOut_payload_0_7693;
    _zz_dataOut_payload_0_7726 <= _zz_dataOut_payload_0_7694;
    _zz_dataOut_payload_0_7727 <= _zz_dataOut_payload_0_7695;
    _zz_dataOut_payload_0_7820 <= (_zz_dataOut_payload_0_7818 ? _zz_dataOut_payload_0_7813 : _zz_dataOut_payload_0_7816);
    _zz_dataOut_payload_0_7821 <= (_zz_dataOut_payload_0_7818 ? _zz_dataOut_payload_0_7816 : _zz_dataOut_payload_0_7813);
    _zz_dataOut_payload_0_7822 <= (_zz_dataOut_payload_0_7819 ? _zz_dataOut_payload_0_7814 : _zz_dataOut_payload_0_7817);
    _zz_dataOut_payload_0_7823 <= (_zz_dataOut_payload_0_7819 ? _zz_dataOut_payload_0_7817 : _zz_dataOut_payload_0_7814);
    _zz_dataOut_payload_0_7832 <= (_zz_dataOut_payload_0_7830 ? _zz_dataOut_payload_0_7825 : _zz_dataOut_payload_0_7828);
    _zz_dataOut_payload_0_7833 <= (_zz_dataOut_payload_0_7830 ? _zz_dataOut_payload_0_7828 : _zz_dataOut_payload_0_7825);
    _zz_dataOut_payload_0_7834 <= (_zz_dataOut_payload_0_7831 ? _zz_dataOut_payload_0_7826 : _zz_dataOut_payload_0_7829);
    _zz_dataOut_payload_0_7835 <= (_zz_dataOut_payload_0_7831 ? _zz_dataOut_payload_0_7829 : _zz_dataOut_payload_0_7826);
    _zz_dataOut_payload_0_7836 <= _zz_dataOut_payload_0_7820;
    _zz_dataOut_payload_0_7837 <= _zz_dataOut_payload_0_7821;
    _zz_dataOut_payload_0_7838 <= _zz_dataOut_payload_0_7822;
    _zz_dataOut_payload_0_7839 <= _zz_dataOut_payload_0_7823;
    _zz_dataOut_payload_0_7840 <= _zz_dataOut_payload_0_7832;
    _zz_dataOut_payload_0_7841 <= _zz_dataOut_payload_0_7833;
    _zz_dataOut_payload_0_7842 <= _zz_dataOut_payload_0_7834;
    _zz_dataOut_payload_0_7843 <= _zz_dataOut_payload_0_7835;
    _zz_dataOut_payload_0_7864 <= (_zz_dataOut_payload_0_7862 ? _zz_dataOut_payload_0_7857 : _zz_dataOut_payload_0_7860);
    _zz_dataOut_payload_0_7865 <= (_zz_dataOut_payload_0_7862 ? _zz_dataOut_payload_0_7860 : _zz_dataOut_payload_0_7857);
    _zz_dataOut_payload_0_7866 <= (_zz_dataOut_payload_0_7863 ? _zz_dataOut_payload_0_7858 : _zz_dataOut_payload_0_7861);
    _zz_dataOut_payload_0_7867 <= (_zz_dataOut_payload_0_7863 ? _zz_dataOut_payload_0_7861 : _zz_dataOut_payload_0_7858);
    _zz_dataOut_payload_0_7876 <= (_zz_dataOut_payload_0_7874 ? _zz_dataOut_payload_0_7869 : _zz_dataOut_payload_0_7872);
    _zz_dataOut_payload_0_7877 <= (_zz_dataOut_payload_0_7874 ? _zz_dataOut_payload_0_7872 : _zz_dataOut_payload_0_7869);
    _zz_dataOut_payload_0_7878 <= (_zz_dataOut_payload_0_7875 ? _zz_dataOut_payload_0_7870 : _zz_dataOut_payload_0_7873);
    _zz_dataOut_payload_0_7879 <= (_zz_dataOut_payload_0_7875 ? _zz_dataOut_payload_0_7873 : _zz_dataOut_payload_0_7870);
    _zz_dataOut_payload_0_7880 <= _zz_dataOut_payload_0_7864;
    _zz_dataOut_payload_0_7881 <= _zz_dataOut_payload_0_7865;
    _zz_dataOut_payload_0_7882 <= _zz_dataOut_payload_0_7866;
    _zz_dataOut_payload_0_7883 <= _zz_dataOut_payload_0_7867;
    _zz_dataOut_payload_0_7884 <= _zz_dataOut_payload_0_7876;
    _zz_dataOut_payload_0_7885 <= _zz_dataOut_payload_0_7877;
    _zz_dataOut_payload_0_7886 <= _zz_dataOut_payload_0_7878;
    _zz_dataOut_payload_0_7887 <= _zz_dataOut_payload_0_7879;
    _zz_dataOut_payload_0_7888 <= _zz_dataOut_payload_0_7836;
    _zz_dataOut_payload_0_7889 <= _zz_dataOut_payload_0_7837;
    _zz_dataOut_payload_0_7890 <= _zz_dataOut_payload_0_7838;
    _zz_dataOut_payload_0_7891 <= _zz_dataOut_payload_0_7839;
    _zz_dataOut_payload_0_7892 <= _zz_dataOut_payload_0_7840;
    _zz_dataOut_payload_0_7893 <= _zz_dataOut_payload_0_7841;
    _zz_dataOut_payload_0_7894 <= _zz_dataOut_payload_0_7842;
    _zz_dataOut_payload_0_7895 <= _zz_dataOut_payload_0_7843;
    _zz_dataOut_payload_0_7896 <= _zz_dataOut_payload_0_7880;
    _zz_dataOut_payload_0_7897 <= _zz_dataOut_payload_0_7881;
    _zz_dataOut_payload_0_7898 <= _zz_dataOut_payload_0_7882;
    _zz_dataOut_payload_0_7899 <= _zz_dataOut_payload_0_7883;
    _zz_dataOut_payload_0_7900 <= _zz_dataOut_payload_0_7884;
    _zz_dataOut_payload_0_7901 <= _zz_dataOut_payload_0_7885;
    _zz_dataOut_payload_0_7902 <= _zz_dataOut_payload_0_7886;
    _zz_dataOut_payload_0_7903 <= _zz_dataOut_payload_0_7887;
    _zz_dataOut_payload_0_7948 <= (_zz_dataOut_payload_0_7946 ? _zz_dataOut_payload_0_7941 : _zz_dataOut_payload_0_7944);
    _zz_dataOut_payload_0_7949 <= (_zz_dataOut_payload_0_7946 ? _zz_dataOut_payload_0_7944 : _zz_dataOut_payload_0_7941);
    _zz_dataOut_payload_0_7950 <= (_zz_dataOut_payload_0_7947 ? _zz_dataOut_payload_0_7942 : _zz_dataOut_payload_0_7945);
    _zz_dataOut_payload_0_7951 <= (_zz_dataOut_payload_0_7947 ? _zz_dataOut_payload_0_7945 : _zz_dataOut_payload_0_7942);
    _zz_dataOut_payload_0_7960 <= (_zz_dataOut_payload_0_7958 ? _zz_dataOut_payload_0_7953 : _zz_dataOut_payload_0_7956);
    _zz_dataOut_payload_0_7961 <= (_zz_dataOut_payload_0_7958 ? _zz_dataOut_payload_0_7956 : _zz_dataOut_payload_0_7953);
    _zz_dataOut_payload_0_7962 <= (_zz_dataOut_payload_0_7959 ? _zz_dataOut_payload_0_7954 : _zz_dataOut_payload_0_7957);
    _zz_dataOut_payload_0_7963 <= (_zz_dataOut_payload_0_7959 ? _zz_dataOut_payload_0_7957 : _zz_dataOut_payload_0_7954);
    _zz_dataOut_payload_0_7964 <= _zz_dataOut_payload_0_7948;
    _zz_dataOut_payload_0_7965 <= _zz_dataOut_payload_0_7949;
    _zz_dataOut_payload_0_7966 <= _zz_dataOut_payload_0_7950;
    _zz_dataOut_payload_0_7967 <= _zz_dataOut_payload_0_7951;
    _zz_dataOut_payload_0_7968 <= _zz_dataOut_payload_0_7960;
    _zz_dataOut_payload_0_7969 <= _zz_dataOut_payload_0_7961;
    _zz_dataOut_payload_0_7970 <= _zz_dataOut_payload_0_7962;
    _zz_dataOut_payload_0_7971 <= _zz_dataOut_payload_0_7963;
    _zz_dataOut_payload_0_7992 <= (_zz_dataOut_payload_0_7990 ? _zz_dataOut_payload_0_7985 : _zz_dataOut_payload_0_7988);
    _zz_dataOut_payload_0_7993 <= (_zz_dataOut_payload_0_7990 ? _zz_dataOut_payload_0_7988 : _zz_dataOut_payload_0_7985);
    _zz_dataOut_payload_0_7994 <= (_zz_dataOut_payload_0_7991 ? _zz_dataOut_payload_0_7986 : _zz_dataOut_payload_0_7989);
    _zz_dataOut_payload_0_7995 <= (_zz_dataOut_payload_0_7991 ? _zz_dataOut_payload_0_7989 : _zz_dataOut_payload_0_7986);
    _zz_dataOut_payload_0_8004 <= (_zz_dataOut_payload_0_8002 ? _zz_dataOut_payload_0_7997 : _zz_dataOut_payload_0_8000);
    _zz_dataOut_payload_0_8005 <= (_zz_dataOut_payload_0_8002 ? _zz_dataOut_payload_0_8000 : _zz_dataOut_payload_0_7997);
    _zz_dataOut_payload_0_8006 <= (_zz_dataOut_payload_0_8003 ? _zz_dataOut_payload_0_7998 : _zz_dataOut_payload_0_8001);
    _zz_dataOut_payload_0_8007 <= (_zz_dataOut_payload_0_8003 ? _zz_dataOut_payload_0_8001 : _zz_dataOut_payload_0_7998);
    _zz_dataOut_payload_0_8008 <= _zz_dataOut_payload_0_7992;
    _zz_dataOut_payload_0_8009 <= _zz_dataOut_payload_0_7993;
    _zz_dataOut_payload_0_8010 <= _zz_dataOut_payload_0_7994;
    _zz_dataOut_payload_0_8011 <= _zz_dataOut_payload_0_7995;
    _zz_dataOut_payload_0_8012 <= _zz_dataOut_payload_0_8004;
    _zz_dataOut_payload_0_8013 <= _zz_dataOut_payload_0_8005;
    _zz_dataOut_payload_0_8014 <= _zz_dataOut_payload_0_8006;
    _zz_dataOut_payload_0_8015 <= _zz_dataOut_payload_0_8007;
    _zz_dataOut_payload_0_8016 <= _zz_dataOut_payload_0_7964;
    _zz_dataOut_payload_0_8017 <= _zz_dataOut_payload_0_7965;
    _zz_dataOut_payload_0_8018 <= _zz_dataOut_payload_0_7966;
    _zz_dataOut_payload_0_8019 <= _zz_dataOut_payload_0_7967;
    _zz_dataOut_payload_0_8020 <= _zz_dataOut_payload_0_7968;
    _zz_dataOut_payload_0_8021 <= _zz_dataOut_payload_0_7969;
    _zz_dataOut_payload_0_8022 <= _zz_dataOut_payload_0_7970;
    _zz_dataOut_payload_0_8023 <= _zz_dataOut_payload_0_7971;
    _zz_dataOut_payload_0_8024 <= _zz_dataOut_payload_0_8008;
    _zz_dataOut_payload_0_8025 <= _zz_dataOut_payload_0_8009;
    _zz_dataOut_payload_0_8026 <= _zz_dataOut_payload_0_8010;
    _zz_dataOut_payload_0_8027 <= _zz_dataOut_payload_0_8011;
    _zz_dataOut_payload_0_8028 <= _zz_dataOut_payload_0_8012;
    _zz_dataOut_payload_0_8029 <= _zz_dataOut_payload_0_8013;
    _zz_dataOut_payload_0_8030 <= _zz_dataOut_payload_0_8014;
    _zz_dataOut_payload_0_8031 <= _zz_dataOut_payload_0_8015;
    _zz_dataOut_payload_0_8032 <= _zz_dataOut_payload_0_7888;
    _zz_dataOut_payload_0_8033 <= _zz_dataOut_payload_0_7889;
    _zz_dataOut_payload_0_8034 <= _zz_dataOut_payload_0_7890;
    _zz_dataOut_payload_0_8035 <= _zz_dataOut_payload_0_7891;
    _zz_dataOut_payload_0_8036 <= _zz_dataOut_payload_0_7892;
    _zz_dataOut_payload_0_8037 <= _zz_dataOut_payload_0_7893;
    _zz_dataOut_payload_0_8038 <= _zz_dataOut_payload_0_7894;
    _zz_dataOut_payload_0_8039 <= _zz_dataOut_payload_0_7895;
    _zz_dataOut_payload_0_8040 <= _zz_dataOut_payload_0_7896;
    _zz_dataOut_payload_0_8041 <= _zz_dataOut_payload_0_7897;
    _zz_dataOut_payload_0_8042 <= _zz_dataOut_payload_0_7898;
    _zz_dataOut_payload_0_8043 <= _zz_dataOut_payload_0_7899;
    _zz_dataOut_payload_0_8044 <= _zz_dataOut_payload_0_7900;
    _zz_dataOut_payload_0_8045 <= _zz_dataOut_payload_0_7901;
    _zz_dataOut_payload_0_8046 <= _zz_dataOut_payload_0_7902;
    _zz_dataOut_payload_0_8047 <= _zz_dataOut_payload_0_7903;
    _zz_dataOut_payload_0_8048 <= _zz_dataOut_payload_0_8016;
    _zz_dataOut_payload_0_8049 <= _zz_dataOut_payload_0_8017;
    _zz_dataOut_payload_0_8050 <= _zz_dataOut_payload_0_8018;
    _zz_dataOut_payload_0_8051 <= _zz_dataOut_payload_0_8019;
    _zz_dataOut_payload_0_8052 <= _zz_dataOut_payload_0_8020;
    _zz_dataOut_payload_0_8053 <= _zz_dataOut_payload_0_8021;
    _zz_dataOut_payload_0_8054 <= _zz_dataOut_payload_0_8022;
    _zz_dataOut_payload_0_8055 <= _zz_dataOut_payload_0_8023;
    _zz_dataOut_payload_0_8056 <= _zz_dataOut_payload_0_8024;
    _zz_dataOut_payload_0_8057 <= _zz_dataOut_payload_0_8025;
    _zz_dataOut_payload_0_8058 <= _zz_dataOut_payload_0_8026;
    _zz_dataOut_payload_0_8059 <= _zz_dataOut_payload_0_8027;
    _zz_dataOut_payload_0_8060 <= _zz_dataOut_payload_0_8028;
    _zz_dataOut_payload_0_8061 <= _zz_dataOut_payload_0_8029;
    _zz_dataOut_payload_0_8062 <= _zz_dataOut_payload_0_8030;
    _zz_dataOut_payload_0_8063 <= _zz_dataOut_payload_0_8031;
    _zz_dataOut_payload_0_8064 <= _zz_dataOut_payload_0_5680;
    _zz_dataOut_payload_0_8065 <= _zz_dataOut_payload_0_5681;
    _zz_dataOut_payload_0_8066 <= _zz_dataOut_payload_0_5682;
    _zz_dataOut_payload_0_8067 <= _zz_dataOut_payload_0_5683;
    _zz_dataOut_payload_0_8068 <= _zz_dataOut_payload_0_5684;
    _zz_dataOut_payload_0_8069 <= _zz_dataOut_payload_0_5685;
    _zz_dataOut_payload_0_8070 <= _zz_dataOut_payload_0_5686;
    _zz_dataOut_payload_0_8071 <= _zz_dataOut_payload_0_5687;
    _zz_dataOut_payload_0_8072 <= _zz_dataOut_payload_0_5688;
    _zz_dataOut_payload_0_8073 <= _zz_dataOut_payload_0_5689;
    _zz_dataOut_payload_0_8074 <= _zz_dataOut_payload_0_5690;
    _zz_dataOut_payload_0_8075 <= _zz_dataOut_payload_0_5691;
    _zz_dataOut_payload_0_8076 <= _zz_dataOut_payload_0_5692;
    _zz_dataOut_payload_0_8077 <= _zz_dataOut_payload_0_5693;
    _zz_dataOut_payload_0_8078 <= _zz_dataOut_payload_0_5694;
    _zz_dataOut_payload_0_8079 <= _zz_dataOut_payload_0_5695;
    _zz_dataOut_payload_0_8080 <= _zz_dataOut_payload_0_5696;
    _zz_dataOut_payload_0_8081 <= _zz_dataOut_payload_0_5697;
    _zz_dataOut_payload_0_8082 <= _zz_dataOut_payload_0_5698;
    _zz_dataOut_payload_0_8083 <= _zz_dataOut_payload_0_5699;
    _zz_dataOut_payload_0_8084 <= _zz_dataOut_payload_0_5700;
    _zz_dataOut_payload_0_8085 <= _zz_dataOut_payload_0_5701;
    _zz_dataOut_payload_0_8086 <= _zz_dataOut_payload_0_5702;
    _zz_dataOut_payload_0_8087 <= _zz_dataOut_payload_0_5703;
    _zz_dataOut_payload_0_8088 <= _zz_dataOut_payload_0_5704;
    _zz_dataOut_payload_0_8089 <= _zz_dataOut_payload_0_5705;
    _zz_dataOut_payload_0_8090 <= _zz_dataOut_payload_0_5706;
    _zz_dataOut_payload_0_8091 <= _zz_dataOut_payload_0_5707;
    _zz_dataOut_payload_0_8092 <= _zz_dataOut_payload_0_5708;
    _zz_dataOut_payload_0_8093 <= _zz_dataOut_payload_0_5709;
    _zz_dataOut_payload_0_8094 <= _zz_dataOut_payload_0_5710;
    _zz_dataOut_payload_0_8095 <= _zz_dataOut_payload_0_5711;
    _zz_dataOut_payload_0_8096 <= _zz_dataOut_payload_0_6016;
    _zz_dataOut_payload_0_8097 <= _zz_dataOut_payload_0_6017;
    _zz_dataOut_payload_0_8098 <= _zz_dataOut_payload_0_6018;
    _zz_dataOut_payload_0_8099 <= _zz_dataOut_payload_0_6019;
    _zz_dataOut_payload_0_8100 <= _zz_dataOut_payload_0_6020;
    _zz_dataOut_payload_0_8101 <= _zz_dataOut_payload_0_6021;
    _zz_dataOut_payload_0_8102 <= _zz_dataOut_payload_0_6022;
    _zz_dataOut_payload_0_8103 <= _zz_dataOut_payload_0_6023;
    _zz_dataOut_payload_0_8104 <= _zz_dataOut_payload_0_6024;
    _zz_dataOut_payload_0_8105 <= _zz_dataOut_payload_0_6025;
    _zz_dataOut_payload_0_8106 <= _zz_dataOut_payload_0_6026;
    _zz_dataOut_payload_0_8107 <= _zz_dataOut_payload_0_6027;
    _zz_dataOut_payload_0_8108 <= _zz_dataOut_payload_0_6028;
    _zz_dataOut_payload_0_8109 <= _zz_dataOut_payload_0_6029;
    _zz_dataOut_payload_0_8110 <= _zz_dataOut_payload_0_6030;
    _zz_dataOut_payload_0_8111 <= _zz_dataOut_payload_0_6031;
    _zz_dataOut_payload_0_8112 <= _zz_dataOut_payload_0_6032;
    _zz_dataOut_payload_0_8113 <= _zz_dataOut_payload_0_6033;
    _zz_dataOut_payload_0_8114 <= _zz_dataOut_payload_0_6034;
    _zz_dataOut_payload_0_8115 <= _zz_dataOut_payload_0_6035;
    _zz_dataOut_payload_0_8116 <= _zz_dataOut_payload_0_6036;
    _zz_dataOut_payload_0_8117 <= _zz_dataOut_payload_0_6037;
    _zz_dataOut_payload_0_8118 <= _zz_dataOut_payload_0_6038;
    _zz_dataOut_payload_0_8119 <= _zz_dataOut_payload_0_6039;
    _zz_dataOut_payload_0_8120 <= _zz_dataOut_payload_0_6040;
    _zz_dataOut_payload_0_8121 <= _zz_dataOut_payload_0_6041;
    _zz_dataOut_payload_0_8122 <= _zz_dataOut_payload_0_6042;
    _zz_dataOut_payload_0_8123 <= _zz_dataOut_payload_0_6043;
    _zz_dataOut_payload_0_8124 <= _zz_dataOut_payload_0_6044;
    _zz_dataOut_payload_0_8125 <= _zz_dataOut_payload_0_6045;
    _zz_dataOut_payload_0_8126 <= _zz_dataOut_payload_0_6046;
    _zz_dataOut_payload_0_8127 <= _zz_dataOut_payload_0_6047;
    _zz_dataOut_payload_0_8128 <= _zz_dataOut_payload_0_6352;
    _zz_dataOut_payload_0_8129 <= _zz_dataOut_payload_0_6353;
    _zz_dataOut_payload_0_8130 <= _zz_dataOut_payload_0_6354;
    _zz_dataOut_payload_0_8131 <= _zz_dataOut_payload_0_6355;
    _zz_dataOut_payload_0_8132 <= _zz_dataOut_payload_0_6356;
    _zz_dataOut_payload_0_8133 <= _zz_dataOut_payload_0_6357;
    _zz_dataOut_payload_0_8134 <= _zz_dataOut_payload_0_6358;
    _zz_dataOut_payload_0_8135 <= _zz_dataOut_payload_0_6359;
    _zz_dataOut_payload_0_8136 <= _zz_dataOut_payload_0_6360;
    _zz_dataOut_payload_0_8137 <= _zz_dataOut_payload_0_6361;
    _zz_dataOut_payload_0_8138 <= _zz_dataOut_payload_0_6362;
    _zz_dataOut_payload_0_8139 <= _zz_dataOut_payload_0_6363;
    _zz_dataOut_payload_0_8140 <= _zz_dataOut_payload_0_6364;
    _zz_dataOut_payload_0_8141 <= _zz_dataOut_payload_0_6365;
    _zz_dataOut_payload_0_8142 <= _zz_dataOut_payload_0_6366;
    _zz_dataOut_payload_0_8143 <= _zz_dataOut_payload_0_6367;
    _zz_dataOut_payload_0_8144 <= _zz_dataOut_payload_0_6368;
    _zz_dataOut_payload_0_8145 <= _zz_dataOut_payload_0_6369;
    _zz_dataOut_payload_0_8146 <= _zz_dataOut_payload_0_6370;
    _zz_dataOut_payload_0_8147 <= _zz_dataOut_payload_0_6371;
    _zz_dataOut_payload_0_8148 <= _zz_dataOut_payload_0_6372;
    _zz_dataOut_payload_0_8149 <= _zz_dataOut_payload_0_6373;
    _zz_dataOut_payload_0_8150 <= _zz_dataOut_payload_0_6374;
    _zz_dataOut_payload_0_8151 <= _zz_dataOut_payload_0_6375;
    _zz_dataOut_payload_0_8152 <= _zz_dataOut_payload_0_6376;
    _zz_dataOut_payload_0_8153 <= _zz_dataOut_payload_0_6377;
    _zz_dataOut_payload_0_8154 <= _zz_dataOut_payload_0_6378;
    _zz_dataOut_payload_0_8155 <= _zz_dataOut_payload_0_6379;
    _zz_dataOut_payload_0_8156 <= _zz_dataOut_payload_0_6380;
    _zz_dataOut_payload_0_8157 <= _zz_dataOut_payload_0_6381;
    _zz_dataOut_payload_0_8158 <= _zz_dataOut_payload_0_6382;
    _zz_dataOut_payload_0_8159 <= _zz_dataOut_payload_0_6383;
    _zz_dataOut_payload_0_8160 <= _zz_dataOut_payload_0_6688;
    _zz_dataOut_payload_0_8161 <= _zz_dataOut_payload_0_6689;
    _zz_dataOut_payload_0_8162 <= _zz_dataOut_payload_0_6690;
    _zz_dataOut_payload_0_8163 <= _zz_dataOut_payload_0_6691;
    _zz_dataOut_payload_0_8164 <= _zz_dataOut_payload_0_6692;
    _zz_dataOut_payload_0_8165 <= _zz_dataOut_payload_0_6693;
    _zz_dataOut_payload_0_8166 <= _zz_dataOut_payload_0_6694;
    _zz_dataOut_payload_0_8167 <= _zz_dataOut_payload_0_6695;
    _zz_dataOut_payload_0_8168 <= _zz_dataOut_payload_0_6696;
    _zz_dataOut_payload_0_8169 <= _zz_dataOut_payload_0_6697;
    _zz_dataOut_payload_0_8170 <= _zz_dataOut_payload_0_6698;
    _zz_dataOut_payload_0_8171 <= _zz_dataOut_payload_0_6699;
    _zz_dataOut_payload_0_8172 <= _zz_dataOut_payload_0_6700;
    _zz_dataOut_payload_0_8173 <= _zz_dataOut_payload_0_6701;
    _zz_dataOut_payload_0_8174 <= _zz_dataOut_payload_0_6702;
    _zz_dataOut_payload_0_8175 <= _zz_dataOut_payload_0_6703;
    _zz_dataOut_payload_0_8176 <= _zz_dataOut_payload_0_6704;
    _zz_dataOut_payload_0_8177 <= _zz_dataOut_payload_0_6705;
    _zz_dataOut_payload_0_8178 <= _zz_dataOut_payload_0_6706;
    _zz_dataOut_payload_0_8179 <= _zz_dataOut_payload_0_6707;
    _zz_dataOut_payload_0_8180 <= _zz_dataOut_payload_0_6708;
    _zz_dataOut_payload_0_8181 <= _zz_dataOut_payload_0_6709;
    _zz_dataOut_payload_0_8182 <= _zz_dataOut_payload_0_6710;
    _zz_dataOut_payload_0_8183 <= _zz_dataOut_payload_0_6711;
    _zz_dataOut_payload_0_8184 <= _zz_dataOut_payload_0_6712;
    _zz_dataOut_payload_0_8185 <= _zz_dataOut_payload_0_6713;
    _zz_dataOut_payload_0_8186 <= _zz_dataOut_payload_0_6714;
    _zz_dataOut_payload_0_8187 <= _zz_dataOut_payload_0_6715;
    _zz_dataOut_payload_0_8188 <= _zz_dataOut_payload_0_6716;
    _zz_dataOut_payload_0_8189 <= _zz_dataOut_payload_0_6717;
    _zz_dataOut_payload_0_8190 <= _zz_dataOut_payload_0_6718;
    _zz_dataOut_payload_0_8191 <= _zz_dataOut_payload_0_6719;
    _zz_dataOut_payload_0_8192 <= _zz_dataOut_payload_0_7024;
    _zz_dataOut_payload_0_8193 <= _zz_dataOut_payload_0_7025;
    _zz_dataOut_payload_0_8194 <= _zz_dataOut_payload_0_7026;
    _zz_dataOut_payload_0_8195 <= _zz_dataOut_payload_0_7027;
    _zz_dataOut_payload_0_8196 <= _zz_dataOut_payload_0_7028;
    _zz_dataOut_payload_0_8197 <= _zz_dataOut_payload_0_7029;
    _zz_dataOut_payload_0_8198 <= _zz_dataOut_payload_0_7030;
    _zz_dataOut_payload_0_8199 <= _zz_dataOut_payload_0_7031;
    _zz_dataOut_payload_0_8200 <= _zz_dataOut_payload_0_7032;
    _zz_dataOut_payload_0_8201 <= _zz_dataOut_payload_0_7033;
    _zz_dataOut_payload_0_8202 <= _zz_dataOut_payload_0_7034;
    _zz_dataOut_payload_0_8203 <= _zz_dataOut_payload_0_7035;
    _zz_dataOut_payload_0_8204 <= _zz_dataOut_payload_0_7036;
    _zz_dataOut_payload_0_8205 <= _zz_dataOut_payload_0_7037;
    _zz_dataOut_payload_0_8206 <= _zz_dataOut_payload_0_7038;
    _zz_dataOut_payload_0_8207 <= _zz_dataOut_payload_0_7039;
    _zz_dataOut_payload_0_8208 <= _zz_dataOut_payload_0_7040;
    _zz_dataOut_payload_0_8209 <= _zz_dataOut_payload_0_7041;
    _zz_dataOut_payload_0_8210 <= _zz_dataOut_payload_0_7042;
    _zz_dataOut_payload_0_8211 <= _zz_dataOut_payload_0_7043;
    _zz_dataOut_payload_0_8212 <= _zz_dataOut_payload_0_7044;
    _zz_dataOut_payload_0_8213 <= _zz_dataOut_payload_0_7045;
    _zz_dataOut_payload_0_8214 <= _zz_dataOut_payload_0_7046;
    _zz_dataOut_payload_0_8215 <= _zz_dataOut_payload_0_7047;
    _zz_dataOut_payload_0_8216 <= _zz_dataOut_payload_0_7048;
    _zz_dataOut_payload_0_8217 <= _zz_dataOut_payload_0_7049;
    _zz_dataOut_payload_0_8218 <= _zz_dataOut_payload_0_7050;
    _zz_dataOut_payload_0_8219 <= _zz_dataOut_payload_0_7051;
    _zz_dataOut_payload_0_8220 <= _zz_dataOut_payload_0_7052;
    _zz_dataOut_payload_0_8221 <= _zz_dataOut_payload_0_7053;
    _zz_dataOut_payload_0_8222 <= _zz_dataOut_payload_0_7054;
    _zz_dataOut_payload_0_8223 <= _zz_dataOut_payload_0_7055;
    _zz_dataOut_payload_0_8224 <= _zz_dataOut_payload_0_7360;
    _zz_dataOut_payload_0_8225 <= _zz_dataOut_payload_0_7361;
    _zz_dataOut_payload_0_8226 <= _zz_dataOut_payload_0_7362;
    _zz_dataOut_payload_0_8227 <= _zz_dataOut_payload_0_7363;
    _zz_dataOut_payload_0_8228 <= _zz_dataOut_payload_0_7364;
    _zz_dataOut_payload_0_8229 <= _zz_dataOut_payload_0_7365;
    _zz_dataOut_payload_0_8230 <= _zz_dataOut_payload_0_7366;
    _zz_dataOut_payload_0_8231 <= _zz_dataOut_payload_0_7367;
    _zz_dataOut_payload_0_8232 <= _zz_dataOut_payload_0_7368;
    _zz_dataOut_payload_0_8233 <= _zz_dataOut_payload_0_7369;
    _zz_dataOut_payload_0_8234 <= _zz_dataOut_payload_0_7370;
    _zz_dataOut_payload_0_8235 <= _zz_dataOut_payload_0_7371;
    _zz_dataOut_payload_0_8236 <= _zz_dataOut_payload_0_7372;
    _zz_dataOut_payload_0_8237 <= _zz_dataOut_payload_0_7373;
    _zz_dataOut_payload_0_8238 <= _zz_dataOut_payload_0_7374;
    _zz_dataOut_payload_0_8239 <= _zz_dataOut_payload_0_7375;
    _zz_dataOut_payload_0_8240 <= _zz_dataOut_payload_0_7376;
    _zz_dataOut_payload_0_8241 <= _zz_dataOut_payload_0_7377;
    _zz_dataOut_payload_0_8242 <= _zz_dataOut_payload_0_7378;
    _zz_dataOut_payload_0_8243 <= _zz_dataOut_payload_0_7379;
    _zz_dataOut_payload_0_8244 <= _zz_dataOut_payload_0_7380;
    _zz_dataOut_payload_0_8245 <= _zz_dataOut_payload_0_7381;
    _zz_dataOut_payload_0_8246 <= _zz_dataOut_payload_0_7382;
    _zz_dataOut_payload_0_8247 <= _zz_dataOut_payload_0_7383;
    _zz_dataOut_payload_0_8248 <= _zz_dataOut_payload_0_7384;
    _zz_dataOut_payload_0_8249 <= _zz_dataOut_payload_0_7385;
    _zz_dataOut_payload_0_8250 <= _zz_dataOut_payload_0_7386;
    _zz_dataOut_payload_0_8251 <= _zz_dataOut_payload_0_7387;
    _zz_dataOut_payload_0_8252 <= _zz_dataOut_payload_0_7388;
    _zz_dataOut_payload_0_8253 <= _zz_dataOut_payload_0_7389;
    _zz_dataOut_payload_0_8254 <= _zz_dataOut_payload_0_7390;
    _zz_dataOut_payload_0_8255 <= _zz_dataOut_payload_0_7391;
    _zz_dataOut_payload_0_8256 <= _zz_dataOut_payload_0_7696;
    _zz_dataOut_payload_0_8257 <= _zz_dataOut_payload_0_7697;
    _zz_dataOut_payload_0_8258 <= _zz_dataOut_payload_0_7698;
    _zz_dataOut_payload_0_8259 <= _zz_dataOut_payload_0_7699;
    _zz_dataOut_payload_0_8260 <= _zz_dataOut_payload_0_7700;
    _zz_dataOut_payload_0_8261 <= _zz_dataOut_payload_0_7701;
    _zz_dataOut_payload_0_8262 <= _zz_dataOut_payload_0_7702;
    _zz_dataOut_payload_0_8263 <= _zz_dataOut_payload_0_7703;
    _zz_dataOut_payload_0_8264 <= _zz_dataOut_payload_0_7704;
    _zz_dataOut_payload_0_8265 <= _zz_dataOut_payload_0_7705;
    _zz_dataOut_payload_0_8266 <= _zz_dataOut_payload_0_7706;
    _zz_dataOut_payload_0_8267 <= _zz_dataOut_payload_0_7707;
    _zz_dataOut_payload_0_8268 <= _zz_dataOut_payload_0_7708;
    _zz_dataOut_payload_0_8269 <= _zz_dataOut_payload_0_7709;
    _zz_dataOut_payload_0_8270 <= _zz_dataOut_payload_0_7710;
    _zz_dataOut_payload_0_8271 <= _zz_dataOut_payload_0_7711;
    _zz_dataOut_payload_0_8272 <= _zz_dataOut_payload_0_7712;
    _zz_dataOut_payload_0_8273 <= _zz_dataOut_payload_0_7713;
    _zz_dataOut_payload_0_8274 <= _zz_dataOut_payload_0_7714;
    _zz_dataOut_payload_0_8275 <= _zz_dataOut_payload_0_7715;
    _zz_dataOut_payload_0_8276 <= _zz_dataOut_payload_0_7716;
    _zz_dataOut_payload_0_8277 <= _zz_dataOut_payload_0_7717;
    _zz_dataOut_payload_0_8278 <= _zz_dataOut_payload_0_7718;
    _zz_dataOut_payload_0_8279 <= _zz_dataOut_payload_0_7719;
    _zz_dataOut_payload_0_8280 <= _zz_dataOut_payload_0_7720;
    _zz_dataOut_payload_0_8281 <= _zz_dataOut_payload_0_7721;
    _zz_dataOut_payload_0_8282 <= _zz_dataOut_payload_0_7722;
    _zz_dataOut_payload_0_8283 <= _zz_dataOut_payload_0_7723;
    _zz_dataOut_payload_0_8284 <= _zz_dataOut_payload_0_7724;
    _zz_dataOut_payload_0_8285 <= _zz_dataOut_payload_0_7725;
    _zz_dataOut_payload_0_8286 <= _zz_dataOut_payload_0_7726;
    _zz_dataOut_payload_0_8287 <= _zz_dataOut_payload_0_7727;
    _zz_dataOut_payload_0_8288 <= _zz_dataOut_payload_0_8032;
    _zz_dataOut_payload_0_8289 <= _zz_dataOut_payload_0_8033;
    _zz_dataOut_payload_0_8290 <= _zz_dataOut_payload_0_8034;
    _zz_dataOut_payload_0_8291 <= _zz_dataOut_payload_0_8035;
    _zz_dataOut_payload_0_8292 <= _zz_dataOut_payload_0_8036;
    _zz_dataOut_payload_0_8293 <= _zz_dataOut_payload_0_8037;
    _zz_dataOut_payload_0_8294 <= _zz_dataOut_payload_0_8038;
    _zz_dataOut_payload_0_8295 <= _zz_dataOut_payload_0_8039;
    _zz_dataOut_payload_0_8296 <= _zz_dataOut_payload_0_8040;
    _zz_dataOut_payload_0_8297 <= _zz_dataOut_payload_0_8041;
    _zz_dataOut_payload_0_8298 <= _zz_dataOut_payload_0_8042;
    _zz_dataOut_payload_0_8299 <= _zz_dataOut_payload_0_8043;
    _zz_dataOut_payload_0_8300 <= _zz_dataOut_payload_0_8044;
    _zz_dataOut_payload_0_8301 <= _zz_dataOut_payload_0_8045;
    _zz_dataOut_payload_0_8302 <= _zz_dataOut_payload_0_8046;
    _zz_dataOut_payload_0_8303 <= _zz_dataOut_payload_0_8047;
    _zz_dataOut_payload_0_8304 <= _zz_dataOut_payload_0_8048;
    _zz_dataOut_payload_0_8305 <= _zz_dataOut_payload_0_8049;
    _zz_dataOut_payload_0_8306 <= _zz_dataOut_payload_0_8050;
    _zz_dataOut_payload_0_8307 <= _zz_dataOut_payload_0_8051;
    _zz_dataOut_payload_0_8308 <= _zz_dataOut_payload_0_8052;
    _zz_dataOut_payload_0_8309 <= _zz_dataOut_payload_0_8053;
    _zz_dataOut_payload_0_8310 <= _zz_dataOut_payload_0_8054;
    _zz_dataOut_payload_0_8311 <= _zz_dataOut_payload_0_8055;
    _zz_dataOut_payload_0_8312 <= _zz_dataOut_payload_0_8056;
    _zz_dataOut_payload_0_8313 <= _zz_dataOut_payload_0_8057;
    _zz_dataOut_payload_0_8314 <= _zz_dataOut_payload_0_8058;
    _zz_dataOut_payload_0_8315 <= _zz_dataOut_payload_0_8059;
    _zz_dataOut_payload_0_8316 <= _zz_dataOut_payload_0_8060;
    _zz_dataOut_payload_0_8317 <= _zz_dataOut_payload_0_8061;
    _zz_dataOut_payload_0_8318 <= _zz_dataOut_payload_0_8062;
    _zz_dataOut_payload_0_8319 <= _zz_dataOut_payload_0_8063;
    _zz_dataOut_payload_0_8508 <= (_zz_dataOut_payload_0_8506 ? _zz_dataOut_payload_0_8501 : _zz_dataOut_payload_0_8504);
    _zz_dataOut_payload_0_8509 <= (_zz_dataOut_payload_0_8506 ? _zz_dataOut_payload_0_8504 : _zz_dataOut_payload_0_8501);
    _zz_dataOut_payload_0_8510 <= (_zz_dataOut_payload_0_8507 ? _zz_dataOut_payload_0_8502 : _zz_dataOut_payload_0_8505);
    _zz_dataOut_payload_0_8511 <= (_zz_dataOut_payload_0_8507 ? _zz_dataOut_payload_0_8505 : _zz_dataOut_payload_0_8502);
    _zz_dataOut_payload_0_8520 <= (_zz_dataOut_payload_0_8518 ? _zz_dataOut_payload_0_8513 : _zz_dataOut_payload_0_8516);
    _zz_dataOut_payload_0_8521 <= (_zz_dataOut_payload_0_8518 ? _zz_dataOut_payload_0_8516 : _zz_dataOut_payload_0_8513);
    _zz_dataOut_payload_0_8522 <= (_zz_dataOut_payload_0_8519 ? _zz_dataOut_payload_0_8514 : _zz_dataOut_payload_0_8517);
    _zz_dataOut_payload_0_8523 <= (_zz_dataOut_payload_0_8519 ? _zz_dataOut_payload_0_8517 : _zz_dataOut_payload_0_8514);
    _zz_dataOut_payload_0_8524 <= _zz_dataOut_payload_0_8508;
    _zz_dataOut_payload_0_8525 <= _zz_dataOut_payload_0_8509;
    _zz_dataOut_payload_0_8526 <= _zz_dataOut_payload_0_8510;
    _zz_dataOut_payload_0_8527 <= _zz_dataOut_payload_0_8511;
    _zz_dataOut_payload_0_8528 <= _zz_dataOut_payload_0_8520;
    _zz_dataOut_payload_0_8529 <= _zz_dataOut_payload_0_8521;
    _zz_dataOut_payload_0_8530 <= _zz_dataOut_payload_0_8522;
    _zz_dataOut_payload_0_8531 <= _zz_dataOut_payload_0_8523;
    _zz_dataOut_payload_0_8552 <= (_zz_dataOut_payload_0_8550 ? _zz_dataOut_payload_0_8545 : _zz_dataOut_payload_0_8548);
    _zz_dataOut_payload_0_8553 <= (_zz_dataOut_payload_0_8550 ? _zz_dataOut_payload_0_8548 : _zz_dataOut_payload_0_8545);
    _zz_dataOut_payload_0_8554 <= (_zz_dataOut_payload_0_8551 ? _zz_dataOut_payload_0_8546 : _zz_dataOut_payload_0_8549);
    _zz_dataOut_payload_0_8555 <= (_zz_dataOut_payload_0_8551 ? _zz_dataOut_payload_0_8549 : _zz_dataOut_payload_0_8546);
    _zz_dataOut_payload_0_8564 <= (_zz_dataOut_payload_0_8562 ? _zz_dataOut_payload_0_8557 : _zz_dataOut_payload_0_8560);
    _zz_dataOut_payload_0_8565 <= (_zz_dataOut_payload_0_8562 ? _zz_dataOut_payload_0_8560 : _zz_dataOut_payload_0_8557);
    _zz_dataOut_payload_0_8566 <= (_zz_dataOut_payload_0_8563 ? _zz_dataOut_payload_0_8558 : _zz_dataOut_payload_0_8561);
    _zz_dataOut_payload_0_8567 <= (_zz_dataOut_payload_0_8563 ? _zz_dataOut_payload_0_8561 : _zz_dataOut_payload_0_8558);
    _zz_dataOut_payload_0_8568 <= _zz_dataOut_payload_0_8552;
    _zz_dataOut_payload_0_8569 <= _zz_dataOut_payload_0_8553;
    _zz_dataOut_payload_0_8570 <= _zz_dataOut_payload_0_8554;
    _zz_dataOut_payload_0_8571 <= _zz_dataOut_payload_0_8555;
    _zz_dataOut_payload_0_8572 <= _zz_dataOut_payload_0_8564;
    _zz_dataOut_payload_0_8573 <= _zz_dataOut_payload_0_8565;
    _zz_dataOut_payload_0_8574 <= _zz_dataOut_payload_0_8566;
    _zz_dataOut_payload_0_8575 <= _zz_dataOut_payload_0_8567;
    _zz_dataOut_payload_0_8576 <= _zz_dataOut_payload_0_8524;
    _zz_dataOut_payload_0_8577 <= _zz_dataOut_payload_0_8525;
    _zz_dataOut_payload_0_8578 <= _zz_dataOut_payload_0_8526;
    _zz_dataOut_payload_0_8579 <= _zz_dataOut_payload_0_8527;
    _zz_dataOut_payload_0_8580 <= _zz_dataOut_payload_0_8528;
    _zz_dataOut_payload_0_8581 <= _zz_dataOut_payload_0_8529;
    _zz_dataOut_payload_0_8582 <= _zz_dataOut_payload_0_8530;
    _zz_dataOut_payload_0_8583 <= _zz_dataOut_payload_0_8531;
    _zz_dataOut_payload_0_8584 <= _zz_dataOut_payload_0_8568;
    _zz_dataOut_payload_0_8585 <= _zz_dataOut_payload_0_8569;
    _zz_dataOut_payload_0_8586 <= _zz_dataOut_payload_0_8570;
    _zz_dataOut_payload_0_8587 <= _zz_dataOut_payload_0_8571;
    _zz_dataOut_payload_0_8588 <= _zz_dataOut_payload_0_8572;
    _zz_dataOut_payload_0_8589 <= _zz_dataOut_payload_0_8573;
    _zz_dataOut_payload_0_8590 <= _zz_dataOut_payload_0_8574;
    _zz_dataOut_payload_0_8591 <= _zz_dataOut_payload_0_8575;
    _zz_dataOut_payload_0_8636 <= (_zz_dataOut_payload_0_8634 ? _zz_dataOut_payload_0_8629 : _zz_dataOut_payload_0_8632);
    _zz_dataOut_payload_0_8637 <= (_zz_dataOut_payload_0_8634 ? _zz_dataOut_payload_0_8632 : _zz_dataOut_payload_0_8629);
    _zz_dataOut_payload_0_8638 <= (_zz_dataOut_payload_0_8635 ? _zz_dataOut_payload_0_8630 : _zz_dataOut_payload_0_8633);
    _zz_dataOut_payload_0_8639 <= (_zz_dataOut_payload_0_8635 ? _zz_dataOut_payload_0_8633 : _zz_dataOut_payload_0_8630);
    _zz_dataOut_payload_0_8648 <= (_zz_dataOut_payload_0_8646 ? _zz_dataOut_payload_0_8641 : _zz_dataOut_payload_0_8644);
    _zz_dataOut_payload_0_8649 <= (_zz_dataOut_payload_0_8646 ? _zz_dataOut_payload_0_8644 : _zz_dataOut_payload_0_8641);
    _zz_dataOut_payload_0_8650 <= (_zz_dataOut_payload_0_8647 ? _zz_dataOut_payload_0_8642 : _zz_dataOut_payload_0_8645);
    _zz_dataOut_payload_0_8651 <= (_zz_dataOut_payload_0_8647 ? _zz_dataOut_payload_0_8645 : _zz_dataOut_payload_0_8642);
    _zz_dataOut_payload_0_8652 <= _zz_dataOut_payload_0_8636;
    _zz_dataOut_payload_0_8653 <= _zz_dataOut_payload_0_8637;
    _zz_dataOut_payload_0_8654 <= _zz_dataOut_payload_0_8638;
    _zz_dataOut_payload_0_8655 <= _zz_dataOut_payload_0_8639;
    _zz_dataOut_payload_0_8656 <= _zz_dataOut_payload_0_8648;
    _zz_dataOut_payload_0_8657 <= _zz_dataOut_payload_0_8649;
    _zz_dataOut_payload_0_8658 <= _zz_dataOut_payload_0_8650;
    _zz_dataOut_payload_0_8659 <= _zz_dataOut_payload_0_8651;
    _zz_dataOut_payload_0_8680 <= (_zz_dataOut_payload_0_8678 ? _zz_dataOut_payload_0_8673 : _zz_dataOut_payload_0_8676);
    _zz_dataOut_payload_0_8681 <= (_zz_dataOut_payload_0_8678 ? _zz_dataOut_payload_0_8676 : _zz_dataOut_payload_0_8673);
    _zz_dataOut_payload_0_8682 <= (_zz_dataOut_payload_0_8679 ? _zz_dataOut_payload_0_8674 : _zz_dataOut_payload_0_8677);
    _zz_dataOut_payload_0_8683 <= (_zz_dataOut_payload_0_8679 ? _zz_dataOut_payload_0_8677 : _zz_dataOut_payload_0_8674);
    _zz_dataOut_payload_0_8692 <= (_zz_dataOut_payload_0_8690 ? _zz_dataOut_payload_0_8685 : _zz_dataOut_payload_0_8688);
    _zz_dataOut_payload_0_8693 <= (_zz_dataOut_payload_0_8690 ? _zz_dataOut_payload_0_8688 : _zz_dataOut_payload_0_8685);
    _zz_dataOut_payload_0_8694 <= (_zz_dataOut_payload_0_8691 ? _zz_dataOut_payload_0_8686 : _zz_dataOut_payload_0_8689);
    _zz_dataOut_payload_0_8695 <= (_zz_dataOut_payload_0_8691 ? _zz_dataOut_payload_0_8689 : _zz_dataOut_payload_0_8686);
    _zz_dataOut_payload_0_8696 <= _zz_dataOut_payload_0_8680;
    _zz_dataOut_payload_0_8697 <= _zz_dataOut_payload_0_8681;
    _zz_dataOut_payload_0_8698 <= _zz_dataOut_payload_0_8682;
    _zz_dataOut_payload_0_8699 <= _zz_dataOut_payload_0_8683;
    _zz_dataOut_payload_0_8700 <= _zz_dataOut_payload_0_8692;
    _zz_dataOut_payload_0_8701 <= _zz_dataOut_payload_0_8693;
    _zz_dataOut_payload_0_8702 <= _zz_dataOut_payload_0_8694;
    _zz_dataOut_payload_0_8703 <= _zz_dataOut_payload_0_8695;
    _zz_dataOut_payload_0_8704 <= _zz_dataOut_payload_0_8652;
    _zz_dataOut_payload_0_8705 <= _zz_dataOut_payload_0_8653;
    _zz_dataOut_payload_0_8706 <= _zz_dataOut_payload_0_8654;
    _zz_dataOut_payload_0_8707 <= _zz_dataOut_payload_0_8655;
    _zz_dataOut_payload_0_8708 <= _zz_dataOut_payload_0_8656;
    _zz_dataOut_payload_0_8709 <= _zz_dataOut_payload_0_8657;
    _zz_dataOut_payload_0_8710 <= _zz_dataOut_payload_0_8658;
    _zz_dataOut_payload_0_8711 <= _zz_dataOut_payload_0_8659;
    _zz_dataOut_payload_0_8712 <= _zz_dataOut_payload_0_8696;
    _zz_dataOut_payload_0_8713 <= _zz_dataOut_payload_0_8697;
    _zz_dataOut_payload_0_8714 <= _zz_dataOut_payload_0_8698;
    _zz_dataOut_payload_0_8715 <= _zz_dataOut_payload_0_8699;
    _zz_dataOut_payload_0_8716 <= _zz_dataOut_payload_0_8700;
    _zz_dataOut_payload_0_8717 <= _zz_dataOut_payload_0_8701;
    _zz_dataOut_payload_0_8718 <= _zz_dataOut_payload_0_8702;
    _zz_dataOut_payload_0_8719 <= _zz_dataOut_payload_0_8703;
    _zz_dataOut_payload_0_8720 <= _zz_dataOut_payload_0_8576;
    _zz_dataOut_payload_0_8721 <= _zz_dataOut_payload_0_8577;
    _zz_dataOut_payload_0_8722 <= _zz_dataOut_payload_0_8578;
    _zz_dataOut_payload_0_8723 <= _zz_dataOut_payload_0_8579;
    _zz_dataOut_payload_0_8724 <= _zz_dataOut_payload_0_8580;
    _zz_dataOut_payload_0_8725 <= _zz_dataOut_payload_0_8581;
    _zz_dataOut_payload_0_8726 <= _zz_dataOut_payload_0_8582;
    _zz_dataOut_payload_0_8727 <= _zz_dataOut_payload_0_8583;
    _zz_dataOut_payload_0_8728 <= _zz_dataOut_payload_0_8584;
    _zz_dataOut_payload_0_8729 <= _zz_dataOut_payload_0_8585;
    _zz_dataOut_payload_0_8730 <= _zz_dataOut_payload_0_8586;
    _zz_dataOut_payload_0_8731 <= _zz_dataOut_payload_0_8587;
    _zz_dataOut_payload_0_8732 <= _zz_dataOut_payload_0_8588;
    _zz_dataOut_payload_0_8733 <= _zz_dataOut_payload_0_8589;
    _zz_dataOut_payload_0_8734 <= _zz_dataOut_payload_0_8590;
    _zz_dataOut_payload_0_8735 <= _zz_dataOut_payload_0_8591;
    _zz_dataOut_payload_0_8736 <= _zz_dataOut_payload_0_8704;
    _zz_dataOut_payload_0_8737 <= _zz_dataOut_payload_0_8705;
    _zz_dataOut_payload_0_8738 <= _zz_dataOut_payload_0_8706;
    _zz_dataOut_payload_0_8739 <= _zz_dataOut_payload_0_8707;
    _zz_dataOut_payload_0_8740 <= _zz_dataOut_payload_0_8708;
    _zz_dataOut_payload_0_8741 <= _zz_dataOut_payload_0_8709;
    _zz_dataOut_payload_0_8742 <= _zz_dataOut_payload_0_8710;
    _zz_dataOut_payload_0_8743 <= _zz_dataOut_payload_0_8711;
    _zz_dataOut_payload_0_8744 <= _zz_dataOut_payload_0_8712;
    _zz_dataOut_payload_0_8745 <= _zz_dataOut_payload_0_8713;
    _zz_dataOut_payload_0_8746 <= _zz_dataOut_payload_0_8714;
    _zz_dataOut_payload_0_8747 <= _zz_dataOut_payload_0_8715;
    _zz_dataOut_payload_0_8748 <= _zz_dataOut_payload_0_8716;
    _zz_dataOut_payload_0_8749 <= _zz_dataOut_payload_0_8717;
    _zz_dataOut_payload_0_8750 <= _zz_dataOut_payload_0_8718;
    _zz_dataOut_payload_0_8751 <= _zz_dataOut_payload_0_8719;
    _zz_dataOut_payload_0_8844 <= (_zz_dataOut_payload_0_8842 ? _zz_dataOut_payload_0_8837 : _zz_dataOut_payload_0_8840);
    _zz_dataOut_payload_0_8845 <= (_zz_dataOut_payload_0_8842 ? _zz_dataOut_payload_0_8840 : _zz_dataOut_payload_0_8837);
    _zz_dataOut_payload_0_8846 <= (_zz_dataOut_payload_0_8843 ? _zz_dataOut_payload_0_8838 : _zz_dataOut_payload_0_8841);
    _zz_dataOut_payload_0_8847 <= (_zz_dataOut_payload_0_8843 ? _zz_dataOut_payload_0_8841 : _zz_dataOut_payload_0_8838);
    _zz_dataOut_payload_0_8856 <= (_zz_dataOut_payload_0_8854 ? _zz_dataOut_payload_0_8849 : _zz_dataOut_payload_0_8852);
    _zz_dataOut_payload_0_8857 <= (_zz_dataOut_payload_0_8854 ? _zz_dataOut_payload_0_8852 : _zz_dataOut_payload_0_8849);
    _zz_dataOut_payload_0_8858 <= (_zz_dataOut_payload_0_8855 ? _zz_dataOut_payload_0_8850 : _zz_dataOut_payload_0_8853);
    _zz_dataOut_payload_0_8859 <= (_zz_dataOut_payload_0_8855 ? _zz_dataOut_payload_0_8853 : _zz_dataOut_payload_0_8850);
    _zz_dataOut_payload_0_8860 <= _zz_dataOut_payload_0_8844;
    _zz_dataOut_payload_0_8861 <= _zz_dataOut_payload_0_8845;
    _zz_dataOut_payload_0_8862 <= _zz_dataOut_payload_0_8846;
    _zz_dataOut_payload_0_8863 <= _zz_dataOut_payload_0_8847;
    _zz_dataOut_payload_0_8864 <= _zz_dataOut_payload_0_8856;
    _zz_dataOut_payload_0_8865 <= _zz_dataOut_payload_0_8857;
    _zz_dataOut_payload_0_8866 <= _zz_dataOut_payload_0_8858;
    _zz_dataOut_payload_0_8867 <= _zz_dataOut_payload_0_8859;
    _zz_dataOut_payload_0_8888 <= (_zz_dataOut_payload_0_8886 ? _zz_dataOut_payload_0_8881 : _zz_dataOut_payload_0_8884);
    _zz_dataOut_payload_0_8889 <= (_zz_dataOut_payload_0_8886 ? _zz_dataOut_payload_0_8884 : _zz_dataOut_payload_0_8881);
    _zz_dataOut_payload_0_8890 <= (_zz_dataOut_payload_0_8887 ? _zz_dataOut_payload_0_8882 : _zz_dataOut_payload_0_8885);
    _zz_dataOut_payload_0_8891 <= (_zz_dataOut_payload_0_8887 ? _zz_dataOut_payload_0_8885 : _zz_dataOut_payload_0_8882);
    _zz_dataOut_payload_0_8900 <= (_zz_dataOut_payload_0_8898 ? _zz_dataOut_payload_0_8893 : _zz_dataOut_payload_0_8896);
    _zz_dataOut_payload_0_8901 <= (_zz_dataOut_payload_0_8898 ? _zz_dataOut_payload_0_8896 : _zz_dataOut_payload_0_8893);
    _zz_dataOut_payload_0_8902 <= (_zz_dataOut_payload_0_8899 ? _zz_dataOut_payload_0_8894 : _zz_dataOut_payload_0_8897);
    _zz_dataOut_payload_0_8903 <= (_zz_dataOut_payload_0_8899 ? _zz_dataOut_payload_0_8897 : _zz_dataOut_payload_0_8894);
    _zz_dataOut_payload_0_8904 <= _zz_dataOut_payload_0_8888;
    _zz_dataOut_payload_0_8905 <= _zz_dataOut_payload_0_8889;
    _zz_dataOut_payload_0_8906 <= _zz_dataOut_payload_0_8890;
    _zz_dataOut_payload_0_8907 <= _zz_dataOut_payload_0_8891;
    _zz_dataOut_payload_0_8908 <= _zz_dataOut_payload_0_8900;
    _zz_dataOut_payload_0_8909 <= _zz_dataOut_payload_0_8901;
    _zz_dataOut_payload_0_8910 <= _zz_dataOut_payload_0_8902;
    _zz_dataOut_payload_0_8911 <= _zz_dataOut_payload_0_8903;
    _zz_dataOut_payload_0_8912 <= _zz_dataOut_payload_0_8860;
    _zz_dataOut_payload_0_8913 <= _zz_dataOut_payload_0_8861;
    _zz_dataOut_payload_0_8914 <= _zz_dataOut_payload_0_8862;
    _zz_dataOut_payload_0_8915 <= _zz_dataOut_payload_0_8863;
    _zz_dataOut_payload_0_8916 <= _zz_dataOut_payload_0_8864;
    _zz_dataOut_payload_0_8917 <= _zz_dataOut_payload_0_8865;
    _zz_dataOut_payload_0_8918 <= _zz_dataOut_payload_0_8866;
    _zz_dataOut_payload_0_8919 <= _zz_dataOut_payload_0_8867;
    _zz_dataOut_payload_0_8920 <= _zz_dataOut_payload_0_8904;
    _zz_dataOut_payload_0_8921 <= _zz_dataOut_payload_0_8905;
    _zz_dataOut_payload_0_8922 <= _zz_dataOut_payload_0_8906;
    _zz_dataOut_payload_0_8923 <= _zz_dataOut_payload_0_8907;
    _zz_dataOut_payload_0_8924 <= _zz_dataOut_payload_0_8908;
    _zz_dataOut_payload_0_8925 <= _zz_dataOut_payload_0_8909;
    _zz_dataOut_payload_0_8926 <= _zz_dataOut_payload_0_8910;
    _zz_dataOut_payload_0_8927 <= _zz_dataOut_payload_0_8911;
    _zz_dataOut_payload_0_8972 <= (_zz_dataOut_payload_0_8970 ? _zz_dataOut_payload_0_8965 : _zz_dataOut_payload_0_8968);
    _zz_dataOut_payload_0_8973 <= (_zz_dataOut_payload_0_8970 ? _zz_dataOut_payload_0_8968 : _zz_dataOut_payload_0_8965);
    _zz_dataOut_payload_0_8974 <= (_zz_dataOut_payload_0_8971 ? _zz_dataOut_payload_0_8966 : _zz_dataOut_payload_0_8969);
    _zz_dataOut_payload_0_8975 <= (_zz_dataOut_payload_0_8971 ? _zz_dataOut_payload_0_8969 : _zz_dataOut_payload_0_8966);
    _zz_dataOut_payload_0_8984 <= (_zz_dataOut_payload_0_8982 ? _zz_dataOut_payload_0_8977 : _zz_dataOut_payload_0_8980);
    _zz_dataOut_payload_0_8985 <= (_zz_dataOut_payload_0_8982 ? _zz_dataOut_payload_0_8980 : _zz_dataOut_payload_0_8977);
    _zz_dataOut_payload_0_8986 <= (_zz_dataOut_payload_0_8983 ? _zz_dataOut_payload_0_8978 : _zz_dataOut_payload_0_8981);
    _zz_dataOut_payload_0_8987 <= (_zz_dataOut_payload_0_8983 ? _zz_dataOut_payload_0_8981 : _zz_dataOut_payload_0_8978);
    _zz_dataOut_payload_0_8988 <= _zz_dataOut_payload_0_8972;
    _zz_dataOut_payload_0_8989 <= _zz_dataOut_payload_0_8973;
    _zz_dataOut_payload_0_8990 <= _zz_dataOut_payload_0_8974;
    _zz_dataOut_payload_0_8991 <= _zz_dataOut_payload_0_8975;
    _zz_dataOut_payload_0_8992 <= _zz_dataOut_payload_0_8984;
    _zz_dataOut_payload_0_8993 <= _zz_dataOut_payload_0_8985;
    _zz_dataOut_payload_0_8994 <= _zz_dataOut_payload_0_8986;
    _zz_dataOut_payload_0_8995 <= _zz_dataOut_payload_0_8987;
    _zz_dataOut_payload_0_9016 <= (_zz_dataOut_payload_0_9014 ? _zz_dataOut_payload_0_9009 : _zz_dataOut_payload_0_9012);
    _zz_dataOut_payload_0_9017 <= (_zz_dataOut_payload_0_9014 ? _zz_dataOut_payload_0_9012 : _zz_dataOut_payload_0_9009);
    _zz_dataOut_payload_0_9018 <= (_zz_dataOut_payload_0_9015 ? _zz_dataOut_payload_0_9010 : _zz_dataOut_payload_0_9013);
    _zz_dataOut_payload_0_9019 <= (_zz_dataOut_payload_0_9015 ? _zz_dataOut_payload_0_9013 : _zz_dataOut_payload_0_9010);
    _zz_dataOut_payload_0_9028 <= (_zz_dataOut_payload_0_9026 ? _zz_dataOut_payload_0_9021 : _zz_dataOut_payload_0_9024);
    _zz_dataOut_payload_0_9029 <= (_zz_dataOut_payload_0_9026 ? _zz_dataOut_payload_0_9024 : _zz_dataOut_payload_0_9021);
    _zz_dataOut_payload_0_9030 <= (_zz_dataOut_payload_0_9027 ? _zz_dataOut_payload_0_9022 : _zz_dataOut_payload_0_9025);
    _zz_dataOut_payload_0_9031 <= (_zz_dataOut_payload_0_9027 ? _zz_dataOut_payload_0_9025 : _zz_dataOut_payload_0_9022);
    _zz_dataOut_payload_0_9032 <= _zz_dataOut_payload_0_9016;
    _zz_dataOut_payload_0_9033 <= _zz_dataOut_payload_0_9017;
    _zz_dataOut_payload_0_9034 <= _zz_dataOut_payload_0_9018;
    _zz_dataOut_payload_0_9035 <= _zz_dataOut_payload_0_9019;
    _zz_dataOut_payload_0_9036 <= _zz_dataOut_payload_0_9028;
    _zz_dataOut_payload_0_9037 <= _zz_dataOut_payload_0_9029;
    _zz_dataOut_payload_0_9038 <= _zz_dataOut_payload_0_9030;
    _zz_dataOut_payload_0_9039 <= _zz_dataOut_payload_0_9031;
    _zz_dataOut_payload_0_9040 <= _zz_dataOut_payload_0_8988;
    _zz_dataOut_payload_0_9041 <= _zz_dataOut_payload_0_8989;
    _zz_dataOut_payload_0_9042 <= _zz_dataOut_payload_0_8990;
    _zz_dataOut_payload_0_9043 <= _zz_dataOut_payload_0_8991;
    _zz_dataOut_payload_0_9044 <= _zz_dataOut_payload_0_8992;
    _zz_dataOut_payload_0_9045 <= _zz_dataOut_payload_0_8993;
    _zz_dataOut_payload_0_9046 <= _zz_dataOut_payload_0_8994;
    _zz_dataOut_payload_0_9047 <= _zz_dataOut_payload_0_8995;
    _zz_dataOut_payload_0_9048 <= _zz_dataOut_payload_0_9032;
    _zz_dataOut_payload_0_9049 <= _zz_dataOut_payload_0_9033;
    _zz_dataOut_payload_0_9050 <= _zz_dataOut_payload_0_9034;
    _zz_dataOut_payload_0_9051 <= _zz_dataOut_payload_0_9035;
    _zz_dataOut_payload_0_9052 <= _zz_dataOut_payload_0_9036;
    _zz_dataOut_payload_0_9053 <= _zz_dataOut_payload_0_9037;
    _zz_dataOut_payload_0_9054 <= _zz_dataOut_payload_0_9038;
    _zz_dataOut_payload_0_9055 <= _zz_dataOut_payload_0_9039;
    _zz_dataOut_payload_0_9056 <= _zz_dataOut_payload_0_8912;
    _zz_dataOut_payload_0_9057 <= _zz_dataOut_payload_0_8913;
    _zz_dataOut_payload_0_9058 <= _zz_dataOut_payload_0_8914;
    _zz_dataOut_payload_0_9059 <= _zz_dataOut_payload_0_8915;
    _zz_dataOut_payload_0_9060 <= _zz_dataOut_payload_0_8916;
    _zz_dataOut_payload_0_9061 <= _zz_dataOut_payload_0_8917;
    _zz_dataOut_payload_0_9062 <= _zz_dataOut_payload_0_8918;
    _zz_dataOut_payload_0_9063 <= _zz_dataOut_payload_0_8919;
    _zz_dataOut_payload_0_9064 <= _zz_dataOut_payload_0_8920;
    _zz_dataOut_payload_0_9065 <= _zz_dataOut_payload_0_8921;
    _zz_dataOut_payload_0_9066 <= _zz_dataOut_payload_0_8922;
    _zz_dataOut_payload_0_9067 <= _zz_dataOut_payload_0_8923;
    _zz_dataOut_payload_0_9068 <= _zz_dataOut_payload_0_8924;
    _zz_dataOut_payload_0_9069 <= _zz_dataOut_payload_0_8925;
    _zz_dataOut_payload_0_9070 <= _zz_dataOut_payload_0_8926;
    _zz_dataOut_payload_0_9071 <= _zz_dataOut_payload_0_8927;
    _zz_dataOut_payload_0_9072 <= _zz_dataOut_payload_0_9040;
    _zz_dataOut_payload_0_9073 <= _zz_dataOut_payload_0_9041;
    _zz_dataOut_payload_0_9074 <= _zz_dataOut_payload_0_9042;
    _zz_dataOut_payload_0_9075 <= _zz_dataOut_payload_0_9043;
    _zz_dataOut_payload_0_9076 <= _zz_dataOut_payload_0_9044;
    _zz_dataOut_payload_0_9077 <= _zz_dataOut_payload_0_9045;
    _zz_dataOut_payload_0_9078 <= _zz_dataOut_payload_0_9046;
    _zz_dataOut_payload_0_9079 <= _zz_dataOut_payload_0_9047;
    _zz_dataOut_payload_0_9080 <= _zz_dataOut_payload_0_9048;
    _zz_dataOut_payload_0_9081 <= _zz_dataOut_payload_0_9049;
    _zz_dataOut_payload_0_9082 <= _zz_dataOut_payload_0_9050;
    _zz_dataOut_payload_0_9083 <= _zz_dataOut_payload_0_9051;
    _zz_dataOut_payload_0_9084 <= _zz_dataOut_payload_0_9052;
    _zz_dataOut_payload_0_9085 <= _zz_dataOut_payload_0_9053;
    _zz_dataOut_payload_0_9086 <= _zz_dataOut_payload_0_9054;
    _zz_dataOut_payload_0_9087 <= _zz_dataOut_payload_0_9055;
    _zz_dataOut_payload_0_9088 <= _zz_dataOut_payload_0_8720;
    _zz_dataOut_payload_0_9089 <= _zz_dataOut_payload_0_8721;
    _zz_dataOut_payload_0_9090 <= _zz_dataOut_payload_0_8722;
    _zz_dataOut_payload_0_9091 <= _zz_dataOut_payload_0_8723;
    _zz_dataOut_payload_0_9092 <= _zz_dataOut_payload_0_8724;
    _zz_dataOut_payload_0_9093 <= _zz_dataOut_payload_0_8725;
    _zz_dataOut_payload_0_9094 <= _zz_dataOut_payload_0_8726;
    _zz_dataOut_payload_0_9095 <= _zz_dataOut_payload_0_8727;
    _zz_dataOut_payload_0_9096 <= _zz_dataOut_payload_0_8728;
    _zz_dataOut_payload_0_9097 <= _zz_dataOut_payload_0_8729;
    _zz_dataOut_payload_0_9098 <= _zz_dataOut_payload_0_8730;
    _zz_dataOut_payload_0_9099 <= _zz_dataOut_payload_0_8731;
    _zz_dataOut_payload_0_9100 <= _zz_dataOut_payload_0_8732;
    _zz_dataOut_payload_0_9101 <= _zz_dataOut_payload_0_8733;
    _zz_dataOut_payload_0_9102 <= _zz_dataOut_payload_0_8734;
    _zz_dataOut_payload_0_9103 <= _zz_dataOut_payload_0_8735;
    _zz_dataOut_payload_0_9104 <= _zz_dataOut_payload_0_8736;
    _zz_dataOut_payload_0_9105 <= _zz_dataOut_payload_0_8737;
    _zz_dataOut_payload_0_9106 <= _zz_dataOut_payload_0_8738;
    _zz_dataOut_payload_0_9107 <= _zz_dataOut_payload_0_8739;
    _zz_dataOut_payload_0_9108 <= _zz_dataOut_payload_0_8740;
    _zz_dataOut_payload_0_9109 <= _zz_dataOut_payload_0_8741;
    _zz_dataOut_payload_0_9110 <= _zz_dataOut_payload_0_8742;
    _zz_dataOut_payload_0_9111 <= _zz_dataOut_payload_0_8743;
    _zz_dataOut_payload_0_9112 <= _zz_dataOut_payload_0_8744;
    _zz_dataOut_payload_0_9113 <= _zz_dataOut_payload_0_8745;
    _zz_dataOut_payload_0_9114 <= _zz_dataOut_payload_0_8746;
    _zz_dataOut_payload_0_9115 <= _zz_dataOut_payload_0_8747;
    _zz_dataOut_payload_0_9116 <= _zz_dataOut_payload_0_8748;
    _zz_dataOut_payload_0_9117 <= _zz_dataOut_payload_0_8749;
    _zz_dataOut_payload_0_9118 <= _zz_dataOut_payload_0_8750;
    _zz_dataOut_payload_0_9119 <= _zz_dataOut_payload_0_8751;
    _zz_dataOut_payload_0_9120 <= _zz_dataOut_payload_0_9056;
    _zz_dataOut_payload_0_9121 <= _zz_dataOut_payload_0_9057;
    _zz_dataOut_payload_0_9122 <= _zz_dataOut_payload_0_9058;
    _zz_dataOut_payload_0_9123 <= _zz_dataOut_payload_0_9059;
    _zz_dataOut_payload_0_9124 <= _zz_dataOut_payload_0_9060;
    _zz_dataOut_payload_0_9125 <= _zz_dataOut_payload_0_9061;
    _zz_dataOut_payload_0_9126 <= _zz_dataOut_payload_0_9062;
    _zz_dataOut_payload_0_9127 <= _zz_dataOut_payload_0_9063;
    _zz_dataOut_payload_0_9128 <= _zz_dataOut_payload_0_9064;
    _zz_dataOut_payload_0_9129 <= _zz_dataOut_payload_0_9065;
    _zz_dataOut_payload_0_9130 <= _zz_dataOut_payload_0_9066;
    _zz_dataOut_payload_0_9131 <= _zz_dataOut_payload_0_9067;
    _zz_dataOut_payload_0_9132 <= _zz_dataOut_payload_0_9068;
    _zz_dataOut_payload_0_9133 <= _zz_dataOut_payload_0_9069;
    _zz_dataOut_payload_0_9134 <= _zz_dataOut_payload_0_9070;
    _zz_dataOut_payload_0_9135 <= _zz_dataOut_payload_0_9071;
    _zz_dataOut_payload_0_9136 <= _zz_dataOut_payload_0_9072;
    _zz_dataOut_payload_0_9137 <= _zz_dataOut_payload_0_9073;
    _zz_dataOut_payload_0_9138 <= _zz_dataOut_payload_0_9074;
    _zz_dataOut_payload_0_9139 <= _zz_dataOut_payload_0_9075;
    _zz_dataOut_payload_0_9140 <= _zz_dataOut_payload_0_9076;
    _zz_dataOut_payload_0_9141 <= _zz_dataOut_payload_0_9077;
    _zz_dataOut_payload_0_9142 <= _zz_dataOut_payload_0_9078;
    _zz_dataOut_payload_0_9143 <= _zz_dataOut_payload_0_9079;
    _zz_dataOut_payload_0_9144 <= _zz_dataOut_payload_0_9080;
    _zz_dataOut_payload_0_9145 <= _zz_dataOut_payload_0_9081;
    _zz_dataOut_payload_0_9146 <= _zz_dataOut_payload_0_9082;
    _zz_dataOut_payload_0_9147 <= _zz_dataOut_payload_0_9083;
    _zz_dataOut_payload_0_9148 <= _zz_dataOut_payload_0_9084;
    _zz_dataOut_payload_0_9149 <= _zz_dataOut_payload_0_9085;
    _zz_dataOut_payload_0_9150 <= _zz_dataOut_payload_0_9086;
    _zz_dataOut_payload_0_9151 <= _zz_dataOut_payload_0_9087;
    _zz_dataOut_payload_0_9340 <= (_zz_dataOut_payload_0_9338 ? _zz_dataOut_payload_0_9333 : _zz_dataOut_payload_0_9336);
    _zz_dataOut_payload_0_9341 <= (_zz_dataOut_payload_0_9338 ? _zz_dataOut_payload_0_9336 : _zz_dataOut_payload_0_9333);
    _zz_dataOut_payload_0_9342 <= (_zz_dataOut_payload_0_9339 ? _zz_dataOut_payload_0_9334 : _zz_dataOut_payload_0_9337);
    _zz_dataOut_payload_0_9343 <= (_zz_dataOut_payload_0_9339 ? _zz_dataOut_payload_0_9337 : _zz_dataOut_payload_0_9334);
    _zz_dataOut_payload_0_9352 <= (_zz_dataOut_payload_0_9350 ? _zz_dataOut_payload_0_9345 : _zz_dataOut_payload_0_9348);
    _zz_dataOut_payload_0_9353 <= (_zz_dataOut_payload_0_9350 ? _zz_dataOut_payload_0_9348 : _zz_dataOut_payload_0_9345);
    _zz_dataOut_payload_0_9354 <= (_zz_dataOut_payload_0_9351 ? _zz_dataOut_payload_0_9346 : _zz_dataOut_payload_0_9349);
    _zz_dataOut_payload_0_9355 <= (_zz_dataOut_payload_0_9351 ? _zz_dataOut_payload_0_9349 : _zz_dataOut_payload_0_9346);
    _zz_dataOut_payload_0_9356 <= _zz_dataOut_payload_0_9340;
    _zz_dataOut_payload_0_9357 <= _zz_dataOut_payload_0_9341;
    _zz_dataOut_payload_0_9358 <= _zz_dataOut_payload_0_9342;
    _zz_dataOut_payload_0_9359 <= _zz_dataOut_payload_0_9343;
    _zz_dataOut_payload_0_9360 <= _zz_dataOut_payload_0_9352;
    _zz_dataOut_payload_0_9361 <= _zz_dataOut_payload_0_9353;
    _zz_dataOut_payload_0_9362 <= _zz_dataOut_payload_0_9354;
    _zz_dataOut_payload_0_9363 <= _zz_dataOut_payload_0_9355;
    _zz_dataOut_payload_0_9384 <= (_zz_dataOut_payload_0_9382 ? _zz_dataOut_payload_0_9377 : _zz_dataOut_payload_0_9380);
    _zz_dataOut_payload_0_9385 <= (_zz_dataOut_payload_0_9382 ? _zz_dataOut_payload_0_9380 : _zz_dataOut_payload_0_9377);
    _zz_dataOut_payload_0_9386 <= (_zz_dataOut_payload_0_9383 ? _zz_dataOut_payload_0_9378 : _zz_dataOut_payload_0_9381);
    _zz_dataOut_payload_0_9387 <= (_zz_dataOut_payload_0_9383 ? _zz_dataOut_payload_0_9381 : _zz_dataOut_payload_0_9378);
    _zz_dataOut_payload_0_9396 <= (_zz_dataOut_payload_0_9394 ? _zz_dataOut_payload_0_9389 : _zz_dataOut_payload_0_9392);
    _zz_dataOut_payload_0_9397 <= (_zz_dataOut_payload_0_9394 ? _zz_dataOut_payload_0_9392 : _zz_dataOut_payload_0_9389);
    _zz_dataOut_payload_0_9398 <= (_zz_dataOut_payload_0_9395 ? _zz_dataOut_payload_0_9390 : _zz_dataOut_payload_0_9393);
    _zz_dataOut_payload_0_9399 <= (_zz_dataOut_payload_0_9395 ? _zz_dataOut_payload_0_9393 : _zz_dataOut_payload_0_9390);
    _zz_dataOut_payload_0_9400 <= _zz_dataOut_payload_0_9384;
    _zz_dataOut_payload_0_9401 <= _zz_dataOut_payload_0_9385;
    _zz_dataOut_payload_0_9402 <= _zz_dataOut_payload_0_9386;
    _zz_dataOut_payload_0_9403 <= _zz_dataOut_payload_0_9387;
    _zz_dataOut_payload_0_9404 <= _zz_dataOut_payload_0_9396;
    _zz_dataOut_payload_0_9405 <= _zz_dataOut_payload_0_9397;
    _zz_dataOut_payload_0_9406 <= _zz_dataOut_payload_0_9398;
    _zz_dataOut_payload_0_9407 <= _zz_dataOut_payload_0_9399;
    _zz_dataOut_payload_0_9408 <= _zz_dataOut_payload_0_9356;
    _zz_dataOut_payload_0_9409 <= _zz_dataOut_payload_0_9357;
    _zz_dataOut_payload_0_9410 <= _zz_dataOut_payload_0_9358;
    _zz_dataOut_payload_0_9411 <= _zz_dataOut_payload_0_9359;
    _zz_dataOut_payload_0_9412 <= _zz_dataOut_payload_0_9360;
    _zz_dataOut_payload_0_9413 <= _zz_dataOut_payload_0_9361;
    _zz_dataOut_payload_0_9414 <= _zz_dataOut_payload_0_9362;
    _zz_dataOut_payload_0_9415 <= _zz_dataOut_payload_0_9363;
    _zz_dataOut_payload_0_9416 <= _zz_dataOut_payload_0_9400;
    _zz_dataOut_payload_0_9417 <= _zz_dataOut_payload_0_9401;
    _zz_dataOut_payload_0_9418 <= _zz_dataOut_payload_0_9402;
    _zz_dataOut_payload_0_9419 <= _zz_dataOut_payload_0_9403;
    _zz_dataOut_payload_0_9420 <= _zz_dataOut_payload_0_9404;
    _zz_dataOut_payload_0_9421 <= _zz_dataOut_payload_0_9405;
    _zz_dataOut_payload_0_9422 <= _zz_dataOut_payload_0_9406;
    _zz_dataOut_payload_0_9423 <= _zz_dataOut_payload_0_9407;
    _zz_dataOut_payload_0_9468 <= (_zz_dataOut_payload_0_9466 ? _zz_dataOut_payload_0_9461 : _zz_dataOut_payload_0_9464);
    _zz_dataOut_payload_0_9469 <= (_zz_dataOut_payload_0_9466 ? _zz_dataOut_payload_0_9464 : _zz_dataOut_payload_0_9461);
    _zz_dataOut_payload_0_9470 <= (_zz_dataOut_payload_0_9467 ? _zz_dataOut_payload_0_9462 : _zz_dataOut_payload_0_9465);
    _zz_dataOut_payload_0_9471 <= (_zz_dataOut_payload_0_9467 ? _zz_dataOut_payload_0_9465 : _zz_dataOut_payload_0_9462);
    _zz_dataOut_payload_0_9480 <= (_zz_dataOut_payload_0_9478 ? _zz_dataOut_payload_0_9473 : _zz_dataOut_payload_0_9476);
    _zz_dataOut_payload_0_9481 <= (_zz_dataOut_payload_0_9478 ? _zz_dataOut_payload_0_9476 : _zz_dataOut_payload_0_9473);
    _zz_dataOut_payload_0_9482 <= (_zz_dataOut_payload_0_9479 ? _zz_dataOut_payload_0_9474 : _zz_dataOut_payload_0_9477);
    _zz_dataOut_payload_0_9483 <= (_zz_dataOut_payload_0_9479 ? _zz_dataOut_payload_0_9477 : _zz_dataOut_payload_0_9474);
    _zz_dataOut_payload_0_9484 <= _zz_dataOut_payload_0_9468;
    _zz_dataOut_payload_0_9485 <= _zz_dataOut_payload_0_9469;
    _zz_dataOut_payload_0_9486 <= _zz_dataOut_payload_0_9470;
    _zz_dataOut_payload_0_9487 <= _zz_dataOut_payload_0_9471;
    _zz_dataOut_payload_0_9488 <= _zz_dataOut_payload_0_9480;
    _zz_dataOut_payload_0_9489 <= _zz_dataOut_payload_0_9481;
    _zz_dataOut_payload_0_9490 <= _zz_dataOut_payload_0_9482;
    _zz_dataOut_payload_0_9491 <= _zz_dataOut_payload_0_9483;
    _zz_dataOut_payload_0_9512 <= (_zz_dataOut_payload_0_9510 ? _zz_dataOut_payload_0_9505 : _zz_dataOut_payload_0_9508);
    _zz_dataOut_payload_0_9513 <= (_zz_dataOut_payload_0_9510 ? _zz_dataOut_payload_0_9508 : _zz_dataOut_payload_0_9505);
    _zz_dataOut_payload_0_9514 <= (_zz_dataOut_payload_0_9511 ? _zz_dataOut_payload_0_9506 : _zz_dataOut_payload_0_9509);
    _zz_dataOut_payload_0_9515 <= (_zz_dataOut_payload_0_9511 ? _zz_dataOut_payload_0_9509 : _zz_dataOut_payload_0_9506);
    _zz_dataOut_payload_0_9524 <= (_zz_dataOut_payload_0_9522 ? _zz_dataOut_payload_0_9517 : _zz_dataOut_payload_0_9520);
    _zz_dataOut_payload_0_9525 <= (_zz_dataOut_payload_0_9522 ? _zz_dataOut_payload_0_9520 : _zz_dataOut_payload_0_9517);
    _zz_dataOut_payload_0_9526 <= (_zz_dataOut_payload_0_9523 ? _zz_dataOut_payload_0_9518 : _zz_dataOut_payload_0_9521);
    _zz_dataOut_payload_0_9527 <= (_zz_dataOut_payload_0_9523 ? _zz_dataOut_payload_0_9521 : _zz_dataOut_payload_0_9518);
    _zz_dataOut_payload_0_9528 <= _zz_dataOut_payload_0_9512;
    _zz_dataOut_payload_0_9529 <= _zz_dataOut_payload_0_9513;
    _zz_dataOut_payload_0_9530 <= _zz_dataOut_payload_0_9514;
    _zz_dataOut_payload_0_9531 <= _zz_dataOut_payload_0_9515;
    _zz_dataOut_payload_0_9532 <= _zz_dataOut_payload_0_9524;
    _zz_dataOut_payload_0_9533 <= _zz_dataOut_payload_0_9525;
    _zz_dataOut_payload_0_9534 <= _zz_dataOut_payload_0_9526;
    _zz_dataOut_payload_0_9535 <= _zz_dataOut_payload_0_9527;
    _zz_dataOut_payload_0_9536 <= _zz_dataOut_payload_0_9484;
    _zz_dataOut_payload_0_9537 <= _zz_dataOut_payload_0_9485;
    _zz_dataOut_payload_0_9538 <= _zz_dataOut_payload_0_9486;
    _zz_dataOut_payload_0_9539 <= _zz_dataOut_payload_0_9487;
    _zz_dataOut_payload_0_9540 <= _zz_dataOut_payload_0_9488;
    _zz_dataOut_payload_0_9541 <= _zz_dataOut_payload_0_9489;
    _zz_dataOut_payload_0_9542 <= _zz_dataOut_payload_0_9490;
    _zz_dataOut_payload_0_9543 <= _zz_dataOut_payload_0_9491;
    _zz_dataOut_payload_0_9544 <= _zz_dataOut_payload_0_9528;
    _zz_dataOut_payload_0_9545 <= _zz_dataOut_payload_0_9529;
    _zz_dataOut_payload_0_9546 <= _zz_dataOut_payload_0_9530;
    _zz_dataOut_payload_0_9547 <= _zz_dataOut_payload_0_9531;
    _zz_dataOut_payload_0_9548 <= _zz_dataOut_payload_0_9532;
    _zz_dataOut_payload_0_9549 <= _zz_dataOut_payload_0_9533;
    _zz_dataOut_payload_0_9550 <= _zz_dataOut_payload_0_9534;
    _zz_dataOut_payload_0_9551 <= _zz_dataOut_payload_0_9535;
    _zz_dataOut_payload_0_9552 <= _zz_dataOut_payload_0_9408;
    _zz_dataOut_payload_0_9553 <= _zz_dataOut_payload_0_9409;
    _zz_dataOut_payload_0_9554 <= _zz_dataOut_payload_0_9410;
    _zz_dataOut_payload_0_9555 <= _zz_dataOut_payload_0_9411;
    _zz_dataOut_payload_0_9556 <= _zz_dataOut_payload_0_9412;
    _zz_dataOut_payload_0_9557 <= _zz_dataOut_payload_0_9413;
    _zz_dataOut_payload_0_9558 <= _zz_dataOut_payload_0_9414;
    _zz_dataOut_payload_0_9559 <= _zz_dataOut_payload_0_9415;
    _zz_dataOut_payload_0_9560 <= _zz_dataOut_payload_0_9416;
    _zz_dataOut_payload_0_9561 <= _zz_dataOut_payload_0_9417;
    _zz_dataOut_payload_0_9562 <= _zz_dataOut_payload_0_9418;
    _zz_dataOut_payload_0_9563 <= _zz_dataOut_payload_0_9419;
    _zz_dataOut_payload_0_9564 <= _zz_dataOut_payload_0_9420;
    _zz_dataOut_payload_0_9565 <= _zz_dataOut_payload_0_9421;
    _zz_dataOut_payload_0_9566 <= _zz_dataOut_payload_0_9422;
    _zz_dataOut_payload_0_9567 <= _zz_dataOut_payload_0_9423;
    _zz_dataOut_payload_0_9568 <= _zz_dataOut_payload_0_9536;
    _zz_dataOut_payload_0_9569 <= _zz_dataOut_payload_0_9537;
    _zz_dataOut_payload_0_9570 <= _zz_dataOut_payload_0_9538;
    _zz_dataOut_payload_0_9571 <= _zz_dataOut_payload_0_9539;
    _zz_dataOut_payload_0_9572 <= _zz_dataOut_payload_0_9540;
    _zz_dataOut_payload_0_9573 <= _zz_dataOut_payload_0_9541;
    _zz_dataOut_payload_0_9574 <= _zz_dataOut_payload_0_9542;
    _zz_dataOut_payload_0_9575 <= _zz_dataOut_payload_0_9543;
    _zz_dataOut_payload_0_9576 <= _zz_dataOut_payload_0_9544;
    _zz_dataOut_payload_0_9577 <= _zz_dataOut_payload_0_9545;
    _zz_dataOut_payload_0_9578 <= _zz_dataOut_payload_0_9546;
    _zz_dataOut_payload_0_9579 <= _zz_dataOut_payload_0_9547;
    _zz_dataOut_payload_0_9580 <= _zz_dataOut_payload_0_9548;
    _zz_dataOut_payload_0_9581 <= _zz_dataOut_payload_0_9549;
    _zz_dataOut_payload_0_9582 <= _zz_dataOut_payload_0_9550;
    _zz_dataOut_payload_0_9583 <= _zz_dataOut_payload_0_9551;
    _zz_dataOut_payload_0_9676 <= (_zz_dataOut_payload_0_9674 ? _zz_dataOut_payload_0_9669 : _zz_dataOut_payload_0_9672);
    _zz_dataOut_payload_0_9677 <= (_zz_dataOut_payload_0_9674 ? _zz_dataOut_payload_0_9672 : _zz_dataOut_payload_0_9669);
    _zz_dataOut_payload_0_9678 <= (_zz_dataOut_payload_0_9675 ? _zz_dataOut_payload_0_9670 : _zz_dataOut_payload_0_9673);
    _zz_dataOut_payload_0_9679 <= (_zz_dataOut_payload_0_9675 ? _zz_dataOut_payload_0_9673 : _zz_dataOut_payload_0_9670);
    _zz_dataOut_payload_0_9688 <= (_zz_dataOut_payload_0_9686 ? _zz_dataOut_payload_0_9681 : _zz_dataOut_payload_0_9684);
    _zz_dataOut_payload_0_9689 <= (_zz_dataOut_payload_0_9686 ? _zz_dataOut_payload_0_9684 : _zz_dataOut_payload_0_9681);
    _zz_dataOut_payload_0_9690 <= (_zz_dataOut_payload_0_9687 ? _zz_dataOut_payload_0_9682 : _zz_dataOut_payload_0_9685);
    _zz_dataOut_payload_0_9691 <= (_zz_dataOut_payload_0_9687 ? _zz_dataOut_payload_0_9685 : _zz_dataOut_payload_0_9682);
    _zz_dataOut_payload_0_9692 <= _zz_dataOut_payload_0_9676;
    _zz_dataOut_payload_0_9693 <= _zz_dataOut_payload_0_9677;
    _zz_dataOut_payload_0_9694 <= _zz_dataOut_payload_0_9678;
    _zz_dataOut_payload_0_9695 <= _zz_dataOut_payload_0_9679;
    _zz_dataOut_payload_0_9696 <= _zz_dataOut_payload_0_9688;
    _zz_dataOut_payload_0_9697 <= _zz_dataOut_payload_0_9689;
    _zz_dataOut_payload_0_9698 <= _zz_dataOut_payload_0_9690;
    _zz_dataOut_payload_0_9699 <= _zz_dataOut_payload_0_9691;
    _zz_dataOut_payload_0_9720 <= (_zz_dataOut_payload_0_9718 ? _zz_dataOut_payload_0_9713 : _zz_dataOut_payload_0_9716);
    _zz_dataOut_payload_0_9721 <= (_zz_dataOut_payload_0_9718 ? _zz_dataOut_payload_0_9716 : _zz_dataOut_payload_0_9713);
    _zz_dataOut_payload_0_9722 <= (_zz_dataOut_payload_0_9719 ? _zz_dataOut_payload_0_9714 : _zz_dataOut_payload_0_9717);
    _zz_dataOut_payload_0_9723 <= (_zz_dataOut_payload_0_9719 ? _zz_dataOut_payload_0_9717 : _zz_dataOut_payload_0_9714);
    _zz_dataOut_payload_0_9732 <= (_zz_dataOut_payload_0_9730 ? _zz_dataOut_payload_0_9725 : _zz_dataOut_payload_0_9728);
    _zz_dataOut_payload_0_9733 <= (_zz_dataOut_payload_0_9730 ? _zz_dataOut_payload_0_9728 : _zz_dataOut_payload_0_9725);
    _zz_dataOut_payload_0_9734 <= (_zz_dataOut_payload_0_9731 ? _zz_dataOut_payload_0_9726 : _zz_dataOut_payload_0_9729);
    _zz_dataOut_payload_0_9735 <= (_zz_dataOut_payload_0_9731 ? _zz_dataOut_payload_0_9729 : _zz_dataOut_payload_0_9726);
    _zz_dataOut_payload_0_9736 <= _zz_dataOut_payload_0_9720;
    _zz_dataOut_payload_0_9737 <= _zz_dataOut_payload_0_9721;
    _zz_dataOut_payload_0_9738 <= _zz_dataOut_payload_0_9722;
    _zz_dataOut_payload_0_9739 <= _zz_dataOut_payload_0_9723;
    _zz_dataOut_payload_0_9740 <= _zz_dataOut_payload_0_9732;
    _zz_dataOut_payload_0_9741 <= _zz_dataOut_payload_0_9733;
    _zz_dataOut_payload_0_9742 <= _zz_dataOut_payload_0_9734;
    _zz_dataOut_payload_0_9743 <= _zz_dataOut_payload_0_9735;
    _zz_dataOut_payload_0_9744 <= _zz_dataOut_payload_0_9692;
    _zz_dataOut_payload_0_9745 <= _zz_dataOut_payload_0_9693;
    _zz_dataOut_payload_0_9746 <= _zz_dataOut_payload_0_9694;
    _zz_dataOut_payload_0_9747 <= _zz_dataOut_payload_0_9695;
    _zz_dataOut_payload_0_9748 <= _zz_dataOut_payload_0_9696;
    _zz_dataOut_payload_0_9749 <= _zz_dataOut_payload_0_9697;
    _zz_dataOut_payload_0_9750 <= _zz_dataOut_payload_0_9698;
    _zz_dataOut_payload_0_9751 <= _zz_dataOut_payload_0_9699;
    _zz_dataOut_payload_0_9752 <= _zz_dataOut_payload_0_9736;
    _zz_dataOut_payload_0_9753 <= _zz_dataOut_payload_0_9737;
    _zz_dataOut_payload_0_9754 <= _zz_dataOut_payload_0_9738;
    _zz_dataOut_payload_0_9755 <= _zz_dataOut_payload_0_9739;
    _zz_dataOut_payload_0_9756 <= _zz_dataOut_payload_0_9740;
    _zz_dataOut_payload_0_9757 <= _zz_dataOut_payload_0_9741;
    _zz_dataOut_payload_0_9758 <= _zz_dataOut_payload_0_9742;
    _zz_dataOut_payload_0_9759 <= _zz_dataOut_payload_0_9743;
    _zz_dataOut_payload_0_9804 <= (_zz_dataOut_payload_0_9802 ? _zz_dataOut_payload_0_9797 : _zz_dataOut_payload_0_9800);
    _zz_dataOut_payload_0_9805 <= (_zz_dataOut_payload_0_9802 ? _zz_dataOut_payload_0_9800 : _zz_dataOut_payload_0_9797);
    _zz_dataOut_payload_0_9806 <= (_zz_dataOut_payload_0_9803 ? _zz_dataOut_payload_0_9798 : _zz_dataOut_payload_0_9801);
    _zz_dataOut_payload_0_9807 <= (_zz_dataOut_payload_0_9803 ? _zz_dataOut_payload_0_9801 : _zz_dataOut_payload_0_9798);
    _zz_dataOut_payload_0_9816 <= (_zz_dataOut_payload_0_9814 ? _zz_dataOut_payload_0_9809 : _zz_dataOut_payload_0_9812);
    _zz_dataOut_payload_0_9817 <= (_zz_dataOut_payload_0_9814 ? _zz_dataOut_payload_0_9812 : _zz_dataOut_payload_0_9809);
    _zz_dataOut_payload_0_9818 <= (_zz_dataOut_payload_0_9815 ? _zz_dataOut_payload_0_9810 : _zz_dataOut_payload_0_9813);
    _zz_dataOut_payload_0_9819 <= (_zz_dataOut_payload_0_9815 ? _zz_dataOut_payload_0_9813 : _zz_dataOut_payload_0_9810);
    _zz_dataOut_payload_0_9820 <= _zz_dataOut_payload_0_9804;
    _zz_dataOut_payload_0_9821 <= _zz_dataOut_payload_0_9805;
    _zz_dataOut_payload_0_9822 <= _zz_dataOut_payload_0_9806;
    _zz_dataOut_payload_0_9823 <= _zz_dataOut_payload_0_9807;
    _zz_dataOut_payload_0_9824 <= _zz_dataOut_payload_0_9816;
    _zz_dataOut_payload_0_9825 <= _zz_dataOut_payload_0_9817;
    _zz_dataOut_payload_0_9826 <= _zz_dataOut_payload_0_9818;
    _zz_dataOut_payload_0_9827 <= _zz_dataOut_payload_0_9819;
    _zz_dataOut_payload_0_9848 <= (_zz_dataOut_payload_0_9846 ? _zz_dataOut_payload_0_9841 : _zz_dataOut_payload_0_9844);
    _zz_dataOut_payload_0_9849 <= (_zz_dataOut_payload_0_9846 ? _zz_dataOut_payload_0_9844 : _zz_dataOut_payload_0_9841);
    _zz_dataOut_payload_0_9850 <= (_zz_dataOut_payload_0_9847 ? _zz_dataOut_payload_0_9842 : _zz_dataOut_payload_0_9845);
    _zz_dataOut_payload_0_9851 <= (_zz_dataOut_payload_0_9847 ? _zz_dataOut_payload_0_9845 : _zz_dataOut_payload_0_9842);
    _zz_dataOut_payload_0_9860 <= (_zz_dataOut_payload_0_9858 ? _zz_dataOut_payload_0_9853 : _zz_dataOut_payload_0_9856);
    _zz_dataOut_payload_0_9861 <= (_zz_dataOut_payload_0_9858 ? _zz_dataOut_payload_0_9856 : _zz_dataOut_payload_0_9853);
    _zz_dataOut_payload_0_9862 <= (_zz_dataOut_payload_0_9859 ? _zz_dataOut_payload_0_9854 : _zz_dataOut_payload_0_9857);
    _zz_dataOut_payload_0_9863 <= (_zz_dataOut_payload_0_9859 ? _zz_dataOut_payload_0_9857 : _zz_dataOut_payload_0_9854);
    _zz_dataOut_payload_0_9864 <= _zz_dataOut_payload_0_9848;
    _zz_dataOut_payload_0_9865 <= _zz_dataOut_payload_0_9849;
    _zz_dataOut_payload_0_9866 <= _zz_dataOut_payload_0_9850;
    _zz_dataOut_payload_0_9867 <= _zz_dataOut_payload_0_9851;
    _zz_dataOut_payload_0_9868 <= _zz_dataOut_payload_0_9860;
    _zz_dataOut_payload_0_9869 <= _zz_dataOut_payload_0_9861;
    _zz_dataOut_payload_0_9870 <= _zz_dataOut_payload_0_9862;
    _zz_dataOut_payload_0_9871 <= _zz_dataOut_payload_0_9863;
    _zz_dataOut_payload_0_9872 <= _zz_dataOut_payload_0_9820;
    _zz_dataOut_payload_0_9873 <= _zz_dataOut_payload_0_9821;
    _zz_dataOut_payload_0_9874 <= _zz_dataOut_payload_0_9822;
    _zz_dataOut_payload_0_9875 <= _zz_dataOut_payload_0_9823;
    _zz_dataOut_payload_0_9876 <= _zz_dataOut_payload_0_9824;
    _zz_dataOut_payload_0_9877 <= _zz_dataOut_payload_0_9825;
    _zz_dataOut_payload_0_9878 <= _zz_dataOut_payload_0_9826;
    _zz_dataOut_payload_0_9879 <= _zz_dataOut_payload_0_9827;
    _zz_dataOut_payload_0_9880 <= _zz_dataOut_payload_0_9864;
    _zz_dataOut_payload_0_9881 <= _zz_dataOut_payload_0_9865;
    _zz_dataOut_payload_0_9882 <= _zz_dataOut_payload_0_9866;
    _zz_dataOut_payload_0_9883 <= _zz_dataOut_payload_0_9867;
    _zz_dataOut_payload_0_9884 <= _zz_dataOut_payload_0_9868;
    _zz_dataOut_payload_0_9885 <= _zz_dataOut_payload_0_9869;
    _zz_dataOut_payload_0_9886 <= _zz_dataOut_payload_0_9870;
    _zz_dataOut_payload_0_9887 <= _zz_dataOut_payload_0_9871;
    _zz_dataOut_payload_0_9888 <= _zz_dataOut_payload_0_9744;
    _zz_dataOut_payload_0_9889 <= _zz_dataOut_payload_0_9745;
    _zz_dataOut_payload_0_9890 <= _zz_dataOut_payload_0_9746;
    _zz_dataOut_payload_0_9891 <= _zz_dataOut_payload_0_9747;
    _zz_dataOut_payload_0_9892 <= _zz_dataOut_payload_0_9748;
    _zz_dataOut_payload_0_9893 <= _zz_dataOut_payload_0_9749;
    _zz_dataOut_payload_0_9894 <= _zz_dataOut_payload_0_9750;
    _zz_dataOut_payload_0_9895 <= _zz_dataOut_payload_0_9751;
    _zz_dataOut_payload_0_9896 <= _zz_dataOut_payload_0_9752;
    _zz_dataOut_payload_0_9897 <= _zz_dataOut_payload_0_9753;
    _zz_dataOut_payload_0_9898 <= _zz_dataOut_payload_0_9754;
    _zz_dataOut_payload_0_9899 <= _zz_dataOut_payload_0_9755;
    _zz_dataOut_payload_0_9900 <= _zz_dataOut_payload_0_9756;
    _zz_dataOut_payload_0_9901 <= _zz_dataOut_payload_0_9757;
    _zz_dataOut_payload_0_9902 <= _zz_dataOut_payload_0_9758;
    _zz_dataOut_payload_0_9903 <= _zz_dataOut_payload_0_9759;
    _zz_dataOut_payload_0_9904 <= _zz_dataOut_payload_0_9872;
    _zz_dataOut_payload_0_9905 <= _zz_dataOut_payload_0_9873;
    _zz_dataOut_payload_0_9906 <= _zz_dataOut_payload_0_9874;
    _zz_dataOut_payload_0_9907 <= _zz_dataOut_payload_0_9875;
    _zz_dataOut_payload_0_9908 <= _zz_dataOut_payload_0_9876;
    _zz_dataOut_payload_0_9909 <= _zz_dataOut_payload_0_9877;
    _zz_dataOut_payload_0_9910 <= _zz_dataOut_payload_0_9878;
    _zz_dataOut_payload_0_9911 <= _zz_dataOut_payload_0_9879;
    _zz_dataOut_payload_0_9912 <= _zz_dataOut_payload_0_9880;
    _zz_dataOut_payload_0_9913 <= _zz_dataOut_payload_0_9881;
    _zz_dataOut_payload_0_9914 <= _zz_dataOut_payload_0_9882;
    _zz_dataOut_payload_0_9915 <= _zz_dataOut_payload_0_9883;
    _zz_dataOut_payload_0_9916 <= _zz_dataOut_payload_0_9884;
    _zz_dataOut_payload_0_9917 <= _zz_dataOut_payload_0_9885;
    _zz_dataOut_payload_0_9918 <= _zz_dataOut_payload_0_9886;
    _zz_dataOut_payload_0_9919 <= _zz_dataOut_payload_0_9887;
    _zz_dataOut_payload_0_9920 <= _zz_dataOut_payload_0_9552;
    _zz_dataOut_payload_0_9921 <= _zz_dataOut_payload_0_9553;
    _zz_dataOut_payload_0_9922 <= _zz_dataOut_payload_0_9554;
    _zz_dataOut_payload_0_9923 <= _zz_dataOut_payload_0_9555;
    _zz_dataOut_payload_0_9924 <= _zz_dataOut_payload_0_9556;
    _zz_dataOut_payload_0_9925 <= _zz_dataOut_payload_0_9557;
    _zz_dataOut_payload_0_9926 <= _zz_dataOut_payload_0_9558;
    _zz_dataOut_payload_0_9927 <= _zz_dataOut_payload_0_9559;
    _zz_dataOut_payload_0_9928 <= _zz_dataOut_payload_0_9560;
    _zz_dataOut_payload_0_9929 <= _zz_dataOut_payload_0_9561;
    _zz_dataOut_payload_0_9930 <= _zz_dataOut_payload_0_9562;
    _zz_dataOut_payload_0_9931 <= _zz_dataOut_payload_0_9563;
    _zz_dataOut_payload_0_9932 <= _zz_dataOut_payload_0_9564;
    _zz_dataOut_payload_0_9933 <= _zz_dataOut_payload_0_9565;
    _zz_dataOut_payload_0_9934 <= _zz_dataOut_payload_0_9566;
    _zz_dataOut_payload_0_9935 <= _zz_dataOut_payload_0_9567;
    _zz_dataOut_payload_0_9936 <= _zz_dataOut_payload_0_9568;
    _zz_dataOut_payload_0_9937 <= _zz_dataOut_payload_0_9569;
    _zz_dataOut_payload_0_9938 <= _zz_dataOut_payload_0_9570;
    _zz_dataOut_payload_0_9939 <= _zz_dataOut_payload_0_9571;
    _zz_dataOut_payload_0_9940 <= _zz_dataOut_payload_0_9572;
    _zz_dataOut_payload_0_9941 <= _zz_dataOut_payload_0_9573;
    _zz_dataOut_payload_0_9942 <= _zz_dataOut_payload_0_9574;
    _zz_dataOut_payload_0_9943 <= _zz_dataOut_payload_0_9575;
    _zz_dataOut_payload_0_9944 <= _zz_dataOut_payload_0_9576;
    _zz_dataOut_payload_0_9945 <= _zz_dataOut_payload_0_9577;
    _zz_dataOut_payload_0_9946 <= _zz_dataOut_payload_0_9578;
    _zz_dataOut_payload_0_9947 <= _zz_dataOut_payload_0_9579;
    _zz_dataOut_payload_0_9948 <= _zz_dataOut_payload_0_9580;
    _zz_dataOut_payload_0_9949 <= _zz_dataOut_payload_0_9581;
    _zz_dataOut_payload_0_9950 <= _zz_dataOut_payload_0_9582;
    _zz_dataOut_payload_0_9951 <= _zz_dataOut_payload_0_9583;
    _zz_dataOut_payload_0_9952 <= _zz_dataOut_payload_0_9888;
    _zz_dataOut_payload_0_9953 <= _zz_dataOut_payload_0_9889;
    _zz_dataOut_payload_0_9954 <= _zz_dataOut_payload_0_9890;
    _zz_dataOut_payload_0_9955 <= _zz_dataOut_payload_0_9891;
    _zz_dataOut_payload_0_9956 <= _zz_dataOut_payload_0_9892;
    _zz_dataOut_payload_0_9957 <= _zz_dataOut_payload_0_9893;
    _zz_dataOut_payload_0_9958 <= _zz_dataOut_payload_0_9894;
    _zz_dataOut_payload_0_9959 <= _zz_dataOut_payload_0_9895;
    _zz_dataOut_payload_0_9960 <= _zz_dataOut_payload_0_9896;
    _zz_dataOut_payload_0_9961 <= _zz_dataOut_payload_0_9897;
    _zz_dataOut_payload_0_9962 <= _zz_dataOut_payload_0_9898;
    _zz_dataOut_payload_0_9963 <= _zz_dataOut_payload_0_9899;
    _zz_dataOut_payload_0_9964 <= _zz_dataOut_payload_0_9900;
    _zz_dataOut_payload_0_9965 <= _zz_dataOut_payload_0_9901;
    _zz_dataOut_payload_0_9966 <= _zz_dataOut_payload_0_9902;
    _zz_dataOut_payload_0_9967 <= _zz_dataOut_payload_0_9903;
    _zz_dataOut_payload_0_9968 <= _zz_dataOut_payload_0_9904;
    _zz_dataOut_payload_0_9969 <= _zz_dataOut_payload_0_9905;
    _zz_dataOut_payload_0_9970 <= _zz_dataOut_payload_0_9906;
    _zz_dataOut_payload_0_9971 <= _zz_dataOut_payload_0_9907;
    _zz_dataOut_payload_0_9972 <= _zz_dataOut_payload_0_9908;
    _zz_dataOut_payload_0_9973 <= _zz_dataOut_payload_0_9909;
    _zz_dataOut_payload_0_9974 <= _zz_dataOut_payload_0_9910;
    _zz_dataOut_payload_0_9975 <= _zz_dataOut_payload_0_9911;
    _zz_dataOut_payload_0_9976 <= _zz_dataOut_payload_0_9912;
    _zz_dataOut_payload_0_9977 <= _zz_dataOut_payload_0_9913;
    _zz_dataOut_payload_0_9978 <= _zz_dataOut_payload_0_9914;
    _zz_dataOut_payload_0_9979 <= _zz_dataOut_payload_0_9915;
    _zz_dataOut_payload_0_9980 <= _zz_dataOut_payload_0_9916;
    _zz_dataOut_payload_0_9981 <= _zz_dataOut_payload_0_9917;
    _zz_dataOut_payload_0_9982 <= _zz_dataOut_payload_0_9918;
    _zz_dataOut_payload_0_9983 <= _zz_dataOut_payload_0_9919;
    _zz_dataOut_payload_0_10172 <= (_zz_dataOut_payload_0_10170 ? _zz_dataOut_payload_0_10165 : _zz_dataOut_payload_0_10168);
    _zz_dataOut_payload_0_10173 <= (_zz_dataOut_payload_0_10170 ? _zz_dataOut_payload_0_10168 : _zz_dataOut_payload_0_10165);
    _zz_dataOut_payload_0_10174 <= (_zz_dataOut_payload_0_10171 ? _zz_dataOut_payload_0_10166 : _zz_dataOut_payload_0_10169);
    _zz_dataOut_payload_0_10175 <= (_zz_dataOut_payload_0_10171 ? _zz_dataOut_payload_0_10169 : _zz_dataOut_payload_0_10166);
    _zz_dataOut_payload_0_10184 <= (_zz_dataOut_payload_0_10182 ? _zz_dataOut_payload_0_10177 : _zz_dataOut_payload_0_10180);
    _zz_dataOut_payload_0_10185 <= (_zz_dataOut_payload_0_10182 ? _zz_dataOut_payload_0_10180 : _zz_dataOut_payload_0_10177);
    _zz_dataOut_payload_0_10186 <= (_zz_dataOut_payload_0_10183 ? _zz_dataOut_payload_0_10178 : _zz_dataOut_payload_0_10181);
    _zz_dataOut_payload_0_10187 <= (_zz_dataOut_payload_0_10183 ? _zz_dataOut_payload_0_10181 : _zz_dataOut_payload_0_10178);
    _zz_dataOut_payload_0_10188 <= _zz_dataOut_payload_0_10172;
    _zz_dataOut_payload_0_10189 <= _zz_dataOut_payload_0_10173;
    _zz_dataOut_payload_0_10190 <= _zz_dataOut_payload_0_10174;
    _zz_dataOut_payload_0_10191 <= _zz_dataOut_payload_0_10175;
    _zz_dataOut_payload_0_10192 <= _zz_dataOut_payload_0_10184;
    _zz_dataOut_payload_0_10193 <= _zz_dataOut_payload_0_10185;
    _zz_dataOut_payload_0_10194 <= _zz_dataOut_payload_0_10186;
    _zz_dataOut_payload_0_10195 <= _zz_dataOut_payload_0_10187;
    _zz_dataOut_payload_0_10216 <= (_zz_dataOut_payload_0_10214 ? _zz_dataOut_payload_0_10209 : _zz_dataOut_payload_0_10212);
    _zz_dataOut_payload_0_10217 <= (_zz_dataOut_payload_0_10214 ? _zz_dataOut_payload_0_10212 : _zz_dataOut_payload_0_10209);
    _zz_dataOut_payload_0_10218 <= (_zz_dataOut_payload_0_10215 ? _zz_dataOut_payload_0_10210 : _zz_dataOut_payload_0_10213);
    _zz_dataOut_payload_0_10219 <= (_zz_dataOut_payload_0_10215 ? _zz_dataOut_payload_0_10213 : _zz_dataOut_payload_0_10210);
    _zz_dataOut_payload_0_10228 <= (_zz_dataOut_payload_0_10226 ? _zz_dataOut_payload_0_10221 : _zz_dataOut_payload_0_10224);
    _zz_dataOut_payload_0_10229 <= (_zz_dataOut_payload_0_10226 ? _zz_dataOut_payload_0_10224 : _zz_dataOut_payload_0_10221);
    _zz_dataOut_payload_0_10230 <= (_zz_dataOut_payload_0_10227 ? _zz_dataOut_payload_0_10222 : _zz_dataOut_payload_0_10225);
    _zz_dataOut_payload_0_10231 <= (_zz_dataOut_payload_0_10227 ? _zz_dataOut_payload_0_10225 : _zz_dataOut_payload_0_10222);
    _zz_dataOut_payload_0_10232 <= _zz_dataOut_payload_0_10216;
    _zz_dataOut_payload_0_10233 <= _zz_dataOut_payload_0_10217;
    _zz_dataOut_payload_0_10234 <= _zz_dataOut_payload_0_10218;
    _zz_dataOut_payload_0_10235 <= _zz_dataOut_payload_0_10219;
    _zz_dataOut_payload_0_10236 <= _zz_dataOut_payload_0_10228;
    _zz_dataOut_payload_0_10237 <= _zz_dataOut_payload_0_10229;
    _zz_dataOut_payload_0_10238 <= _zz_dataOut_payload_0_10230;
    _zz_dataOut_payload_0_10239 <= _zz_dataOut_payload_0_10231;
    _zz_dataOut_payload_0_10240 <= _zz_dataOut_payload_0_10188;
    _zz_dataOut_payload_0_10241 <= _zz_dataOut_payload_0_10189;
    _zz_dataOut_payload_0_10242 <= _zz_dataOut_payload_0_10190;
    _zz_dataOut_payload_0_10243 <= _zz_dataOut_payload_0_10191;
    _zz_dataOut_payload_0_10244 <= _zz_dataOut_payload_0_10192;
    _zz_dataOut_payload_0_10245 <= _zz_dataOut_payload_0_10193;
    _zz_dataOut_payload_0_10246 <= _zz_dataOut_payload_0_10194;
    _zz_dataOut_payload_0_10247 <= _zz_dataOut_payload_0_10195;
    _zz_dataOut_payload_0_10248 <= _zz_dataOut_payload_0_10232;
    _zz_dataOut_payload_0_10249 <= _zz_dataOut_payload_0_10233;
    _zz_dataOut_payload_0_10250 <= _zz_dataOut_payload_0_10234;
    _zz_dataOut_payload_0_10251 <= _zz_dataOut_payload_0_10235;
    _zz_dataOut_payload_0_10252 <= _zz_dataOut_payload_0_10236;
    _zz_dataOut_payload_0_10253 <= _zz_dataOut_payload_0_10237;
    _zz_dataOut_payload_0_10254 <= _zz_dataOut_payload_0_10238;
    _zz_dataOut_payload_0_10255 <= _zz_dataOut_payload_0_10239;
    _zz_dataOut_payload_0_10300 <= (_zz_dataOut_payload_0_10298 ? _zz_dataOut_payload_0_10293 : _zz_dataOut_payload_0_10296);
    _zz_dataOut_payload_0_10301 <= (_zz_dataOut_payload_0_10298 ? _zz_dataOut_payload_0_10296 : _zz_dataOut_payload_0_10293);
    _zz_dataOut_payload_0_10302 <= (_zz_dataOut_payload_0_10299 ? _zz_dataOut_payload_0_10294 : _zz_dataOut_payload_0_10297);
    _zz_dataOut_payload_0_10303 <= (_zz_dataOut_payload_0_10299 ? _zz_dataOut_payload_0_10297 : _zz_dataOut_payload_0_10294);
    _zz_dataOut_payload_0_10312 <= (_zz_dataOut_payload_0_10310 ? _zz_dataOut_payload_0_10305 : _zz_dataOut_payload_0_10308);
    _zz_dataOut_payload_0_10313 <= (_zz_dataOut_payload_0_10310 ? _zz_dataOut_payload_0_10308 : _zz_dataOut_payload_0_10305);
    _zz_dataOut_payload_0_10314 <= (_zz_dataOut_payload_0_10311 ? _zz_dataOut_payload_0_10306 : _zz_dataOut_payload_0_10309);
    _zz_dataOut_payload_0_10315 <= (_zz_dataOut_payload_0_10311 ? _zz_dataOut_payload_0_10309 : _zz_dataOut_payload_0_10306);
    _zz_dataOut_payload_0_10316 <= _zz_dataOut_payload_0_10300;
    _zz_dataOut_payload_0_10317 <= _zz_dataOut_payload_0_10301;
    _zz_dataOut_payload_0_10318 <= _zz_dataOut_payload_0_10302;
    _zz_dataOut_payload_0_10319 <= _zz_dataOut_payload_0_10303;
    _zz_dataOut_payload_0_10320 <= _zz_dataOut_payload_0_10312;
    _zz_dataOut_payload_0_10321 <= _zz_dataOut_payload_0_10313;
    _zz_dataOut_payload_0_10322 <= _zz_dataOut_payload_0_10314;
    _zz_dataOut_payload_0_10323 <= _zz_dataOut_payload_0_10315;
    _zz_dataOut_payload_0_10344 <= (_zz_dataOut_payload_0_10342 ? _zz_dataOut_payload_0_10337 : _zz_dataOut_payload_0_10340);
    _zz_dataOut_payload_0_10345 <= (_zz_dataOut_payload_0_10342 ? _zz_dataOut_payload_0_10340 : _zz_dataOut_payload_0_10337);
    _zz_dataOut_payload_0_10346 <= (_zz_dataOut_payload_0_10343 ? _zz_dataOut_payload_0_10338 : _zz_dataOut_payload_0_10341);
    _zz_dataOut_payload_0_10347 <= (_zz_dataOut_payload_0_10343 ? _zz_dataOut_payload_0_10341 : _zz_dataOut_payload_0_10338);
    _zz_dataOut_payload_0_10356 <= (_zz_dataOut_payload_0_10354 ? _zz_dataOut_payload_0_10349 : _zz_dataOut_payload_0_10352);
    _zz_dataOut_payload_0_10357 <= (_zz_dataOut_payload_0_10354 ? _zz_dataOut_payload_0_10352 : _zz_dataOut_payload_0_10349);
    _zz_dataOut_payload_0_10358 <= (_zz_dataOut_payload_0_10355 ? _zz_dataOut_payload_0_10350 : _zz_dataOut_payload_0_10353);
    _zz_dataOut_payload_0_10359 <= (_zz_dataOut_payload_0_10355 ? _zz_dataOut_payload_0_10353 : _zz_dataOut_payload_0_10350);
    _zz_dataOut_payload_0_10360 <= _zz_dataOut_payload_0_10344;
    _zz_dataOut_payload_0_10361 <= _zz_dataOut_payload_0_10345;
    _zz_dataOut_payload_0_10362 <= _zz_dataOut_payload_0_10346;
    _zz_dataOut_payload_0_10363 <= _zz_dataOut_payload_0_10347;
    _zz_dataOut_payload_0_10364 <= _zz_dataOut_payload_0_10356;
    _zz_dataOut_payload_0_10365 <= _zz_dataOut_payload_0_10357;
    _zz_dataOut_payload_0_10366 <= _zz_dataOut_payload_0_10358;
    _zz_dataOut_payload_0_10367 <= _zz_dataOut_payload_0_10359;
    _zz_dataOut_payload_0_10368 <= _zz_dataOut_payload_0_10316;
    _zz_dataOut_payload_0_10369 <= _zz_dataOut_payload_0_10317;
    _zz_dataOut_payload_0_10370 <= _zz_dataOut_payload_0_10318;
    _zz_dataOut_payload_0_10371 <= _zz_dataOut_payload_0_10319;
    _zz_dataOut_payload_0_10372 <= _zz_dataOut_payload_0_10320;
    _zz_dataOut_payload_0_10373 <= _zz_dataOut_payload_0_10321;
    _zz_dataOut_payload_0_10374 <= _zz_dataOut_payload_0_10322;
    _zz_dataOut_payload_0_10375 <= _zz_dataOut_payload_0_10323;
    _zz_dataOut_payload_0_10376 <= _zz_dataOut_payload_0_10360;
    _zz_dataOut_payload_0_10377 <= _zz_dataOut_payload_0_10361;
    _zz_dataOut_payload_0_10378 <= _zz_dataOut_payload_0_10362;
    _zz_dataOut_payload_0_10379 <= _zz_dataOut_payload_0_10363;
    _zz_dataOut_payload_0_10380 <= _zz_dataOut_payload_0_10364;
    _zz_dataOut_payload_0_10381 <= _zz_dataOut_payload_0_10365;
    _zz_dataOut_payload_0_10382 <= _zz_dataOut_payload_0_10366;
    _zz_dataOut_payload_0_10383 <= _zz_dataOut_payload_0_10367;
    _zz_dataOut_payload_0_10384 <= _zz_dataOut_payload_0_10240;
    _zz_dataOut_payload_0_10385 <= _zz_dataOut_payload_0_10241;
    _zz_dataOut_payload_0_10386 <= _zz_dataOut_payload_0_10242;
    _zz_dataOut_payload_0_10387 <= _zz_dataOut_payload_0_10243;
    _zz_dataOut_payload_0_10388 <= _zz_dataOut_payload_0_10244;
    _zz_dataOut_payload_0_10389 <= _zz_dataOut_payload_0_10245;
    _zz_dataOut_payload_0_10390 <= _zz_dataOut_payload_0_10246;
    _zz_dataOut_payload_0_10391 <= _zz_dataOut_payload_0_10247;
    _zz_dataOut_payload_0_10392 <= _zz_dataOut_payload_0_10248;
    _zz_dataOut_payload_0_10393 <= _zz_dataOut_payload_0_10249;
    _zz_dataOut_payload_0_10394 <= _zz_dataOut_payload_0_10250;
    _zz_dataOut_payload_0_10395 <= _zz_dataOut_payload_0_10251;
    _zz_dataOut_payload_0_10396 <= _zz_dataOut_payload_0_10252;
    _zz_dataOut_payload_0_10397 <= _zz_dataOut_payload_0_10253;
    _zz_dataOut_payload_0_10398 <= _zz_dataOut_payload_0_10254;
    _zz_dataOut_payload_0_10399 <= _zz_dataOut_payload_0_10255;
    _zz_dataOut_payload_0_10400 <= _zz_dataOut_payload_0_10368;
    _zz_dataOut_payload_0_10401 <= _zz_dataOut_payload_0_10369;
    _zz_dataOut_payload_0_10402 <= _zz_dataOut_payload_0_10370;
    _zz_dataOut_payload_0_10403 <= _zz_dataOut_payload_0_10371;
    _zz_dataOut_payload_0_10404 <= _zz_dataOut_payload_0_10372;
    _zz_dataOut_payload_0_10405 <= _zz_dataOut_payload_0_10373;
    _zz_dataOut_payload_0_10406 <= _zz_dataOut_payload_0_10374;
    _zz_dataOut_payload_0_10407 <= _zz_dataOut_payload_0_10375;
    _zz_dataOut_payload_0_10408 <= _zz_dataOut_payload_0_10376;
    _zz_dataOut_payload_0_10409 <= _zz_dataOut_payload_0_10377;
    _zz_dataOut_payload_0_10410 <= _zz_dataOut_payload_0_10378;
    _zz_dataOut_payload_0_10411 <= _zz_dataOut_payload_0_10379;
    _zz_dataOut_payload_0_10412 <= _zz_dataOut_payload_0_10380;
    _zz_dataOut_payload_0_10413 <= _zz_dataOut_payload_0_10381;
    _zz_dataOut_payload_0_10414 <= _zz_dataOut_payload_0_10382;
    _zz_dataOut_payload_0_10415 <= _zz_dataOut_payload_0_10383;
    _zz_dataOut_payload_0_10508 <= (_zz_dataOut_payload_0_10506 ? _zz_dataOut_payload_0_10501 : _zz_dataOut_payload_0_10504);
    _zz_dataOut_payload_0_10509 <= (_zz_dataOut_payload_0_10506 ? _zz_dataOut_payload_0_10504 : _zz_dataOut_payload_0_10501);
    _zz_dataOut_payload_0_10510 <= (_zz_dataOut_payload_0_10507 ? _zz_dataOut_payload_0_10502 : _zz_dataOut_payload_0_10505);
    _zz_dataOut_payload_0_10511 <= (_zz_dataOut_payload_0_10507 ? _zz_dataOut_payload_0_10505 : _zz_dataOut_payload_0_10502);
    _zz_dataOut_payload_0_10520 <= (_zz_dataOut_payload_0_10518 ? _zz_dataOut_payload_0_10513 : _zz_dataOut_payload_0_10516);
    _zz_dataOut_payload_0_10521 <= (_zz_dataOut_payload_0_10518 ? _zz_dataOut_payload_0_10516 : _zz_dataOut_payload_0_10513);
    _zz_dataOut_payload_0_10522 <= (_zz_dataOut_payload_0_10519 ? _zz_dataOut_payload_0_10514 : _zz_dataOut_payload_0_10517);
    _zz_dataOut_payload_0_10523 <= (_zz_dataOut_payload_0_10519 ? _zz_dataOut_payload_0_10517 : _zz_dataOut_payload_0_10514);
    _zz_dataOut_payload_0_10524 <= _zz_dataOut_payload_0_10508;
    _zz_dataOut_payload_0_10525 <= _zz_dataOut_payload_0_10509;
    _zz_dataOut_payload_0_10526 <= _zz_dataOut_payload_0_10510;
    _zz_dataOut_payload_0_10527 <= _zz_dataOut_payload_0_10511;
    _zz_dataOut_payload_0_10528 <= _zz_dataOut_payload_0_10520;
    _zz_dataOut_payload_0_10529 <= _zz_dataOut_payload_0_10521;
    _zz_dataOut_payload_0_10530 <= _zz_dataOut_payload_0_10522;
    _zz_dataOut_payload_0_10531 <= _zz_dataOut_payload_0_10523;
    _zz_dataOut_payload_0_10552 <= (_zz_dataOut_payload_0_10550 ? _zz_dataOut_payload_0_10545 : _zz_dataOut_payload_0_10548);
    _zz_dataOut_payload_0_10553 <= (_zz_dataOut_payload_0_10550 ? _zz_dataOut_payload_0_10548 : _zz_dataOut_payload_0_10545);
    _zz_dataOut_payload_0_10554 <= (_zz_dataOut_payload_0_10551 ? _zz_dataOut_payload_0_10546 : _zz_dataOut_payload_0_10549);
    _zz_dataOut_payload_0_10555 <= (_zz_dataOut_payload_0_10551 ? _zz_dataOut_payload_0_10549 : _zz_dataOut_payload_0_10546);
    _zz_dataOut_payload_0_10564 <= (_zz_dataOut_payload_0_10562 ? _zz_dataOut_payload_0_10557 : _zz_dataOut_payload_0_10560);
    _zz_dataOut_payload_0_10565 <= (_zz_dataOut_payload_0_10562 ? _zz_dataOut_payload_0_10560 : _zz_dataOut_payload_0_10557);
    _zz_dataOut_payload_0_10566 <= (_zz_dataOut_payload_0_10563 ? _zz_dataOut_payload_0_10558 : _zz_dataOut_payload_0_10561);
    _zz_dataOut_payload_0_10567 <= (_zz_dataOut_payload_0_10563 ? _zz_dataOut_payload_0_10561 : _zz_dataOut_payload_0_10558);
    _zz_dataOut_payload_0_10568 <= _zz_dataOut_payload_0_10552;
    _zz_dataOut_payload_0_10569 <= _zz_dataOut_payload_0_10553;
    _zz_dataOut_payload_0_10570 <= _zz_dataOut_payload_0_10554;
    _zz_dataOut_payload_0_10571 <= _zz_dataOut_payload_0_10555;
    _zz_dataOut_payload_0_10572 <= _zz_dataOut_payload_0_10564;
    _zz_dataOut_payload_0_10573 <= _zz_dataOut_payload_0_10565;
    _zz_dataOut_payload_0_10574 <= _zz_dataOut_payload_0_10566;
    _zz_dataOut_payload_0_10575 <= _zz_dataOut_payload_0_10567;
    _zz_dataOut_payload_0_10576 <= _zz_dataOut_payload_0_10524;
    _zz_dataOut_payload_0_10577 <= _zz_dataOut_payload_0_10525;
    _zz_dataOut_payload_0_10578 <= _zz_dataOut_payload_0_10526;
    _zz_dataOut_payload_0_10579 <= _zz_dataOut_payload_0_10527;
    _zz_dataOut_payload_0_10580 <= _zz_dataOut_payload_0_10528;
    _zz_dataOut_payload_0_10581 <= _zz_dataOut_payload_0_10529;
    _zz_dataOut_payload_0_10582 <= _zz_dataOut_payload_0_10530;
    _zz_dataOut_payload_0_10583 <= _zz_dataOut_payload_0_10531;
    _zz_dataOut_payload_0_10584 <= _zz_dataOut_payload_0_10568;
    _zz_dataOut_payload_0_10585 <= _zz_dataOut_payload_0_10569;
    _zz_dataOut_payload_0_10586 <= _zz_dataOut_payload_0_10570;
    _zz_dataOut_payload_0_10587 <= _zz_dataOut_payload_0_10571;
    _zz_dataOut_payload_0_10588 <= _zz_dataOut_payload_0_10572;
    _zz_dataOut_payload_0_10589 <= _zz_dataOut_payload_0_10573;
    _zz_dataOut_payload_0_10590 <= _zz_dataOut_payload_0_10574;
    _zz_dataOut_payload_0_10591 <= _zz_dataOut_payload_0_10575;
    _zz_dataOut_payload_0_10636 <= (_zz_dataOut_payload_0_10634 ? _zz_dataOut_payload_0_10629 : _zz_dataOut_payload_0_10632);
    _zz_dataOut_payload_0_10637 <= (_zz_dataOut_payload_0_10634 ? _zz_dataOut_payload_0_10632 : _zz_dataOut_payload_0_10629);
    _zz_dataOut_payload_0_10638 <= (_zz_dataOut_payload_0_10635 ? _zz_dataOut_payload_0_10630 : _zz_dataOut_payload_0_10633);
    _zz_dataOut_payload_0_10639 <= (_zz_dataOut_payload_0_10635 ? _zz_dataOut_payload_0_10633 : _zz_dataOut_payload_0_10630);
    _zz_dataOut_payload_0_10648 <= (_zz_dataOut_payload_0_10646 ? _zz_dataOut_payload_0_10641 : _zz_dataOut_payload_0_10644);
    _zz_dataOut_payload_0_10649 <= (_zz_dataOut_payload_0_10646 ? _zz_dataOut_payload_0_10644 : _zz_dataOut_payload_0_10641);
    _zz_dataOut_payload_0_10650 <= (_zz_dataOut_payload_0_10647 ? _zz_dataOut_payload_0_10642 : _zz_dataOut_payload_0_10645);
    _zz_dataOut_payload_0_10651 <= (_zz_dataOut_payload_0_10647 ? _zz_dataOut_payload_0_10645 : _zz_dataOut_payload_0_10642);
    _zz_dataOut_payload_0_10652 <= _zz_dataOut_payload_0_10636;
    _zz_dataOut_payload_0_10653 <= _zz_dataOut_payload_0_10637;
    _zz_dataOut_payload_0_10654 <= _zz_dataOut_payload_0_10638;
    _zz_dataOut_payload_0_10655 <= _zz_dataOut_payload_0_10639;
    _zz_dataOut_payload_0_10656 <= _zz_dataOut_payload_0_10648;
    _zz_dataOut_payload_0_10657 <= _zz_dataOut_payload_0_10649;
    _zz_dataOut_payload_0_10658 <= _zz_dataOut_payload_0_10650;
    _zz_dataOut_payload_0_10659 <= _zz_dataOut_payload_0_10651;
    _zz_dataOut_payload_0_10680 <= (_zz_dataOut_payload_0_10678 ? _zz_dataOut_payload_0_10673 : _zz_dataOut_payload_0_10676);
    _zz_dataOut_payload_0_10681 <= (_zz_dataOut_payload_0_10678 ? _zz_dataOut_payload_0_10676 : _zz_dataOut_payload_0_10673);
    _zz_dataOut_payload_0_10682 <= (_zz_dataOut_payload_0_10679 ? _zz_dataOut_payload_0_10674 : _zz_dataOut_payload_0_10677);
    _zz_dataOut_payload_0_10683 <= (_zz_dataOut_payload_0_10679 ? _zz_dataOut_payload_0_10677 : _zz_dataOut_payload_0_10674);
    _zz_dataOut_payload_0_10692 <= (_zz_dataOut_payload_0_10690 ? _zz_dataOut_payload_0_10685 : _zz_dataOut_payload_0_10688);
    _zz_dataOut_payload_0_10693 <= (_zz_dataOut_payload_0_10690 ? _zz_dataOut_payload_0_10688 : _zz_dataOut_payload_0_10685);
    _zz_dataOut_payload_0_10694 <= (_zz_dataOut_payload_0_10691 ? _zz_dataOut_payload_0_10686 : _zz_dataOut_payload_0_10689);
    _zz_dataOut_payload_0_10695 <= (_zz_dataOut_payload_0_10691 ? _zz_dataOut_payload_0_10689 : _zz_dataOut_payload_0_10686);
    _zz_dataOut_payload_0_10696 <= _zz_dataOut_payload_0_10680;
    _zz_dataOut_payload_0_10697 <= _zz_dataOut_payload_0_10681;
    _zz_dataOut_payload_0_10698 <= _zz_dataOut_payload_0_10682;
    _zz_dataOut_payload_0_10699 <= _zz_dataOut_payload_0_10683;
    _zz_dataOut_payload_0_10700 <= _zz_dataOut_payload_0_10692;
    _zz_dataOut_payload_0_10701 <= _zz_dataOut_payload_0_10693;
    _zz_dataOut_payload_0_10702 <= _zz_dataOut_payload_0_10694;
    _zz_dataOut_payload_0_10703 <= _zz_dataOut_payload_0_10695;
    _zz_dataOut_payload_0_10704 <= _zz_dataOut_payload_0_10652;
    _zz_dataOut_payload_0_10705 <= _zz_dataOut_payload_0_10653;
    _zz_dataOut_payload_0_10706 <= _zz_dataOut_payload_0_10654;
    _zz_dataOut_payload_0_10707 <= _zz_dataOut_payload_0_10655;
    _zz_dataOut_payload_0_10708 <= _zz_dataOut_payload_0_10656;
    _zz_dataOut_payload_0_10709 <= _zz_dataOut_payload_0_10657;
    _zz_dataOut_payload_0_10710 <= _zz_dataOut_payload_0_10658;
    _zz_dataOut_payload_0_10711 <= _zz_dataOut_payload_0_10659;
    _zz_dataOut_payload_0_10712 <= _zz_dataOut_payload_0_10696;
    _zz_dataOut_payload_0_10713 <= _zz_dataOut_payload_0_10697;
    _zz_dataOut_payload_0_10714 <= _zz_dataOut_payload_0_10698;
    _zz_dataOut_payload_0_10715 <= _zz_dataOut_payload_0_10699;
    _zz_dataOut_payload_0_10716 <= _zz_dataOut_payload_0_10700;
    _zz_dataOut_payload_0_10717 <= _zz_dataOut_payload_0_10701;
    _zz_dataOut_payload_0_10718 <= _zz_dataOut_payload_0_10702;
    _zz_dataOut_payload_0_10719 <= _zz_dataOut_payload_0_10703;
    _zz_dataOut_payload_0_10720 <= _zz_dataOut_payload_0_10576;
    _zz_dataOut_payload_0_10721 <= _zz_dataOut_payload_0_10577;
    _zz_dataOut_payload_0_10722 <= _zz_dataOut_payload_0_10578;
    _zz_dataOut_payload_0_10723 <= _zz_dataOut_payload_0_10579;
    _zz_dataOut_payload_0_10724 <= _zz_dataOut_payload_0_10580;
    _zz_dataOut_payload_0_10725 <= _zz_dataOut_payload_0_10581;
    _zz_dataOut_payload_0_10726 <= _zz_dataOut_payload_0_10582;
    _zz_dataOut_payload_0_10727 <= _zz_dataOut_payload_0_10583;
    _zz_dataOut_payload_0_10728 <= _zz_dataOut_payload_0_10584;
    _zz_dataOut_payload_0_10729 <= _zz_dataOut_payload_0_10585;
    _zz_dataOut_payload_0_10730 <= _zz_dataOut_payload_0_10586;
    _zz_dataOut_payload_0_10731 <= _zz_dataOut_payload_0_10587;
    _zz_dataOut_payload_0_10732 <= _zz_dataOut_payload_0_10588;
    _zz_dataOut_payload_0_10733 <= _zz_dataOut_payload_0_10589;
    _zz_dataOut_payload_0_10734 <= _zz_dataOut_payload_0_10590;
    _zz_dataOut_payload_0_10735 <= _zz_dataOut_payload_0_10591;
    _zz_dataOut_payload_0_10736 <= _zz_dataOut_payload_0_10704;
    _zz_dataOut_payload_0_10737 <= _zz_dataOut_payload_0_10705;
    _zz_dataOut_payload_0_10738 <= _zz_dataOut_payload_0_10706;
    _zz_dataOut_payload_0_10739 <= _zz_dataOut_payload_0_10707;
    _zz_dataOut_payload_0_10740 <= _zz_dataOut_payload_0_10708;
    _zz_dataOut_payload_0_10741 <= _zz_dataOut_payload_0_10709;
    _zz_dataOut_payload_0_10742 <= _zz_dataOut_payload_0_10710;
    _zz_dataOut_payload_0_10743 <= _zz_dataOut_payload_0_10711;
    _zz_dataOut_payload_0_10744 <= _zz_dataOut_payload_0_10712;
    _zz_dataOut_payload_0_10745 <= _zz_dataOut_payload_0_10713;
    _zz_dataOut_payload_0_10746 <= _zz_dataOut_payload_0_10714;
    _zz_dataOut_payload_0_10747 <= _zz_dataOut_payload_0_10715;
    _zz_dataOut_payload_0_10748 <= _zz_dataOut_payload_0_10716;
    _zz_dataOut_payload_0_10749 <= _zz_dataOut_payload_0_10717;
    _zz_dataOut_payload_0_10750 <= _zz_dataOut_payload_0_10718;
    _zz_dataOut_payload_0_10751 <= _zz_dataOut_payload_0_10719;
    _zz_dataOut_payload_0_10752 <= _zz_dataOut_payload_0_10384;
    _zz_dataOut_payload_0_10753 <= _zz_dataOut_payload_0_10385;
    _zz_dataOut_payload_0_10754 <= _zz_dataOut_payload_0_10386;
    _zz_dataOut_payload_0_10755 <= _zz_dataOut_payload_0_10387;
    _zz_dataOut_payload_0_10756 <= _zz_dataOut_payload_0_10388;
    _zz_dataOut_payload_0_10757 <= _zz_dataOut_payload_0_10389;
    _zz_dataOut_payload_0_10758 <= _zz_dataOut_payload_0_10390;
    _zz_dataOut_payload_0_10759 <= _zz_dataOut_payload_0_10391;
    _zz_dataOut_payload_0_10760 <= _zz_dataOut_payload_0_10392;
    _zz_dataOut_payload_0_10761 <= _zz_dataOut_payload_0_10393;
    _zz_dataOut_payload_0_10762 <= _zz_dataOut_payload_0_10394;
    _zz_dataOut_payload_0_10763 <= _zz_dataOut_payload_0_10395;
    _zz_dataOut_payload_0_10764 <= _zz_dataOut_payload_0_10396;
    _zz_dataOut_payload_0_10765 <= _zz_dataOut_payload_0_10397;
    _zz_dataOut_payload_0_10766 <= _zz_dataOut_payload_0_10398;
    _zz_dataOut_payload_0_10767 <= _zz_dataOut_payload_0_10399;
    _zz_dataOut_payload_0_10768 <= _zz_dataOut_payload_0_10400;
    _zz_dataOut_payload_0_10769 <= _zz_dataOut_payload_0_10401;
    _zz_dataOut_payload_0_10770 <= _zz_dataOut_payload_0_10402;
    _zz_dataOut_payload_0_10771 <= _zz_dataOut_payload_0_10403;
    _zz_dataOut_payload_0_10772 <= _zz_dataOut_payload_0_10404;
    _zz_dataOut_payload_0_10773 <= _zz_dataOut_payload_0_10405;
    _zz_dataOut_payload_0_10774 <= _zz_dataOut_payload_0_10406;
    _zz_dataOut_payload_0_10775 <= _zz_dataOut_payload_0_10407;
    _zz_dataOut_payload_0_10776 <= _zz_dataOut_payload_0_10408;
    _zz_dataOut_payload_0_10777 <= _zz_dataOut_payload_0_10409;
    _zz_dataOut_payload_0_10778 <= _zz_dataOut_payload_0_10410;
    _zz_dataOut_payload_0_10779 <= _zz_dataOut_payload_0_10411;
    _zz_dataOut_payload_0_10780 <= _zz_dataOut_payload_0_10412;
    _zz_dataOut_payload_0_10781 <= _zz_dataOut_payload_0_10413;
    _zz_dataOut_payload_0_10782 <= _zz_dataOut_payload_0_10414;
    _zz_dataOut_payload_0_10783 <= _zz_dataOut_payload_0_10415;
    _zz_dataOut_payload_0_10784 <= _zz_dataOut_payload_0_10720;
    _zz_dataOut_payload_0_10785 <= _zz_dataOut_payload_0_10721;
    _zz_dataOut_payload_0_10786 <= _zz_dataOut_payload_0_10722;
    _zz_dataOut_payload_0_10787 <= _zz_dataOut_payload_0_10723;
    _zz_dataOut_payload_0_10788 <= _zz_dataOut_payload_0_10724;
    _zz_dataOut_payload_0_10789 <= _zz_dataOut_payload_0_10725;
    _zz_dataOut_payload_0_10790 <= _zz_dataOut_payload_0_10726;
    _zz_dataOut_payload_0_10791 <= _zz_dataOut_payload_0_10727;
    _zz_dataOut_payload_0_10792 <= _zz_dataOut_payload_0_10728;
    _zz_dataOut_payload_0_10793 <= _zz_dataOut_payload_0_10729;
    _zz_dataOut_payload_0_10794 <= _zz_dataOut_payload_0_10730;
    _zz_dataOut_payload_0_10795 <= _zz_dataOut_payload_0_10731;
    _zz_dataOut_payload_0_10796 <= _zz_dataOut_payload_0_10732;
    _zz_dataOut_payload_0_10797 <= _zz_dataOut_payload_0_10733;
    _zz_dataOut_payload_0_10798 <= _zz_dataOut_payload_0_10734;
    _zz_dataOut_payload_0_10799 <= _zz_dataOut_payload_0_10735;
    _zz_dataOut_payload_0_10800 <= _zz_dataOut_payload_0_10736;
    _zz_dataOut_payload_0_10801 <= _zz_dataOut_payload_0_10737;
    _zz_dataOut_payload_0_10802 <= _zz_dataOut_payload_0_10738;
    _zz_dataOut_payload_0_10803 <= _zz_dataOut_payload_0_10739;
    _zz_dataOut_payload_0_10804 <= _zz_dataOut_payload_0_10740;
    _zz_dataOut_payload_0_10805 <= _zz_dataOut_payload_0_10741;
    _zz_dataOut_payload_0_10806 <= _zz_dataOut_payload_0_10742;
    _zz_dataOut_payload_0_10807 <= _zz_dataOut_payload_0_10743;
    _zz_dataOut_payload_0_10808 <= _zz_dataOut_payload_0_10744;
    _zz_dataOut_payload_0_10809 <= _zz_dataOut_payload_0_10745;
    _zz_dataOut_payload_0_10810 <= _zz_dataOut_payload_0_10746;
    _zz_dataOut_payload_0_10811 <= _zz_dataOut_payload_0_10747;
    _zz_dataOut_payload_0_10812 <= _zz_dataOut_payload_0_10748;
    _zz_dataOut_payload_0_10813 <= _zz_dataOut_payload_0_10749;
    _zz_dataOut_payload_0_10814 <= _zz_dataOut_payload_0_10750;
    _zz_dataOut_payload_0_10815 <= _zz_dataOut_payload_0_10751;
    _zz_dataOut_payload_0_11004 <= (_zz_dataOut_payload_0_11002 ? _zz_dataOut_payload_0_10997 : _zz_dataOut_payload_0_11000);
    _zz_dataOut_payload_0_11005 <= (_zz_dataOut_payload_0_11002 ? _zz_dataOut_payload_0_11000 : _zz_dataOut_payload_0_10997);
    _zz_dataOut_payload_0_11006 <= (_zz_dataOut_payload_0_11003 ? _zz_dataOut_payload_0_10998 : _zz_dataOut_payload_0_11001);
    _zz_dataOut_payload_0_11007 <= (_zz_dataOut_payload_0_11003 ? _zz_dataOut_payload_0_11001 : _zz_dataOut_payload_0_10998);
    _zz_dataOut_payload_0_11016 <= (_zz_dataOut_payload_0_11014 ? _zz_dataOut_payload_0_11009 : _zz_dataOut_payload_0_11012);
    _zz_dataOut_payload_0_11017 <= (_zz_dataOut_payload_0_11014 ? _zz_dataOut_payload_0_11012 : _zz_dataOut_payload_0_11009);
    _zz_dataOut_payload_0_11018 <= (_zz_dataOut_payload_0_11015 ? _zz_dataOut_payload_0_11010 : _zz_dataOut_payload_0_11013);
    _zz_dataOut_payload_0_11019 <= (_zz_dataOut_payload_0_11015 ? _zz_dataOut_payload_0_11013 : _zz_dataOut_payload_0_11010);
    _zz_dataOut_payload_0_11020 <= _zz_dataOut_payload_0_11004;
    _zz_dataOut_payload_0_11021 <= _zz_dataOut_payload_0_11005;
    _zz_dataOut_payload_0_11022 <= _zz_dataOut_payload_0_11006;
    _zz_dataOut_payload_0_11023 <= _zz_dataOut_payload_0_11007;
    _zz_dataOut_payload_0_11024 <= _zz_dataOut_payload_0_11016;
    _zz_dataOut_payload_0_11025 <= _zz_dataOut_payload_0_11017;
    _zz_dataOut_payload_0_11026 <= _zz_dataOut_payload_0_11018;
    _zz_dataOut_payload_0_11027 <= _zz_dataOut_payload_0_11019;
    _zz_dataOut_payload_0_11048 <= (_zz_dataOut_payload_0_11046 ? _zz_dataOut_payload_0_11041 : _zz_dataOut_payload_0_11044);
    _zz_dataOut_payload_0_11049 <= (_zz_dataOut_payload_0_11046 ? _zz_dataOut_payload_0_11044 : _zz_dataOut_payload_0_11041);
    _zz_dataOut_payload_0_11050 <= (_zz_dataOut_payload_0_11047 ? _zz_dataOut_payload_0_11042 : _zz_dataOut_payload_0_11045);
    _zz_dataOut_payload_0_11051 <= (_zz_dataOut_payload_0_11047 ? _zz_dataOut_payload_0_11045 : _zz_dataOut_payload_0_11042);
    _zz_dataOut_payload_0_11060 <= (_zz_dataOut_payload_0_11058 ? _zz_dataOut_payload_0_11053 : _zz_dataOut_payload_0_11056);
    _zz_dataOut_payload_0_11061 <= (_zz_dataOut_payload_0_11058 ? _zz_dataOut_payload_0_11056 : _zz_dataOut_payload_0_11053);
    _zz_dataOut_payload_0_11062 <= (_zz_dataOut_payload_0_11059 ? _zz_dataOut_payload_0_11054 : _zz_dataOut_payload_0_11057);
    _zz_dataOut_payload_0_11063 <= (_zz_dataOut_payload_0_11059 ? _zz_dataOut_payload_0_11057 : _zz_dataOut_payload_0_11054);
    _zz_dataOut_payload_0_11064 <= _zz_dataOut_payload_0_11048;
    _zz_dataOut_payload_0_11065 <= _zz_dataOut_payload_0_11049;
    _zz_dataOut_payload_0_11066 <= _zz_dataOut_payload_0_11050;
    _zz_dataOut_payload_0_11067 <= _zz_dataOut_payload_0_11051;
    _zz_dataOut_payload_0_11068 <= _zz_dataOut_payload_0_11060;
    _zz_dataOut_payload_0_11069 <= _zz_dataOut_payload_0_11061;
    _zz_dataOut_payload_0_11070 <= _zz_dataOut_payload_0_11062;
    _zz_dataOut_payload_0_11071 <= _zz_dataOut_payload_0_11063;
    _zz_dataOut_payload_0_11072 <= _zz_dataOut_payload_0_11020;
    _zz_dataOut_payload_0_11073 <= _zz_dataOut_payload_0_11021;
    _zz_dataOut_payload_0_11074 <= _zz_dataOut_payload_0_11022;
    _zz_dataOut_payload_0_11075 <= _zz_dataOut_payload_0_11023;
    _zz_dataOut_payload_0_11076 <= _zz_dataOut_payload_0_11024;
    _zz_dataOut_payload_0_11077 <= _zz_dataOut_payload_0_11025;
    _zz_dataOut_payload_0_11078 <= _zz_dataOut_payload_0_11026;
    _zz_dataOut_payload_0_11079 <= _zz_dataOut_payload_0_11027;
    _zz_dataOut_payload_0_11080 <= _zz_dataOut_payload_0_11064;
    _zz_dataOut_payload_0_11081 <= _zz_dataOut_payload_0_11065;
    _zz_dataOut_payload_0_11082 <= _zz_dataOut_payload_0_11066;
    _zz_dataOut_payload_0_11083 <= _zz_dataOut_payload_0_11067;
    _zz_dataOut_payload_0_11084 <= _zz_dataOut_payload_0_11068;
    _zz_dataOut_payload_0_11085 <= _zz_dataOut_payload_0_11069;
    _zz_dataOut_payload_0_11086 <= _zz_dataOut_payload_0_11070;
    _zz_dataOut_payload_0_11087 <= _zz_dataOut_payload_0_11071;
    _zz_dataOut_payload_0_11132 <= (_zz_dataOut_payload_0_11130 ? _zz_dataOut_payload_0_11125 : _zz_dataOut_payload_0_11128);
    _zz_dataOut_payload_0_11133 <= (_zz_dataOut_payload_0_11130 ? _zz_dataOut_payload_0_11128 : _zz_dataOut_payload_0_11125);
    _zz_dataOut_payload_0_11134 <= (_zz_dataOut_payload_0_11131 ? _zz_dataOut_payload_0_11126 : _zz_dataOut_payload_0_11129);
    _zz_dataOut_payload_0_11135 <= (_zz_dataOut_payload_0_11131 ? _zz_dataOut_payload_0_11129 : _zz_dataOut_payload_0_11126);
    _zz_dataOut_payload_0_11144 <= (_zz_dataOut_payload_0_11142 ? _zz_dataOut_payload_0_11137 : _zz_dataOut_payload_0_11140);
    _zz_dataOut_payload_0_11145 <= (_zz_dataOut_payload_0_11142 ? _zz_dataOut_payload_0_11140 : _zz_dataOut_payload_0_11137);
    _zz_dataOut_payload_0_11146 <= (_zz_dataOut_payload_0_11143 ? _zz_dataOut_payload_0_11138 : _zz_dataOut_payload_0_11141);
    _zz_dataOut_payload_0_11147 <= (_zz_dataOut_payload_0_11143 ? _zz_dataOut_payload_0_11141 : _zz_dataOut_payload_0_11138);
    _zz_dataOut_payload_0_11148 <= _zz_dataOut_payload_0_11132;
    _zz_dataOut_payload_0_11149 <= _zz_dataOut_payload_0_11133;
    _zz_dataOut_payload_0_11150 <= _zz_dataOut_payload_0_11134;
    _zz_dataOut_payload_0_11151 <= _zz_dataOut_payload_0_11135;
    _zz_dataOut_payload_0_11152 <= _zz_dataOut_payload_0_11144;
    _zz_dataOut_payload_0_11153 <= _zz_dataOut_payload_0_11145;
    _zz_dataOut_payload_0_11154 <= _zz_dataOut_payload_0_11146;
    _zz_dataOut_payload_0_11155 <= _zz_dataOut_payload_0_11147;
    _zz_dataOut_payload_0_11176 <= (_zz_dataOut_payload_0_11174 ? _zz_dataOut_payload_0_11169 : _zz_dataOut_payload_0_11172);
    _zz_dataOut_payload_0_11177 <= (_zz_dataOut_payload_0_11174 ? _zz_dataOut_payload_0_11172 : _zz_dataOut_payload_0_11169);
    _zz_dataOut_payload_0_11178 <= (_zz_dataOut_payload_0_11175 ? _zz_dataOut_payload_0_11170 : _zz_dataOut_payload_0_11173);
    _zz_dataOut_payload_0_11179 <= (_zz_dataOut_payload_0_11175 ? _zz_dataOut_payload_0_11173 : _zz_dataOut_payload_0_11170);
    _zz_dataOut_payload_0_11188 <= (_zz_dataOut_payload_0_11186 ? _zz_dataOut_payload_0_11181 : _zz_dataOut_payload_0_11184);
    _zz_dataOut_payload_0_11189 <= (_zz_dataOut_payload_0_11186 ? _zz_dataOut_payload_0_11184 : _zz_dataOut_payload_0_11181);
    _zz_dataOut_payload_0_11190 <= (_zz_dataOut_payload_0_11187 ? _zz_dataOut_payload_0_11182 : _zz_dataOut_payload_0_11185);
    _zz_dataOut_payload_0_11191 <= (_zz_dataOut_payload_0_11187 ? _zz_dataOut_payload_0_11185 : _zz_dataOut_payload_0_11182);
    _zz_dataOut_payload_0_11192 <= _zz_dataOut_payload_0_11176;
    _zz_dataOut_payload_0_11193 <= _zz_dataOut_payload_0_11177;
    _zz_dataOut_payload_0_11194 <= _zz_dataOut_payload_0_11178;
    _zz_dataOut_payload_0_11195 <= _zz_dataOut_payload_0_11179;
    _zz_dataOut_payload_0_11196 <= _zz_dataOut_payload_0_11188;
    _zz_dataOut_payload_0_11197 <= _zz_dataOut_payload_0_11189;
    _zz_dataOut_payload_0_11198 <= _zz_dataOut_payload_0_11190;
    _zz_dataOut_payload_0_11199 <= _zz_dataOut_payload_0_11191;
    _zz_dataOut_payload_0_11200 <= _zz_dataOut_payload_0_11148;
    _zz_dataOut_payload_0_11201 <= _zz_dataOut_payload_0_11149;
    _zz_dataOut_payload_0_11202 <= _zz_dataOut_payload_0_11150;
    _zz_dataOut_payload_0_11203 <= _zz_dataOut_payload_0_11151;
    _zz_dataOut_payload_0_11204 <= _zz_dataOut_payload_0_11152;
    _zz_dataOut_payload_0_11205 <= _zz_dataOut_payload_0_11153;
    _zz_dataOut_payload_0_11206 <= _zz_dataOut_payload_0_11154;
    _zz_dataOut_payload_0_11207 <= _zz_dataOut_payload_0_11155;
    _zz_dataOut_payload_0_11208 <= _zz_dataOut_payload_0_11192;
    _zz_dataOut_payload_0_11209 <= _zz_dataOut_payload_0_11193;
    _zz_dataOut_payload_0_11210 <= _zz_dataOut_payload_0_11194;
    _zz_dataOut_payload_0_11211 <= _zz_dataOut_payload_0_11195;
    _zz_dataOut_payload_0_11212 <= _zz_dataOut_payload_0_11196;
    _zz_dataOut_payload_0_11213 <= _zz_dataOut_payload_0_11197;
    _zz_dataOut_payload_0_11214 <= _zz_dataOut_payload_0_11198;
    _zz_dataOut_payload_0_11215 <= _zz_dataOut_payload_0_11199;
    _zz_dataOut_payload_0_11216 <= _zz_dataOut_payload_0_11072;
    _zz_dataOut_payload_0_11217 <= _zz_dataOut_payload_0_11073;
    _zz_dataOut_payload_0_11218 <= _zz_dataOut_payload_0_11074;
    _zz_dataOut_payload_0_11219 <= _zz_dataOut_payload_0_11075;
    _zz_dataOut_payload_0_11220 <= _zz_dataOut_payload_0_11076;
    _zz_dataOut_payload_0_11221 <= _zz_dataOut_payload_0_11077;
    _zz_dataOut_payload_0_11222 <= _zz_dataOut_payload_0_11078;
    _zz_dataOut_payload_0_11223 <= _zz_dataOut_payload_0_11079;
    _zz_dataOut_payload_0_11224 <= _zz_dataOut_payload_0_11080;
    _zz_dataOut_payload_0_11225 <= _zz_dataOut_payload_0_11081;
    _zz_dataOut_payload_0_11226 <= _zz_dataOut_payload_0_11082;
    _zz_dataOut_payload_0_11227 <= _zz_dataOut_payload_0_11083;
    _zz_dataOut_payload_0_11228 <= _zz_dataOut_payload_0_11084;
    _zz_dataOut_payload_0_11229 <= _zz_dataOut_payload_0_11085;
    _zz_dataOut_payload_0_11230 <= _zz_dataOut_payload_0_11086;
    _zz_dataOut_payload_0_11231 <= _zz_dataOut_payload_0_11087;
    _zz_dataOut_payload_0_11232 <= _zz_dataOut_payload_0_11200;
    _zz_dataOut_payload_0_11233 <= _zz_dataOut_payload_0_11201;
    _zz_dataOut_payload_0_11234 <= _zz_dataOut_payload_0_11202;
    _zz_dataOut_payload_0_11235 <= _zz_dataOut_payload_0_11203;
    _zz_dataOut_payload_0_11236 <= _zz_dataOut_payload_0_11204;
    _zz_dataOut_payload_0_11237 <= _zz_dataOut_payload_0_11205;
    _zz_dataOut_payload_0_11238 <= _zz_dataOut_payload_0_11206;
    _zz_dataOut_payload_0_11239 <= _zz_dataOut_payload_0_11207;
    _zz_dataOut_payload_0_11240 <= _zz_dataOut_payload_0_11208;
    _zz_dataOut_payload_0_11241 <= _zz_dataOut_payload_0_11209;
    _zz_dataOut_payload_0_11242 <= _zz_dataOut_payload_0_11210;
    _zz_dataOut_payload_0_11243 <= _zz_dataOut_payload_0_11211;
    _zz_dataOut_payload_0_11244 <= _zz_dataOut_payload_0_11212;
    _zz_dataOut_payload_0_11245 <= _zz_dataOut_payload_0_11213;
    _zz_dataOut_payload_0_11246 <= _zz_dataOut_payload_0_11214;
    _zz_dataOut_payload_0_11247 <= _zz_dataOut_payload_0_11215;
    _zz_dataOut_payload_0_11340 <= (_zz_dataOut_payload_0_11338 ? _zz_dataOut_payload_0_11333 : _zz_dataOut_payload_0_11336);
    _zz_dataOut_payload_0_11341 <= (_zz_dataOut_payload_0_11338 ? _zz_dataOut_payload_0_11336 : _zz_dataOut_payload_0_11333);
    _zz_dataOut_payload_0_11342 <= (_zz_dataOut_payload_0_11339 ? _zz_dataOut_payload_0_11334 : _zz_dataOut_payload_0_11337);
    _zz_dataOut_payload_0_11343 <= (_zz_dataOut_payload_0_11339 ? _zz_dataOut_payload_0_11337 : _zz_dataOut_payload_0_11334);
    _zz_dataOut_payload_0_11352 <= (_zz_dataOut_payload_0_11350 ? _zz_dataOut_payload_0_11345 : _zz_dataOut_payload_0_11348);
    _zz_dataOut_payload_0_11353 <= (_zz_dataOut_payload_0_11350 ? _zz_dataOut_payload_0_11348 : _zz_dataOut_payload_0_11345);
    _zz_dataOut_payload_0_11354 <= (_zz_dataOut_payload_0_11351 ? _zz_dataOut_payload_0_11346 : _zz_dataOut_payload_0_11349);
    _zz_dataOut_payload_0_11355 <= (_zz_dataOut_payload_0_11351 ? _zz_dataOut_payload_0_11349 : _zz_dataOut_payload_0_11346);
    _zz_dataOut_payload_0_11356 <= _zz_dataOut_payload_0_11340;
    _zz_dataOut_payload_0_11357 <= _zz_dataOut_payload_0_11341;
    _zz_dataOut_payload_0_11358 <= _zz_dataOut_payload_0_11342;
    _zz_dataOut_payload_0_11359 <= _zz_dataOut_payload_0_11343;
    _zz_dataOut_payload_0_11360 <= _zz_dataOut_payload_0_11352;
    _zz_dataOut_payload_0_11361 <= _zz_dataOut_payload_0_11353;
    _zz_dataOut_payload_0_11362 <= _zz_dataOut_payload_0_11354;
    _zz_dataOut_payload_0_11363 <= _zz_dataOut_payload_0_11355;
    _zz_dataOut_payload_0_11384 <= (_zz_dataOut_payload_0_11382 ? _zz_dataOut_payload_0_11377 : _zz_dataOut_payload_0_11380);
    _zz_dataOut_payload_0_11385 <= (_zz_dataOut_payload_0_11382 ? _zz_dataOut_payload_0_11380 : _zz_dataOut_payload_0_11377);
    _zz_dataOut_payload_0_11386 <= (_zz_dataOut_payload_0_11383 ? _zz_dataOut_payload_0_11378 : _zz_dataOut_payload_0_11381);
    _zz_dataOut_payload_0_11387 <= (_zz_dataOut_payload_0_11383 ? _zz_dataOut_payload_0_11381 : _zz_dataOut_payload_0_11378);
    _zz_dataOut_payload_0_11396 <= (_zz_dataOut_payload_0_11394 ? _zz_dataOut_payload_0_11389 : _zz_dataOut_payload_0_11392);
    _zz_dataOut_payload_0_11397 <= (_zz_dataOut_payload_0_11394 ? _zz_dataOut_payload_0_11392 : _zz_dataOut_payload_0_11389);
    _zz_dataOut_payload_0_11398 <= (_zz_dataOut_payload_0_11395 ? _zz_dataOut_payload_0_11390 : _zz_dataOut_payload_0_11393);
    _zz_dataOut_payload_0_11399 <= (_zz_dataOut_payload_0_11395 ? _zz_dataOut_payload_0_11393 : _zz_dataOut_payload_0_11390);
    _zz_dataOut_payload_0_11400 <= _zz_dataOut_payload_0_11384;
    _zz_dataOut_payload_0_11401 <= _zz_dataOut_payload_0_11385;
    _zz_dataOut_payload_0_11402 <= _zz_dataOut_payload_0_11386;
    _zz_dataOut_payload_0_11403 <= _zz_dataOut_payload_0_11387;
    _zz_dataOut_payload_0_11404 <= _zz_dataOut_payload_0_11396;
    _zz_dataOut_payload_0_11405 <= _zz_dataOut_payload_0_11397;
    _zz_dataOut_payload_0_11406 <= _zz_dataOut_payload_0_11398;
    _zz_dataOut_payload_0_11407 <= _zz_dataOut_payload_0_11399;
    _zz_dataOut_payload_0_11408 <= _zz_dataOut_payload_0_11356;
    _zz_dataOut_payload_0_11409 <= _zz_dataOut_payload_0_11357;
    _zz_dataOut_payload_0_11410 <= _zz_dataOut_payload_0_11358;
    _zz_dataOut_payload_0_11411 <= _zz_dataOut_payload_0_11359;
    _zz_dataOut_payload_0_11412 <= _zz_dataOut_payload_0_11360;
    _zz_dataOut_payload_0_11413 <= _zz_dataOut_payload_0_11361;
    _zz_dataOut_payload_0_11414 <= _zz_dataOut_payload_0_11362;
    _zz_dataOut_payload_0_11415 <= _zz_dataOut_payload_0_11363;
    _zz_dataOut_payload_0_11416 <= _zz_dataOut_payload_0_11400;
    _zz_dataOut_payload_0_11417 <= _zz_dataOut_payload_0_11401;
    _zz_dataOut_payload_0_11418 <= _zz_dataOut_payload_0_11402;
    _zz_dataOut_payload_0_11419 <= _zz_dataOut_payload_0_11403;
    _zz_dataOut_payload_0_11420 <= _zz_dataOut_payload_0_11404;
    _zz_dataOut_payload_0_11421 <= _zz_dataOut_payload_0_11405;
    _zz_dataOut_payload_0_11422 <= _zz_dataOut_payload_0_11406;
    _zz_dataOut_payload_0_11423 <= _zz_dataOut_payload_0_11407;
    _zz_dataOut_payload_0_11468 <= (_zz_dataOut_payload_0_11466 ? _zz_dataOut_payload_0_11461 : _zz_dataOut_payload_0_11464);
    _zz_dataOut_payload_0_11469 <= (_zz_dataOut_payload_0_11466 ? _zz_dataOut_payload_0_11464 : _zz_dataOut_payload_0_11461);
    _zz_dataOut_payload_0_11470 <= (_zz_dataOut_payload_0_11467 ? _zz_dataOut_payload_0_11462 : _zz_dataOut_payload_0_11465);
    _zz_dataOut_payload_0_11471 <= (_zz_dataOut_payload_0_11467 ? _zz_dataOut_payload_0_11465 : _zz_dataOut_payload_0_11462);
    _zz_dataOut_payload_0_11480 <= (_zz_dataOut_payload_0_11478 ? _zz_dataOut_payload_0_11473 : _zz_dataOut_payload_0_11476);
    _zz_dataOut_payload_0_11481 <= (_zz_dataOut_payload_0_11478 ? _zz_dataOut_payload_0_11476 : _zz_dataOut_payload_0_11473);
    _zz_dataOut_payload_0_11482 <= (_zz_dataOut_payload_0_11479 ? _zz_dataOut_payload_0_11474 : _zz_dataOut_payload_0_11477);
    _zz_dataOut_payload_0_11483 <= (_zz_dataOut_payload_0_11479 ? _zz_dataOut_payload_0_11477 : _zz_dataOut_payload_0_11474);
    _zz_dataOut_payload_0_11484 <= _zz_dataOut_payload_0_11468;
    _zz_dataOut_payload_0_11485 <= _zz_dataOut_payload_0_11469;
    _zz_dataOut_payload_0_11486 <= _zz_dataOut_payload_0_11470;
    _zz_dataOut_payload_0_11487 <= _zz_dataOut_payload_0_11471;
    _zz_dataOut_payload_0_11488 <= _zz_dataOut_payload_0_11480;
    _zz_dataOut_payload_0_11489 <= _zz_dataOut_payload_0_11481;
    _zz_dataOut_payload_0_11490 <= _zz_dataOut_payload_0_11482;
    _zz_dataOut_payload_0_11491 <= _zz_dataOut_payload_0_11483;
    _zz_dataOut_payload_0_11512 <= (_zz_dataOut_payload_0_11510 ? _zz_dataOut_payload_0_11505 : _zz_dataOut_payload_0_11508);
    _zz_dataOut_payload_0_11513 <= (_zz_dataOut_payload_0_11510 ? _zz_dataOut_payload_0_11508 : _zz_dataOut_payload_0_11505);
    _zz_dataOut_payload_0_11514 <= (_zz_dataOut_payload_0_11511 ? _zz_dataOut_payload_0_11506 : _zz_dataOut_payload_0_11509);
    _zz_dataOut_payload_0_11515 <= (_zz_dataOut_payload_0_11511 ? _zz_dataOut_payload_0_11509 : _zz_dataOut_payload_0_11506);
    _zz_dataOut_payload_0_11524 <= (_zz_dataOut_payload_0_11522 ? _zz_dataOut_payload_0_11517 : _zz_dataOut_payload_0_11520);
    _zz_dataOut_payload_0_11525 <= (_zz_dataOut_payload_0_11522 ? _zz_dataOut_payload_0_11520 : _zz_dataOut_payload_0_11517);
    _zz_dataOut_payload_0_11526 <= (_zz_dataOut_payload_0_11523 ? _zz_dataOut_payload_0_11518 : _zz_dataOut_payload_0_11521);
    _zz_dataOut_payload_0_11527 <= (_zz_dataOut_payload_0_11523 ? _zz_dataOut_payload_0_11521 : _zz_dataOut_payload_0_11518);
    _zz_dataOut_payload_0_11528 <= _zz_dataOut_payload_0_11512;
    _zz_dataOut_payload_0_11529 <= _zz_dataOut_payload_0_11513;
    _zz_dataOut_payload_0_11530 <= _zz_dataOut_payload_0_11514;
    _zz_dataOut_payload_0_11531 <= _zz_dataOut_payload_0_11515;
    _zz_dataOut_payload_0_11532 <= _zz_dataOut_payload_0_11524;
    _zz_dataOut_payload_0_11533 <= _zz_dataOut_payload_0_11525;
    _zz_dataOut_payload_0_11534 <= _zz_dataOut_payload_0_11526;
    _zz_dataOut_payload_0_11535 <= _zz_dataOut_payload_0_11527;
    _zz_dataOut_payload_0_11536 <= _zz_dataOut_payload_0_11484;
    _zz_dataOut_payload_0_11537 <= _zz_dataOut_payload_0_11485;
    _zz_dataOut_payload_0_11538 <= _zz_dataOut_payload_0_11486;
    _zz_dataOut_payload_0_11539 <= _zz_dataOut_payload_0_11487;
    _zz_dataOut_payload_0_11540 <= _zz_dataOut_payload_0_11488;
    _zz_dataOut_payload_0_11541 <= _zz_dataOut_payload_0_11489;
    _zz_dataOut_payload_0_11542 <= _zz_dataOut_payload_0_11490;
    _zz_dataOut_payload_0_11543 <= _zz_dataOut_payload_0_11491;
    _zz_dataOut_payload_0_11544 <= _zz_dataOut_payload_0_11528;
    _zz_dataOut_payload_0_11545 <= _zz_dataOut_payload_0_11529;
    _zz_dataOut_payload_0_11546 <= _zz_dataOut_payload_0_11530;
    _zz_dataOut_payload_0_11547 <= _zz_dataOut_payload_0_11531;
    _zz_dataOut_payload_0_11548 <= _zz_dataOut_payload_0_11532;
    _zz_dataOut_payload_0_11549 <= _zz_dataOut_payload_0_11533;
    _zz_dataOut_payload_0_11550 <= _zz_dataOut_payload_0_11534;
    _zz_dataOut_payload_0_11551 <= _zz_dataOut_payload_0_11535;
    _zz_dataOut_payload_0_11552 <= _zz_dataOut_payload_0_11408;
    _zz_dataOut_payload_0_11553 <= _zz_dataOut_payload_0_11409;
    _zz_dataOut_payload_0_11554 <= _zz_dataOut_payload_0_11410;
    _zz_dataOut_payload_0_11555 <= _zz_dataOut_payload_0_11411;
    _zz_dataOut_payload_0_11556 <= _zz_dataOut_payload_0_11412;
    _zz_dataOut_payload_0_11557 <= _zz_dataOut_payload_0_11413;
    _zz_dataOut_payload_0_11558 <= _zz_dataOut_payload_0_11414;
    _zz_dataOut_payload_0_11559 <= _zz_dataOut_payload_0_11415;
    _zz_dataOut_payload_0_11560 <= _zz_dataOut_payload_0_11416;
    _zz_dataOut_payload_0_11561 <= _zz_dataOut_payload_0_11417;
    _zz_dataOut_payload_0_11562 <= _zz_dataOut_payload_0_11418;
    _zz_dataOut_payload_0_11563 <= _zz_dataOut_payload_0_11419;
    _zz_dataOut_payload_0_11564 <= _zz_dataOut_payload_0_11420;
    _zz_dataOut_payload_0_11565 <= _zz_dataOut_payload_0_11421;
    _zz_dataOut_payload_0_11566 <= _zz_dataOut_payload_0_11422;
    _zz_dataOut_payload_0_11567 <= _zz_dataOut_payload_0_11423;
    _zz_dataOut_payload_0_11568 <= _zz_dataOut_payload_0_11536;
    _zz_dataOut_payload_0_11569 <= _zz_dataOut_payload_0_11537;
    _zz_dataOut_payload_0_11570 <= _zz_dataOut_payload_0_11538;
    _zz_dataOut_payload_0_11571 <= _zz_dataOut_payload_0_11539;
    _zz_dataOut_payload_0_11572 <= _zz_dataOut_payload_0_11540;
    _zz_dataOut_payload_0_11573 <= _zz_dataOut_payload_0_11541;
    _zz_dataOut_payload_0_11574 <= _zz_dataOut_payload_0_11542;
    _zz_dataOut_payload_0_11575 <= _zz_dataOut_payload_0_11543;
    _zz_dataOut_payload_0_11576 <= _zz_dataOut_payload_0_11544;
    _zz_dataOut_payload_0_11577 <= _zz_dataOut_payload_0_11545;
    _zz_dataOut_payload_0_11578 <= _zz_dataOut_payload_0_11546;
    _zz_dataOut_payload_0_11579 <= _zz_dataOut_payload_0_11547;
    _zz_dataOut_payload_0_11580 <= _zz_dataOut_payload_0_11548;
    _zz_dataOut_payload_0_11581 <= _zz_dataOut_payload_0_11549;
    _zz_dataOut_payload_0_11582 <= _zz_dataOut_payload_0_11550;
    _zz_dataOut_payload_0_11583 <= _zz_dataOut_payload_0_11551;
    _zz_dataOut_payload_0_11584 <= _zz_dataOut_payload_0_11216;
    _zz_dataOut_payload_0_11585 <= _zz_dataOut_payload_0_11217;
    _zz_dataOut_payload_0_11586 <= _zz_dataOut_payload_0_11218;
    _zz_dataOut_payload_0_11587 <= _zz_dataOut_payload_0_11219;
    _zz_dataOut_payload_0_11588 <= _zz_dataOut_payload_0_11220;
    _zz_dataOut_payload_0_11589 <= _zz_dataOut_payload_0_11221;
    _zz_dataOut_payload_0_11590 <= _zz_dataOut_payload_0_11222;
    _zz_dataOut_payload_0_11591 <= _zz_dataOut_payload_0_11223;
    _zz_dataOut_payload_0_11592 <= _zz_dataOut_payload_0_11224;
    _zz_dataOut_payload_0_11593 <= _zz_dataOut_payload_0_11225;
    _zz_dataOut_payload_0_11594 <= _zz_dataOut_payload_0_11226;
    _zz_dataOut_payload_0_11595 <= _zz_dataOut_payload_0_11227;
    _zz_dataOut_payload_0_11596 <= _zz_dataOut_payload_0_11228;
    _zz_dataOut_payload_0_11597 <= _zz_dataOut_payload_0_11229;
    _zz_dataOut_payload_0_11598 <= _zz_dataOut_payload_0_11230;
    _zz_dataOut_payload_0_11599 <= _zz_dataOut_payload_0_11231;
    _zz_dataOut_payload_0_11600 <= _zz_dataOut_payload_0_11232;
    _zz_dataOut_payload_0_11601 <= _zz_dataOut_payload_0_11233;
    _zz_dataOut_payload_0_11602 <= _zz_dataOut_payload_0_11234;
    _zz_dataOut_payload_0_11603 <= _zz_dataOut_payload_0_11235;
    _zz_dataOut_payload_0_11604 <= _zz_dataOut_payload_0_11236;
    _zz_dataOut_payload_0_11605 <= _zz_dataOut_payload_0_11237;
    _zz_dataOut_payload_0_11606 <= _zz_dataOut_payload_0_11238;
    _zz_dataOut_payload_0_11607 <= _zz_dataOut_payload_0_11239;
    _zz_dataOut_payload_0_11608 <= _zz_dataOut_payload_0_11240;
    _zz_dataOut_payload_0_11609 <= _zz_dataOut_payload_0_11241;
    _zz_dataOut_payload_0_11610 <= _zz_dataOut_payload_0_11242;
    _zz_dataOut_payload_0_11611 <= _zz_dataOut_payload_0_11243;
    _zz_dataOut_payload_0_11612 <= _zz_dataOut_payload_0_11244;
    _zz_dataOut_payload_0_11613 <= _zz_dataOut_payload_0_11245;
    _zz_dataOut_payload_0_11614 <= _zz_dataOut_payload_0_11246;
    _zz_dataOut_payload_0_11615 <= _zz_dataOut_payload_0_11247;
    _zz_dataOut_payload_0_11616 <= _zz_dataOut_payload_0_11552;
    _zz_dataOut_payload_0_11617 <= _zz_dataOut_payload_0_11553;
    _zz_dataOut_payload_0_11618 <= _zz_dataOut_payload_0_11554;
    _zz_dataOut_payload_0_11619 <= _zz_dataOut_payload_0_11555;
    _zz_dataOut_payload_0_11620 <= _zz_dataOut_payload_0_11556;
    _zz_dataOut_payload_0_11621 <= _zz_dataOut_payload_0_11557;
    _zz_dataOut_payload_0_11622 <= _zz_dataOut_payload_0_11558;
    _zz_dataOut_payload_0_11623 <= _zz_dataOut_payload_0_11559;
    _zz_dataOut_payload_0_11624 <= _zz_dataOut_payload_0_11560;
    _zz_dataOut_payload_0_11625 <= _zz_dataOut_payload_0_11561;
    _zz_dataOut_payload_0_11626 <= _zz_dataOut_payload_0_11562;
    _zz_dataOut_payload_0_11627 <= _zz_dataOut_payload_0_11563;
    _zz_dataOut_payload_0_11628 <= _zz_dataOut_payload_0_11564;
    _zz_dataOut_payload_0_11629 <= _zz_dataOut_payload_0_11565;
    _zz_dataOut_payload_0_11630 <= _zz_dataOut_payload_0_11566;
    _zz_dataOut_payload_0_11631 <= _zz_dataOut_payload_0_11567;
    _zz_dataOut_payload_0_11632 <= _zz_dataOut_payload_0_11568;
    _zz_dataOut_payload_0_11633 <= _zz_dataOut_payload_0_11569;
    _zz_dataOut_payload_0_11634 <= _zz_dataOut_payload_0_11570;
    _zz_dataOut_payload_0_11635 <= _zz_dataOut_payload_0_11571;
    _zz_dataOut_payload_0_11636 <= _zz_dataOut_payload_0_11572;
    _zz_dataOut_payload_0_11637 <= _zz_dataOut_payload_0_11573;
    _zz_dataOut_payload_0_11638 <= _zz_dataOut_payload_0_11574;
    _zz_dataOut_payload_0_11639 <= _zz_dataOut_payload_0_11575;
    _zz_dataOut_payload_0_11640 <= _zz_dataOut_payload_0_11576;
    _zz_dataOut_payload_0_11641 <= _zz_dataOut_payload_0_11577;
    _zz_dataOut_payload_0_11642 <= _zz_dataOut_payload_0_11578;
    _zz_dataOut_payload_0_11643 <= _zz_dataOut_payload_0_11579;
    _zz_dataOut_payload_0_11644 <= _zz_dataOut_payload_0_11580;
    _zz_dataOut_payload_0_11645 <= _zz_dataOut_payload_0_11581;
    _zz_dataOut_payload_0_11646 <= _zz_dataOut_payload_0_11582;
    _zz_dataOut_payload_0_11647 <= _zz_dataOut_payload_0_11583;
    _zz_dataOut_payload_0_11648 <= _zz_dataOut_payload_0_9088;
    _zz_dataOut_payload_0_11649 <= _zz_dataOut_payload_0_9089;
    _zz_dataOut_payload_0_11650 <= _zz_dataOut_payload_0_9090;
    _zz_dataOut_payload_0_11651 <= _zz_dataOut_payload_0_9091;
    _zz_dataOut_payload_0_11652 <= _zz_dataOut_payload_0_9092;
    _zz_dataOut_payload_0_11653 <= _zz_dataOut_payload_0_9093;
    _zz_dataOut_payload_0_11654 <= _zz_dataOut_payload_0_9094;
    _zz_dataOut_payload_0_11655 <= _zz_dataOut_payload_0_9095;
    _zz_dataOut_payload_0_11656 <= _zz_dataOut_payload_0_9096;
    _zz_dataOut_payload_0_11657 <= _zz_dataOut_payload_0_9097;
    _zz_dataOut_payload_0_11658 <= _zz_dataOut_payload_0_9098;
    _zz_dataOut_payload_0_11659 <= _zz_dataOut_payload_0_9099;
    _zz_dataOut_payload_0_11660 <= _zz_dataOut_payload_0_9100;
    _zz_dataOut_payload_0_11661 <= _zz_dataOut_payload_0_9101;
    _zz_dataOut_payload_0_11662 <= _zz_dataOut_payload_0_9102;
    _zz_dataOut_payload_0_11663 <= _zz_dataOut_payload_0_9103;
    _zz_dataOut_payload_0_11664 <= _zz_dataOut_payload_0_9104;
    _zz_dataOut_payload_0_11665 <= _zz_dataOut_payload_0_9105;
    _zz_dataOut_payload_0_11666 <= _zz_dataOut_payload_0_9106;
    _zz_dataOut_payload_0_11667 <= _zz_dataOut_payload_0_9107;
    _zz_dataOut_payload_0_11668 <= _zz_dataOut_payload_0_9108;
    _zz_dataOut_payload_0_11669 <= _zz_dataOut_payload_0_9109;
    _zz_dataOut_payload_0_11670 <= _zz_dataOut_payload_0_9110;
    _zz_dataOut_payload_0_11671 <= _zz_dataOut_payload_0_9111;
    _zz_dataOut_payload_0_11672 <= _zz_dataOut_payload_0_9112;
    _zz_dataOut_payload_0_11673 <= _zz_dataOut_payload_0_9113;
    _zz_dataOut_payload_0_11674 <= _zz_dataOut_payload_0_9114;
    _zz_dataOut_payload_0_11675 <= _zz_dataOut_payload_0_9115;
    _zz_dataOut_payload_0_11676 <= _zz_dataOut_payload_0_9116;
    _zz_dataOut_payload_0_11677 <= _zz_dataOut_payload_0_9117;
    _zz_dataOut_payload_0_11678 <= _zz_dataOut_payload_0_9118;
    _zz_dataOut_payload_0_11679 <= _zz_dataOut_payload_0_9119;
    _zz_dataOut_payload_0_11680 <= _zz_dataOut_payload_0_9120;
    _zz_dataOut_payload_0_11681 <= _zz_dataOut_payload_0_9121;
    _zz_dataOut_payload_0_11682 <= _zz_dataOut_payload_0_9122;
    _zz_dataOut_payload_0_11683 <= _zz_dataOut_payload_0_9123;
    _zz_dataOut_payload_0_11684 <= _zz_dataOut_payload_0_9124;
    _zz_dataOut_payload_0_11685 <= _zz_dataOut_payload_0_9125;
    _zz_dataOut_payload_0_11686 <= _zz_dataOut_payload_0_9126;
    _zz_dataOut_payload_0_11687 <= _zz_dataOut_payload_0_9127;
    _zz_dataOut_payload_0_11688 <= _zz_dataOut_payload_0_9128;
    _zz_dataOut_payload_0_11689 <= _zz_dataOut_payload_0_9129;
    _zz_dataOut_payload_0_11690 <= _zz_dataOut_payload_0_9130;
    _zz_dataOut_payload_0_11691 <= _zz_dataOut_payload_0_9131;
    _zz_dataOut_payload_0_11692 <= _zz_dataOut_payload_0_9132;
    _zz_dataOut_payload_0_11693 <= _zz_dataOut_payload_0_9133;
    _zz_dataOut_payload_0_11694 <= _zz_dataOut_payload_0_9134;
    _zz_dataOut_payload_0_11695 <= _zz_dataOut_payload_0_9135;
    _zz_dataOut_payload_0_11696 <= _zz_dataOut_payload_0_9136;
    _zz_dataOut_payload_0_11697 <= _zz_dataOut_payload_0_9137;
    _zz_dataOut_payload_0_11698 <= _zz_dataOut_payload_0_9138;
    _zz_dataOut_payload_0_11699 <= _zz_dataOut_payload_0_9139;
    _zz_dataOut_payload_0_11700 <= _zz_dataOut_payload_0_9140;
    _zz_dataOut_payload_0_11701 <= _zz_dataOut_payload_0_9141;
    _zz_dataOut_payload_0_11702 <= _zz_dataOut_payload_0_9142;
    _zz_dataOut_payload_0_11703 <= _zz_dataOut_payload_0_9143;
    _zz_dataOut_payload_0_11704 <= _zz_dataOut_payload_0_9144;
    _zz_dataOut_payload_0_11705 <= _zz_dataOut_payload_0_9145;
    _zz_dataOut_payload_0_11706 <= _zz_dataOut_payload_0_9146;
    _zz_dataOut_payload_0_11707 <= _zz_dataOut_payload_0_9147;
    _zz_dataOut_payload_0_11708 <= _zz_dataOut_payload_0_9148;
    _zz_dataOut_payload_0_11709 <= _zz_dataOut_payload_0_9149;
    _zz_dataOut_payload_0_11710 <= _zz_dataOut_payload_0_9150;
    _zz_dataOut_payload_0_11711 <= _zz_dataOut_payload_0_9151;
    _zz_dataOut_payload_0_11712 <= _zz_dataOut_payload_0_9920;
    _zz_dataOut_payload_0_11713 <= _zz_dataOut_payload_0_9921;
    _zz_dataOut_payload_0_11714 <= _zz_dataOut_payload_0_9922;
    _zz_dataOut_payload_0_11715 <= _zz_dataOut_payload_0_9923;
    _zz_dataOut_payload_0_11716 <= _zz_dataOut_payload_0_9924;
    _zz_dataOut_payload_0_11717 <= _zz_dataOut_payload_0_9925;
    _zz_dataOut_payload_0_11718 <= _zz_dataOut_payload_0_9926;
    _zz_dataOut_payload_0_11719 <= _zz_dataOut_payload_0_9927;
    _zz_dataOut_payload_0_11720 <= _zz_dataOut_payload_0_9928;
    _zz_dataOut_payload_0_11721 <= _zz_dataOut_payload_0_9929;
    _zz_dataOut_payload_0_11722 <= _zz_dataOut_payload_0_9930;
    _zz_dataOut_payload_0_11723 <= _zz_dataOut_payload_0_9931;
    _zz_dataOut_payload_0_11724 <= _zz_dataOut_payload_0_9932;
    _zz_dataOut_payload_0_11725 <= _zz_dataOut_payload_0_9933;
    _zz_dataOut_payload_0_11726 <= _zz_dataOut_payload_0_9934;
    _zz_dataOut_payload_0_11727 <= _zz_dataOut_payload_0_9935;
    _zz_dataOut_payload_0_11728 <= _zz_dataOut_payload_0_9936;
    _zz_dataOut_payload_0_11729 <= _zz_dataOut_payload_0_9937;
    _zz_dataOut_payload_0_11730 <= _zz_dataOut_payload_0_9938;
    _zz_dataOut_payload_0_11731 <= _zz_dataOut_payload_0_9939;
    _zz_dataOut_payload_0_11732 <= _zz_dataOut_payload_0_9940;
    _zz_dataOut_payload_0_11733 <= _zz_dataOut_payload_0_9941;
    _zz_dataOut_payload_0_11734 <= _zz_dataOut_payload_0_9942;
    _zz_dataOut_payload_0_11735 <= _zz_dataOut_payload_0_9943;
    _zz_dataOut_payload_0_11736 <= _zz_dataOut_payload_0_9944;
    _zz_dataOut_payload_0_11737 <= _zz_dataOut_payload_0_9945;
    _zz_dataOut_payload_0_11738 <= _zz_dataOut_payload_0_9946;
    _zz_dataOut_payload_0_11739 <= _zz_dataOut_payload_0_9947;
    _zz_dataOut_payload_0_11740 <= _zz_dataOut_payload_0_9948;
    _zz_dataOut_payload_0_11741 <= _zz_dataOut_payload_0_9949;
    _zz_dataOut_payload_0_11742 <= _zz_dataOut_payload_0_9950;
    _zz_dataOut_payload_0_11743 <= _zz_dataOut_payload_0_9951;
    _zz_dataOut_payload_0_11744 <= _zz_dataOut_payload_0_9952;
    _zz_dataOut_payload_0_11745 <= _zz_dataOut_payload_0_9953;
    _zz_dataOut_payload_0_11746 <= _zz_dataOut_payload_0_9954;
    _zz_dataOut_payload_0_11747 <= _zz_dataOut_payload_0_9955;
    _zz_dataOut_payload_0_11748 <= _zz_dataOut_payload_0_9956;
    _zz_dataOut_payload_0_11749 <= _zz_dataOut_payload_0_9957;
    _zz_dataOut_payload_0_11750 <= _zz_dataOut_payload_0_9958;
    _zz_dataOut_payload_0_11751 <= _zz_dataOut_payload_0_9959;
    _zz_dataOut_payload_0_11752 <= _zz_dataOut_payload_0_9960;
    _zz_dataOut_payload_0_11753 <= _zz_dataOut_payload_0_9961;
    _zz_dataOut_payload_0_11754 <= _zz_dataOut_payload_0_9962;
    _zz_dataOut_payload_0_11755 <= _zz_dataOut_payload_0_9963;
    _zz_dataOut_payload_0_11756 <= _zz_dataOut_payload_0_9964;
    _zz_dataOut_payload_0_11757 <= _zz_dataOut_payload_0_9965;
    _zz_dataOut_payload_0_11758 <= _zz_dataOut_payload_0_9966;
    _zz_dataOut_payload_0_11759 <= _zz_dataOut_payload_0_9967;
    _zz_dataOut_payload_0_11760 <= _zz_dataOut_payload_0_9968;
    _zz_dataOut_payload_0_11761 <= _zz_dataOut_payload_0_9969;
    _zz_dataOut_payload_0_11762 <= _zz_dataOut_payload_0_9970;
    _zz_dataOut_payload_0_11763 <= _zz_dataOut_payload_0_9971;
    _zz_dataOut_payload_0_11764 <= _zz_dataOut_payload_0_9972;
    _zz_dataOut_payload_0_11765 <= _zz_dataOut_payload_0_9973;
    _zz_dataOut_payload_0_11766 <= _zz_dataOut_payload_0_9974;
    _zz_dataOut_payload_0_11767 <= _zz_dataOut_payload_0_9975;
    _zz_dataOut_payload_0_11768 <= _zz_dataOut_payload_0_9976;
    _zz_dataOut_payload_0_11769 <= _zz_dataOut_payload_0_9977;
    _zz_dataOut_payload_0_11770 <= _zz_dataOut_payload_0_9978;
    _zz_dataOut_payload_0_11771 <= _zz_dataOut_payload_0_9979;
    _zz_dataOut_payload_0_11772 <= _zz_dataOut_payload_0_9980;
    _zz_dataOut_payload_0_11773 <= _zz_dataOut_payload_0_9981;
    _zz_dataOut_payload_0_11774 <= _zz_dataOut_payload_0_9982;
    _zz_dataOut_payload_0_11775 <= _zz_dataOut_payload_0_9983;
    _zz_dataOut_payload_0_11776 <= _zz_dataOut_payload_0_10752;
    _zz_dataOut_payload_0_11777 <= _zz_dataOut_payload_0_10753;
    _zz_dataOut_payload_0_11778 <= _zz_dataOut_payload_0_10754;
    _zz_dataOut_payload_0_11779 <= _zz_dataOut_payload_0_10755;
    _zz_dataOut_payload_0_11780 <= _zz_dataOut_payload_0_10756;
    _zz_dataOut_payload_0_11781 <= _zz_dataOut_payload_0_10757;
    _zz_dataOut_payload_0_11782 <= _zz_dataOut_payload_0_10758;
    _zz_dataOut_payload_0_11783 <= _zz_dataOut_payload_0_10759;
    _zz_dataOut_payload_0_11784 <= _zz_dataOut_payload_0_10760;
    _zz_dataOut_payload_0_11785 <= _zz_dataOut_payload_0_10761;
    _zz_dataOut_payload_0_11786 <= _zz_dataOut_payload_0_10762;
    _zz_dataOut_payload_0_11787 <= _zz_dataOut_payload_0_10763;
    _zz_dataOut_payload_0_11788 <= _zz_dataOut_payload_0_10764;
    _zz_dataOut_payload_0_11789 <= _zz_dataOut_payload_0_10765;
    _zz_dataOut_payload_0_11790 <= _zz_dataOut_payload_0_10766;
    _zz_dataOut_payload_0_11791 <= _zz_dataOut_payload_0_10767;
    _zz_dataOut_payload_0_11792 <= _zz_dataOut_payload_0_10768;
    _zz_dataOut_payload_0_11793 <= _zz_dataOut_payload_0_10769;
    _zz_dataOut_payload_0_11794 <= _zz_dataOut_payload_0_10770;
    _zz_dataOut_payload_0_11795 <= _zz_dataOut_payload_0_10771;
    _zz_dataOut_payload_0_11796 <= _zz_dataOut_payload_0_10772;
    _zz_dataOut_payload_0_11797 <= _zz_dataOut_payload_0_10773;
    _zz_dataOut_payload_0_11798 <= _zz_dataOut_payload_0_10774;
    _zz_dataOut_payload_0_11799 <= _zz_dataOut_payload_0_10775;
    _zz_dataOut_payload_0_11800 <= _zz_dataOut_payload_0_10776;
    _zz_dataOut_payload_0_11801 <= _zz_dataOut_payload_0_10777;
    _zz_dataOut_payload_0_11802 <= _zz_dataOut_payload_0_10778;
    _zz_dataOut_payload_0_11803 <= _zz_dataOut_payload_0_10779;
    _zz_dataOut_payload_0_11804 <= _zz_dataOut_payload_0_10780;
    _zz_dataOut_payload_0_11805 <= _zz_dataOut_payload_0_10781;
    _zz_dataOut_payload_0_11806 <= _zz_dataOut_payload_0_10782;
    _zz_dataOut_payload_0_11807 <= _zz_dataOut_payload_0_10783;
    _zz_dataOut_payload_0_11808 <= _zz_dataOut_payload_0_10784;
    _zz_dataOut_payload_0_11809 <= _zz_dataOut_payload_0_10785;
    _zz_dataOut_payload_0_11810 <= _zz_dataOut_payload_0_10786;
    _zz_dataOut_payload_0_11811 <= _zz_dataOut_payload_0_10787;
    _zz_dataOut_payload_0_11812 <= _zz_dataOut_payload_0_10788;
    _zz_dataOut_payload_0_11813 <= _zz_dataOut_payload_0_10789;
    _zz_dataOut_payload_0_11814 <= _zz_dataOut_payload_0_10790;
    _zz_dataOut_payload_0_11815 <= _zz_dataOut_payload_0_10791;
    _zz_dataOut_payload_0_11816 <= _zz_dataOut_payload_0_10792;
    _zz_dataOut_payload_0_11817 <= _zz_dataOut_payload_0_10793;
    _zz_dataOut_payload_0_11818 <= _zz_dataOut_payload_0_10794;
    _zz_dataOut_payload_0_11819 <= _zz_dataOut_payload_0_10795;
    _zz_dataOut_payload_0_11820 <= _zz_dataOut_payload_0_10796;
    _zz_dataOut_payload_0_11821 <= _zz_dataOut_payload_0_10797;
    _zz_dataOut_payload_0_11822 <= _zz_dataOut_payload_0_10798;
    _zz_dataOut_payload_0_11823 <= _zz_dataOut_payload_0_10799;
    _zz_dataOut_payload_0_11824 <= _zz_dataOut_payload_0_10800;
    _zz_dataOut_payload_0_11825 <= _zz_dataOut_payload_0_10801;
    _zz_dataOut_payload_0_11826 <= _zz_dataOut_payload_0_10802;
    _zz_dataOut_payload_0_11827 <= _zz_dataOut_payload_0_10803;
    _zz_dataOut_payload_0_11828 <= _zz_dataOut_payload_0_10804;
    _zz_dataOut_payload_0_11829 <= _zz_dataOut_payload_0_10805;
    _zz_dataOut_payload_0_11830 <= _zz_dataOut_payload_0_10806;
    _zz_dataOut_payload_0_11831 <= _zz_dataOut_payload_0_10807;
    _zz_dataOut_payload_0_11832 <= _zz_dataOut_payload_0_10808;
    _zz_dataOut_payload_0_11833 <= _zz_dataOut_payload_0_10809;
    _zz_dataOut_payload_0_11834 <= _zz_dataOut_payload_0_10810;
    _zz_dataOut_payload_0_11835 <= _zz_dataOut_payload_0_10811;
    _zz_dataOut_payload_0_11836 <= _zz_dataOut_payload_0_10812;
    _zz_dataOut_payload_0_11837 <= _zz_dataOut_payload_0_10813;
    _zz_dataOut_payload_0_11838 <= _zz_dataOut_payload_0_10814;
    _zz_dataOut_payload_0_11839 <= _zz_dataOut_payload_0_10815;
    _zz_dataOut_payload_0_11840 <= _zz_dataOut_payload_0_11584;
    _zz_dataOut_payload_0_11841 <= _zz_dataOut_payload_0_11585;
    _zz_dataOut_payload_0_11842 <= _zz_dataOut_payload_0_11586;
    _zz_dataOut_payload_0_11843 <= _zz_dataOut_payload_0_11587;
    _zz_dataOut_payload_0_11844 <= _zz_dataOut_payload_0_11588;
    _zz_dataOut_payload_0_11845 <= _zz_dataOut_payload_0_11589;
    _zz_dataOut_payload_0_11846 <= _zz_dataOut_payload_0_11590;
    _zz_dataOut_payload_0_11847 <= _zz_dataOut_payload_0_11591;
    _zz_dataOut_payload_0_11848 <= _zz_dataOut_payload_0_11592;
    _zz_dataOut_payload_0_11849 <= _zz_dataOut_payload_0_11593;
    _zz_dataOut_payload_0_11850 <= _zz_dataOut_payload_0_11594;
    _zz_dataOut_payload_0_11851 <= _zz_dataOut_payload_0_11595;
    _zz_dataOut_payload_0_11852 <= _zz_dataOut_payload_0_11596;
    _zz_dataOut_payload_0_11853 <= _zz_dataOut_payload_0_11597;
    _zz_dataOut_payload_0_11854 <= _zz_dataOut_payload_0_11598;
    _zz_dataOut_payload_0_11855 <= _zz_dataOut_payload_0_11599;
    _zz_dataOut_payload_0_11856 <= _zz_dataOut_payload_0_11600;
    _zz_dataOut_payload_0_11857 <= _zz_dataOut_payload_0_11601;
    _zz_dataOut_payload_0_11858 <= _zz_dataOut_payload_0_11602;
    _zz_dataOut_payload_0_11859 <= _zz_dataOut_payload_0_11603;
    _zz_dataOut_payload_0_11860 <= _zz_dataOut_payload_0_11604;
    _zz_dataOut_payload_0_11861 <= _zz_dataOut_payload_0_11605;
    _zz_dataOut_payload_0_11862 <= _zz_dataOut_payload_0_11606;
    _zz_dataOut_payload_0_11863 <= _zz_dataOut_payload_0_11607;
    _zz_dataOut_payload_0_11864 <= _zz_dataOut_payload_0_11608;
    _zz_dataOut_payload_0_11865 <= _zz_dataOut_payload_0_11609;
    _zz_dataOut_payload_0_11866 <= _zz_dataOut_payload_0_11610;
    _zz_dataOut_payload_0_11867 <= _zz_dataOut_payload_0_11611;
    _zz_dataOut_payload_0_11868 <= _zz_dataOut_payload_0_11612;
    _zz_dataOut_payload_0_11869 <= _zz_dataOut_payload_0_11613;
    _zz_dataOut_payload_0_11870 <= _zz_dataOut_payload_0_11614;
    _zz_dataOut_payload_0_11871 <= _zz_dataOut_payload_0_11615;
    _zz_dataOut_payload_0_11872 <= _zz_dataOut_payload_0_11616;
    _zz_dataOut_payload_0_11873 <= _zz_dataOut_payload_0_11617;
    _zz_dataOut_payload_0_11874 <= _zz_dataOut_payload_0_11618;
    _zz_dataOut_payload_0_11875 <= _zz_dataOut_payload_0_11619;
    _zz_dataOut_payload_0_11876 <= _zz_dataOut_payload_0_11620;
    _zz_dataOut_payload_0_11877 <= _zz_dataOut_payload_0_11621;
    _zz_dataOut_payload_0_11878 <= _zz_dataOut_payload_0_11622;
    _zz_dataOut_payload_0_11879 <= _zz_dataOut_payload_0_11623;
    _zz_dataOut_payload_0_11880 <= _zz_dataOut_payload_0_11624;
    _zz_dataOut_payload_0_11881 <= _zz_dataOut_payload_0_11625;
    _zz_dataOut_payload_0_11882 <= _zz_dataOut_payload_0_11626;
    _zz_dataOut_payload_0_11883 <= _zz_dataOut_payload_0_11627;
    _zz_dataOut_payload_0_11884 <= _zz_dataOut_payload_0_11628;
    _zz_dataOut_payload_0_11885 <= _zz_dataOut_payload_0_11629;
    _zz_dataOut_payload_0_11886 <= _zz_dataOut_payload_0_11630;
    _zz_dataOut_payload_0_11887 <= _zz_dataOut_payload_0_11631;
    _zz_dataOut_payload_0_11888 <= _zz_dataOut_payload_0_11632;
    _zz_dataOut_payload_0_11889 <= _zz_dataOut_payload_0_11633;
    _zz_dataOut_payload_0_11890 <= _zz_dataOut_payload_0_11634;
    _zz_dataOut_payload_0_11891 <= _zz_dataOut_payload_0_11635;
    _zz_dataOut_payload_0_11892 <= _zz_dataOut_payload_0_11636;
    _zz_dataOut_payload_0_11893 <= _zz_dataOut_payload_0_11637;
    _zz_dataOut_payload_0_11894 <= _zz_dataOut_payload_0_11638;
    _zz_dataOut_payload_0_11895 <= _zz_dataOut_payload_0_11639;
    _zz_dataOut_payload_0_11896 <= _zz_dataOut_payload_0_11640;
    _zz_dataOut_payload_0_11897 <= _zz_dataOut_payload_0_11641;
    _zz_dataOut_payload_0_11898 <= _zz_dataOut_payload_0_11642;
    _zz_dataOut_payload_0_11899 <= _zz_dataOut_payload_0_11643;
    _zz_dataOut_payload_0_11900 <= _zz_dataOut_payload_0_11644;
    _zz_dataOut_payload_0_11901 <= _zz_dataOut_payload_0_11645;
    _zz_dataOut_payload_0_11902 <= _zz_dataOut_payload_0_11646;
    _zz_dataOut_payload_0_11903 <= _zz_dataOut_payload_0_11647;
    _zz_dataOut_payload_0_12284 <= (_zz_dataOut_payload_0_12282 ? _zz_dataOut_payload_0_12277 : _zz_dataOut_payload_0_12280);
    _zz_dataOut_payload_0_12285 <= (_zz_dataOut_payload_0_12282 ? _zz_dataOut_payload_0_12280 : _zz_dataOut_payload_0_12277);
    _zz_dataOut_payload_0_12286 <= (_zz_dataOut_payload_0_12283 ? _zz_dataOut_payload_0_12278 : _zz_dataOut_payload_0_12281);
    _zz_dataOut_payload_0_12287 <= (_zz_dataOut_payload_0_12283 ? _zz_dataOut_payload_0_12281 : _zz_dataOut_payload_0_12278);
    _zz_dataOut_payload_0_12296 <= (_zz_dataOut_payload_0_12294 ? _zz_dataOut_payload_0_12289 : _zz_dataOut_payload_0_12292);
    _zz_dataOut_payload_0_12297 <= (_zz_dataOut_payload_0_12294 ? _zz_dataOut_payload_0_12292 : _zz_dataOut_payload_0_12289);
    _zz_dataOut_payload_0_12298 <= (_zz_dataOut_payload_0_12295 ? _zz_dataOut_payload_0_12290 : _zz_dataOut_payload_0_12293);
    _zz_dataOut_payload_0_12299 <= (_zz_dataOut_payload_0_12295 ? _zz_dataOut_payload_0_12293 : _zz_dataOut_payload_0_12290);
    _zz_dataOut_payload_0_12300 <= _zz_dataOut_payload_0_12284;
    _zz_dataOut_payload_0_12301 <= _zz_dataOut_payload_0_12285;
    _zz_dataOut_payload_0_12302 <= _zz_dataOut_payload_0_12286;
    _zz_dataOut_payload_0_12303 <= _zz_dataOut_payload_0_12287;
    _zz_dataOut_payload_0_12304 <= _zz_dataOut_payload_0_12296;
    _zz_dataOut_payload_0_12305 <= _zz_dataOut_payload_0_12297;
    _zz_dataOut_payload_0_12306 <= _zz_dataOut_payload_0_12298;
    _zz_dataOut_payload_0_12307 <= _zz_dataOut_payload_0_12299;
    _zz_dataOut_payload_0_12328 <= (_zz_dataOut_payload_0_12326 ? _zz_dataOut_payload_0_12321 : _zz_dataOut_payload_0_12324);
    _zz_dataOut_payload_0_12329 <= (_zz_dataOut_payload_0_12326 ? _zz_dataOut_payload_0_12324 : _zz_dataOut_payload_0_12321);
    _zz_dataOut_payload_0_12330 <= (_zz_dataOut_payload_0_12327 ? _zz_dataOut_payload_0_12322 : _zz_dataOut_payload_0_12325);
    _zz_dataOut_payload_0_12331 <= (_zz_dataOut_payload_0_12327 ? _zz_dataOut_payload_0_12325 : _zz_dataOut_payload_0_12322);
    _zz_dataOut_payload_0_12340 <= (_zz_dataOut_payload_0_12338 ? _zz_dataOut_payload_0_12333 : _zz_dataOut_payload_0_12336);
    _zz_dataOut_payload_0_12341 <= (_zz_dataOut_payload_0_12338 ? _zz_dataOut_payload_0_12336 : _zz_dataOut_payload_0_12333);
    _zz_dataOut_payload_0_12342 <= (_zz_dataOut_payload_0_12339 ? _zz_dataOut_payload_0_12334 : _zz_dataOut_payload_0_12337);
    _zz_dataOut_payload_0_12343 <= (_zz_dataOut_payload_0_12339 ? _zz_dataOut_payload_0_12337 : _zz_dataOut_payload_0_12334);
    _zz_dataOut_payload_0_12344 <= _zz_dataOut_payload_0_12328;
    _zz_dataOut_payload_0_12345 <= _zz_dataOut_payload_0_12329;
    _zz_dataOut_payload_0_12346 <= _zz_dataOut_payload_0_12330;
    _zz_dataOut_payload_0_12347 <= _zz_dataOut_payload_0_12331;
    _zz_dataOut_payload_0_12348 <= _zz_dataOut_payload_0_12340;
    _zz_dataOut_payload_0_12349 <= _zz_dataOut_payload_0_12341;
    _zz_dataOut_payload_0_12350 <= _zz_dataOut_payload_0_12342;
    _zz_dataOut_payload_0_12351 <= _zz_dataOut_payload_0_12343;
    _zz_dataOut_payload_0_12352 <= _zz_dataOut_payload_0_12300;
    _zz_dataOut_payload_0_12353 <= _zz_dataOut_payload_0_12301;
    _zz_dataOut_payload_0_12354 <= _zz_dataOut_payload_0_12302;
    _zz_dataOut_payload_0_12355 <= _zz_dataOut_payload_0_12303;
    _zz_dataOut_payload_0_12356 <= _zz_dataOut_payload_0_12304;
    _zz_dataOut_payload_0_12357 <= _zz_dataOut_payload_0_12305;
    _zz_dataOut_payload_0_12358 <= _zz_dataOut_payload_0_12306;
    _zz_dataOut_payload_0_12359 <= _zz_dataOut_payload_0_12307;
    _zz_dataOut_payload_0_12360 <= _zz_dataOut_payload_0_12344;
    _zz_dataOut_payload_0_12361 <= _zz_dataOut_payload_0_12345;
    _zz_dataOut_payload_0_12362 <= _zz_dataOut_payload_0_12346;
    _zz_dataOut_payload_0_12363 <= _zz_dataOut_payload_0_12347;
    _zz_dataOut_payload_0_12364 <= _zz_dataOut_payload_0_12348;
    _zz_dataOut_payload_0_12365 <= _zz_dataOut_payload_0_12349;
    _zz_dataOut_payload_0_12366 <= _zz_dataOut_payload_0_12350;
    _zz_dataOut_payload_0_12367 <= _zz_dataOut_payload_0_12351;
    _zz_dataOut_payload_0_12412 <= (_zz_dataOut_payload_0_12410 ? _zz_dataOut_payload_0_12405 : _zz_dataOut_payload_0_12408);
    _zz_dataOut_payload_0_12413 <= (_zz_dataOut_payload_0_12410 ? _zz_dataOut_payload_0_12408 : _zz_dataOut_payload_0_12405);
    _zz_dataOut_payload_0_12414 <= (_zz_dataOut_payload_0_12411 ? _zz_dataOut_payload_0_12406 : _zz_dataOut_payload_0_12409);
    _zz_dataOut_payload_0_12415 <= (_zz_dataOut_payload_0_12411 ? _zz_dataOut_payload_0_12409 : _zz_dataOut_payload_0_12406);
    _zz_dataOut_payload_0_12424 <= (_zz_dataOut_payload_0_12422 ? _zz_dataOut_payload_0_12417 : _zz_dataOut_payload_0_12420);
    _zz_dataOut_payload_0_12425 <= (_zz_dataOut_payload_0_12422 ? _zz_dataOut_payload_0_12420 : _zz_dataOut_payload_0_12417);
    _zz_dataOut_payload_0_12426 <= (_zz_dataOut_payload_0_12423 ? _zz_dataOut_payload_0_12418 : _zz_dataOut_payload_0_12421);
    _zz_dataOut_payload_0_12427 <= (_zz_dataOut_payload_0_12423 ? _zz_dataOut_payload_0_12421 : _zz_dataOut_payload_0_12418);
    _zz_dataOut_payload_0_12428 <= _zz_dataOut_payload_0_12412;
    _zz_dataOut_payload_0_12429 <= _zz_dataOut_payload_0_12413;
    _zz_dataOut_payload_0_12430 <= _zz_dataOut_payload_0_12414;
    _zz_dataOut_payload_0_12431 <= _zz_dataOut_payload_0_12415;
    _zz_dataOut_payload_0_12432 <= _zz_dataOut_payload_0_12424;
    _zz_dataOut_payload_0_12433 <= _zz_dataOut_payload_0_12425;
    _zz_dataOut_payload_0_12434 <= _zz_dataOut_payload_0_12426;
    _zz_dataOut_payload_0_12435 <= _zz_dataOut_payload_0_12427;
    _zz_dataOut_payload_0_12456 <= (_zz_dataOut_payload_0_12454 ? _zz_dataOut_payload_0_12449 : _zz_dataOut_payload_0_12452);
    _zz_dataOut_payload_0_12457 <= (_zz_dataOut_payload_0_12454 ? _zz_dataOut_payload_0_12452 : _zz_dataOut_payload_0_12449);
    _zz_dataOut_payload_0_12458 <= (_zz_dataOut_payload_0_12455 ? _zz_dataOut_payload_0_12450 : _zz_dataOut_payload_0_12453);
    _zz_dataOut_payload_0_12459 <= (_zz_dataOut_payload_0_12455 ? _zz_dataOut_payload_0_12453 : _zz_dataOut_payload_0_12450);
    _zz_dataOut_payload_0_12468 <= (_zz_dataOut_payload_0_12466 ? _zz_dataOut_payload_0_12461 : _zz_dataOut_payload_0_12464);
    _zz_dataOut_payload_0_12469 <= (_zz_dataOut_payload_0_12466 ? _zz_dataOut_payload_0_12464 : _zz_dataOut_payload_0_12461);
    _zz_dataOut_payload_0_12470 <= (_zz_dataOut_payload_0_12467 ? _zz_dataOut_payload_0_12462 : _zz_dataOut_payload_0_12465);
    _zz_dataOut_payload_0_12471 <= (_zz_dataOut_payload_0_12467 ? _zz_dataOut_payload_0_12465 : _zz_dataOut_payload_0_12462);
    _zz_dataOut_payload_0_12472 <= _zz_dataOut_payload_0_12456;
    _zz_dataOut_payload_0_12473 <= _zz_dataOut_payload_0_12457;
    _zz_dataOut_payload_0_12474 <= _zz_dataOut_payload_0_12458;
    _zz_dataOut_payload_0_12475 <= _zz_dataOut_payload_0_12459;
    _zz_dataOut_payload_0_12476 <= _zz_dataOut_payload_0_12468;
    _zz_dataOut_payload_0_12477 <= _zz_dataOut_payload_0_12469;
    _zz_dataOut_payload_0_12478 <= _zz_dataOut_payload_0_12470;
    _zz_dataOut_payload_0_12479 <= _zz_dataOut_payload_0_12471;
    _zz_dataOut_payload_0_12480 <= _zz_dataOut_payload_0_12428;
    _zz_dataOut_payload_0_12481 <= _zz_dataOut_payload_0_12429;
    _zz_dataOut_payload_0_12482 <= _zz_dataOut_payload_0_12430;
    _zz_dataOut_payload_0_12483 <= _zz_dataOut_payload_0_12431;
    _zz_dataOut_payload_0_12484 <= _zz_dataOut_payload_0_12432;
    _zz_dataOut_payload_0_12485 <= _zz_dataOut_payload_0_12433;
    _zz_dataOut_payload_0_12486 <= _zz_dataOut_payload_0_12434;
    _zz_dataOut_payload_0_12487 <= _zz_dataOut_payload_0_12435;
    _zz_dataOut_payload_0_12488 <= _zz_dataOut_payload_0_12472;
    _zz_dataOut_payload_0_12489 <= _zz_dataOut_payload_0_12473;
    _zz_dataOut_payload_0_12490 <= _zz_dataOut_payload_0_12474;
    _zz_dataOut_payload_0_12491 <= _zz_dataOut_payload_0_12475;
    _zz_dataOut_payload_0_12492 <= _zz_dataOut_payload_0_12476;
    _zz_dataOut_payload_0_12493 <= _zz_dataOut_payload_0_12477;
    _zz_dataOut_payload_0_12494 <= _zz_dataOut_payload_0_12478;
    _zz_dataOut_payload_0_12495 <= _zz_dataOut_payload_0_12479;
    _zz_dataOut_payload_0_12496 <= _zz_dataOut_payload_0_12352;
    _zz_dataOut_payload_0_12497 <= _zz_dataOut_payload_0_12353;
    _zz_dataOut_payload_0_12498 <= _zz_dataOut_payload_0_12354;
    _zz_dataOut_payload_0_12499 <= _zz_dataOut_payload_0_12355;
    _zz_dataOut_payload_0_12500 <= _zz_dataOut_payload_0_12356;
    _zz_dataOut_payload_0_12501 <= _zz_dataOut_payload_0_12357;
    _zz_dataOut_payload_0_12502 <= _zz_dataOut_payload_0_12358;
    _zz_dataOut_payload_0_12503 <= _zz_dataOut_payload_0_12359;
    _zz_dataOut_payload_0_12504 <= _zz_dataOut_payload_0_12360;
    _zz_dataOut_payload_0_12505 <= _zz_dataOut_payload_0_12361;
    _zz_dataOut_payload_0_12506 <= _zz_dataOut_payload_0_12362;
    _zz_dataOut_payload_0_12507 <= _zz_dataOut_payload_0_12363;
    _zz_dataOut_payload_0_12508 <= _zz_dataOut_payload_0_12364;
    _zz_dataOut_payload_0_12509 <= _zz_dataOut_payload_0_12365;
    _zz_dataOut_payload_0_12510 <= _zz_dataOut_payload_0_12366;
    _zz_dataOut_payload_0_12511 <= _zz_dataOut_payload_0_12367;
    _zz_dataOut_payload_0_12512 <= _zz_dataOut_payload_0_12480;
    _zz_dataOut_payload_0_12513 <= _zz_dataOut_payload_0_12481;
    _zz_dataOut_payload_0_12514 <= _zz_dataOut_payload_0_12482;
    _zz_dataOut_payload_0_12515 <= _zz_dataOut_payload_0_12483;
    _zz_dataOut_payload_0_12516 <= _zz_dataOut_payload_0_12484;
    _zz_dataOut_payload_0_12517 <= _zz_dataOut_payload_0_12485;
    _zz_dataOut_payload_0_12518 <= _zz_dataOut_payload_0_12486;
    _zz_dataOut_payload_0_12519 <= _zz_dataOut_payload_0_12487;
    _zz_dataOut_payload_0_12520 <= _zz_dataOut_payload_0_12488;
    _zz_dataOut_payload_0_12521 <= _zz_dataOut_payload_0_12489;
    _zz_dataOut_payload_0_12522 <= _zz_dataOut_payload_0_12490;
    _zz_dataOut_payload_0_12523 <= _zz_dataOut_payload_0_12491;
    _zz_dataOut_payload_0_12524 <= _zz_dataOut_payload_0_12492;
    _zz_dataOut_payload_0_12525 <= _zz_dataOut_payload_0_12493;
    _zz_dataOut_payload_0_12526 <= _zz_dataOut_payload_0_12494;
    _zz_dataOut_payload_0_12527 <= _zz_dataOut_payload_0_12495;
    _zz_dataOut_payload_0_12620 <= (_zz_dataOut_payload_0_12618 ? _zz_dataOut_payload_0_12613 : _zz_dataOut_payload_0_12616);
    _zz_dataOut_payload_0_12621 <= (_zz_dataOut_payload_0_12618 ? _zz_dataOut_payload_0_12616 : _zz_dataOut_payload_0_12613);
    _zz_dataOut_payload_0_12622 <= (_zz_dataOut_payload_0_12619 ? _zz_dataOut_payload_0_12614 : _zz_dataOut_payload_0_12617);
    _zz_dataOut_payload_0_12623 <= (_zz_dataOut_payload_0_12619 ? _zz_dataOut_payload_0_12617 : _zz_dataOut_payload_0_12614);
    _zz_dataOut_payload_0_12632 <= (_zz_dataOut_payload_0_12630 ? _zz_dataOut_payload_0_12625 : _zz_dataOut_payload_0_12628);
    _zz_dataOut_payload_0_12633 <= (_zz_dataOut_payload_0_12630 ? _zz_dataOut_payload_0_12628 : _zz_dataOut_payload_0_12625);
    _zz_dataOut_payload_0_12634 <= (_zz_dataOut_payload_0_12631 ? _zz_dataOut_payload_0_12626 : _zz_dataOut_payload_0_12629);
    _zz_dataOut_payload_0_12635 <= (_zz_dataOut_payload_0_12631 ? _zz_dataOut_payload_0_12629 : _zz_dataOut_payload_0_12626);
    _zz_dataOut_payload_0_12636 <= _zz_dataOut_payload_0_12620;
    _zz_dataOut_payload_0_12637 <= _zz_dataOut_payload_0_12621;
    _zz_dataOut_payload_0_12638 <= _zz_dataOut_payload_0_12622;
    _zz_dataOut_payload_0_12639 <= _zz_dataOut_payload_0_12623;
    _zz_dataOut_payload_0_12640 <= _zz_dataOut_payload_0_12632;
    _zz_dataOut_payload_0_12641 <= _zz_dataOut_payload_0_12633;
    _zz_dataOut_payload_0_12642 <= _zz_dataOut_payload_0_12634;
    _zz_dataOut_payload_0_12643 <= _zz_dataOut_payload_0_12635;
    _zz_dataOut_payload_0_12664 <= (_zz_dataOut_payload_0_12662 ? _zz_dataOut_payload_0_12657 : _zz_dataOut_payload_0_12660);
    _zz_dataOut_payload_0_12665 <= (_zz_dataOut_payload_0_12662 ? _zz_dataOut_payload_0_12660 : _zz_dataOut_payload_0_12657);
    _zz_dataOut_payload_0_12666 <= (_zz_dataOut_payload_0_12663 ? _zz_dataOut_payload_0_12658 : _zz_dataOut_payload_0_12661);
    _zz_dataOut_payload_0_12667 <= (_zz_dataOut_payload_0_12663 ? _zz_dataOut_payload_0_12661 : _zz_dataOut_payload_0_12658);
    _zz_dataOut_payload_0_12676 <= (_zz_dataOut_payload_0_12674 ? _zz_dataOut_payload_0_12669 : _zz_dataOut_payload_0_12672);
    _zz_dataOut_payload_0_12677 <= (_zz_dataOut_payload_0_12674 ? _zz_dataOut_payload_0_12672 : _zz_dataOut_payload_0_12669);
    _zz_dataOut_payload_0_12678 <= (_zz_dataOut_payload_0_12675 ? _zz_dataOut_payload_0_12670 : _zz_dataOut_payload_0_12673);
    _zz_dataOut_payload_0_12679 <= (_zz_dataOut_payload_0_12675 ? _zz_dataOut_payload_0_12673 : _zz_dataOut_payload_0_12670);
    _zz_dataOut_payload_0_12680 <= _zz_dataOut_payload_0_12664;
    _zz_dataOut_payload_0_12681 <= _zz_dataOut_payload_0_12665;
    _zz_dataOut_payload_0_12682 <= _zz_dataOut_payload_0_12666;
    _zz_dataOut_payload_0_12683 <= _zz_dataOut_payload_0_12667;
    _zz_dataOut_payload_0_12684 <= _zz_dataOut_payload_0_12676;
    _zz_dataOut_payload_0_12685 <= _zz_dataOut_payload_0_12677;
    _zz_dataOut_payload_0_12686 <= _zz_dataOut_payload_0_12678;
    _zz_dataOut_payload_0_12687 <= _zz_dataOut_payload_0_12679;
    _zz_dataOut_payload_0_12688 <= _zz_dataOut_payload_0_12636;
    _zz_dataOut_payload_0_12689 <= _zz_dataOut_payload_0_12637;
    _zz_dataOut_payload_0_12690 <= _zz_dataOut_payload_0_12638;
    _zz_dataOut_payload_0_12691 <= _zz_dataOut_payload_0_12639;
    _zz_dataOut_payload_0_12692 <= _zz_dataOut_payload_0_12640;
    _zz_dataOut_payload_0_12693 <= _zz_dataOut_payload_0_12641;
    _zz_dataOut_payload_0_12694 <= _zz_dataOut_payload_0_12642;
    _zz_dataOut_payload_0_12695 <= _zz_dataOut_payload_0_12643;
    _zz_dataOut_payload_0_12696 <= _zz_dataOut_payload_0_12680;
    _zz_dataOut_payload_0_12697 <= _zz_dataOut_payload_0_12681;
    _zz_dataOut_payload_0_12698 <= _zz_dataOut_payload_0_12682;
    _zz_dataOut_payload_0_12699 <= _zz_dataOut_payload_0_12683;
    _zz_dataOut_payload_0_12700 <= _zz_dataOut_payload_0_12684;
    _zz_dataOut_payload_0_12701 <= _zz_dataOut_payload_0_12685;
    _zz_dataOut_payload_0_12702 <= _zz_dataOut_payload_0_12686;
    _zz_dataOut_payload_0_12703 <= _zz_dataOut_payload_0_12687;
    _zz_dataOut_payload_0_12748 <= (_zz_dataOut_payload_0_12746 ? _zz_dataOut_payload_0_12741 : _zz_dataOut_payload_0_12744);
    _zz_dataOut_payload_0_12749 <= (_zz_dataOut_payload_0_12746 ? _zz_dataOut_payload_0_12744 : _zz_dataOut_payload_0_12741);
    _zz_dataOut_payload_0_12750 <= (_zz_dataOut_payload_0_12747 ? _zz_dataOut_payload_0_12742 : _zz_dataOut_payload_0_12745);
    _zz_dataOut_payload_0_12751 <= (_zz_dataOut_payload_0_12747 ? _zz_dataOut_payload_0_12745 : _zz_dataOut_payload_0_12742);
    _zz_dataOut_payload_0_12760 <= (_zz_dataOut_payload_0_12758 ? _zz_dataOut_payload_0_12753 : _zz_dataOut_payload_0_12756);
    _zz_dataOut_payload_0_12761 <= (_zz_dataOut_payload_0_12758 ? _zz_dataOut_payload_0_12756 : _zz_dataOut_payload_0_12753);
    _zz_dataOut_payload_0_12762 <= (_zz_dataOut_payload_0_12759 ? _zz_dataOut_payload_0_12754 : _zz_dataOut_payload_0_12757);
    _zz_dataOut_payload_0_12763 <= (_zz_dataOut_payload_0_12759 ? _zz_dataOut_payload_0_12757 : _zz_dataOut_payload_0_12754);
    _zz_dataOut_payload_0_12764 <= _zz_dataOut_payload_0_12748;
    _zz_dataOut_payload_0_12765 <= _zz_dataOut_payload_0_12749;
    _zz_dataOut_payload_0_12766 <= _zz_dataOut_payload_0_12750;
    _zz_dataOut_payload_0_12767 <= _zz_dataOut_payload_0_12751;
    _zz_dataOut_payload_0_12768 <= _zz_dataOut_payload_0_12760;
    _zz_dataOut_payload_0_12769 <= _zz_dataOut_payload_0_12761;
    _zz_dataOut_payload_0_12770 <= _zz_dataOut_payload_0_12762;
    _zz_dataOut_payload_0_12771 <= _zz_dataOut_payload_0_12763;
    _zz_dataOut_payload_0_12792 <= (_zz_dataOut_payload_0_12790 ? _zz_dataOut_payload_0_12785 : _zz_dataOut_payload_0_12788);
    _zz_dataOut_payload_0_12793 <= (_zz_dataOut_payload_0_12790 ? _zz_dataOut_payload_0_12788 : _zz_dataOut_payload_0_12785);
    _zz_dataOut_payload_0_12794 <= (_zz_dataOut_payload_0_12791 ? _zz_dataOut_payload_0_12786 : _zz_dataOut_payload_0_12789);
    _zz_dataOut_payload_0_12795 <= (_zz_dataOut_payload_0_12791 ? _zz_dataOut_payload_0_12789 : _zz_dataOut_payload_0_12786);
    _zz_dataOut_payload_0_12804 <= (_zz_dataOut_payload_0_12802 ? _zz_dataOut_payload_0_12797 : _zz_dataOut_payload_0_12800);
    _zz_dataOut_payload_0_12805 <= (_zz_dataOut_payload_0_12802 ? _zz_dataOut_payload_0_12800 : _zz_dataOut_payload_0_12797);
    _zz_dataOut_payload_0_12806 <= (_zz_dataOut_payload_0_12803 ? _zz_dataOut_payload_0_12798 : _zz_dataOut_payload_0_12801);
    _zz_dataOut_payload_0_12807 <= (_zz_dataOut_payload_0_12803 ? _zz_dataOut_payload_0_12801 : _zz_dataOut_payload_0_12798);
    _zz_dataOut_payload_0_12808 <= _zz_dataOut_payload_0_12792;
    _zz_dataOut_payload_0_12809 <= _zz_dataOut_payload_0_12793;
    _zz_dataOut_payload_0_12810 <= _zz_dataOut_payload_0_12794;
    _zz_dataOut_payload_0_12811 <= _zz_dataOut_payload_0_12795;
    _zz_dataOut_payload_0_12812 <= _zz_dataOut_payload_0_12804;
    _zz_dataOut_payload_0_12813 <= _zz_dataOut_payload_0_12805;
    _zz_dataOut_payload_0_12814 <= _zz_dataOut_payload_0_12806;
    _zz_dataOut_payload_0_12815 <= _zz_dataOut_payload_0_12807;
    _zz_dataOut_payload_0_12816 <= _zz_dataOut_payload_0_12764;
    _zz_dataOut_payload_0_12817 <= _zz_dataOut_payload_0_12765;
    _zz_dataOut_payload_0_12818 <= _zz_dataOut_payload_0_12766;
    _zz_dataOut_payload_0_12819 <= _zz_dataOut_payload_0_12767;
    _zz_dataOut_payload_0_12820 <= _zz_dataOut_payload_0_12768;
    _zz_dataOut_payload_0_12821 <= _zz_dataOut_payload_0_12769;
    _zz_dataOut_payload_0_12822 <= _zz_dataOut_payload_0_12770;
    _zz_dataOut_payload_0_12823 <= _zz_dataOut_payload_0_12771;
    _zz_dataOut_payload_0_12824 <= _zz_dataOut_payload_0_12808;
    _zz_dataOut_payload_0_12825 <= _zz_dataOut_payload_0_12809;
    _zz_dataOut_payload_0_12826 <= _zz_dataOut_payload_0_12810;
    _zz_dataOut_payload_0_12827 <= _zz_dataOut_payload_0_12811;
    _zz_dataOut_payload_0_12828 <= _zz_dataOut_payload_0_12812;
    _zz_dataOut_payload_0_12829 <= _zz_dataOut_payload_0_12813;
    _zz_dataOut_payload_0_12830 <= _zz_dataOut_payload_0_12814;
    _zz_dataOut_payload_0_12831 <= _zz_dataOut_payload_0_12815;
    _zz_dataOut_payload_0_12832 <= _zz_dataOut_payload_0_12688;
    _zz_dataOut_payload_0_12833 <= _zz_dataOut_payload_0_12689;
    _zz_dataOut_payload_0_12834 <= _zz_dataOut_payload_0_12690;
    _zz_dataOut_payload_0_12835 <= _zz_dataOut_payload_0_12691;
    _zz_dataOut_payload_0_12836 <= _zz_dataOut_payload_0_12692;
    _zz_dataOut_payload_0_12837 <= _zz_dataOut_payload_0_12693;
    _zz_dataOut_payload_0_12838 <= _zz_dataOut_payload_0_12694;
    _zz_dataOut_payload_0_12839 <= _zz_dataOut_payload_0_12695;
    _zz_dataOut_payload_0_12840 <= _zz_dataOut_payload_0_12696;
    _zz_dataOut_payload_0_12841 <= _zz_dataOut_payload_0_12697;
    _zz_dataOut_payload_0_12842 <= _zz_dataOut_payload_0_12698;
    _zz_dataOut_payload_0_12843 <= _zz_dataOut_payload_0_12699;
    _zz_dataOut_payload_0_12844 <= _zz_dataOut_payload_0_12700;
    _zz_dataOut_payload_0_12845 <= _zz_dataOut_payload_0_12701;
    _zz_dataOut_payload_0_12846 <= _zz_dataOut_payload_0_12702;
    _zz_dataOut_payload_0_12847 <= _zz_dataOut_payload_0_12703;
    _zz_dataOut_payload_0_12848 <= _zz_dataOut_payload_0_12816;
    _zz_dataOut_payload_0_12849 <= _zz_dataOut_payload_0_12817;
    _zz_dataOut_payload_0_12850 <= _zz_dataOut_payload_0_12818;
    _zz_dataOut_payload_0_12851 <= _zz_dataOut_payload_0_12819;
    _zz_dataOut_payload_0_12852 <= _zz_dataOut_payload_0_12820;
    _zz_dataOut_payload_0_12853 <= _zz_dataOut_payload_0_12821;
    _zz_dataOut_payload_0_12854 <= _zz_dataOut_payload_0_12822;
    _zz_dataOut_payload_0_12855 <= _zz_dataOut_payload_0_12823;
    _zz_dataOut_payload_0_12856 <= _zz_dataOut_payload_0_12824;
    _zz_dataOut_payload_0_12857 <= _zz_dataOut_payload_0_12825;
    _zz_dataOut_payload_0_12858 <= _zz_dataOut_payload_0_12826;
    _zz_dataOut_payload_0_12859 <= _zz_dataOut_payload_0_12827;
    _zz_dataOut_payload_0_12860 <= _zz_dataOut_payload_0_12828;
    _zz_dataOut_payload_0_12861 <= _zz_dataOut_payload_0_12829;
    _zz_dataOut_payload_0_12862 <= _zz_dataOut_payload_0_12830;
    _zz_dataOut_payload_0_12863 <= _zz_dataOut_payload_0_12831;
    _zz_dataOut_payload_0_12864 <= _zz_dataOut_payload_0_12496;
    _zz_dataOut_payload_0_12865 <= _zz_dataOut_payload_0_12497;
    _zz_dataOut_payload_0_12866 <= _zz_dataOut_payload_0_12498;
    _zz_dataOut_payload_0_12867 <= _zz_dataOut_payload_0_12499;
    _zz_dataOut_payload_0_12868 <= _zz_dataOut_payload_0_12500;
    _zz_dataOut_payload_0_12869 <= _zz_dataOut_payload_0_12501;
    _zz_dataOut_payload_0_12870 <= _zz_dataOut_payload_0_12502;
    _zz_dataOut_payload_0_12871 <= _zz_dataOut_payload_0_12503;
    _zz_dataOut_payload_0_12872 <= _zz_dataOut_payload_0_12504;
    _zz_dataOut_payload_0_12873 <= _zz_dataOut_payload_0_12505;
    _zz_dataOut_payload_0_12874 <= _zz_dataOut_payload_0_12506;
    _zz_dataOut_payload_0_12875 <= _zz_dataOut_payload_0_12507;
    _zz_dataOut_payload_0_12876 <= _zz_dataOut_payload_0_12508;
    _zz_dataOut_payload_0_12877 <= _zz_dataOut_payload_0_12509;
    _zz_dataOut_payload_0_12878 <= _zz_dataOut_payload_0_12510;
    _zz_dataOut_payload_0_12879 <= _zz_dataOut_payload_0_12511;
    _zz_dataOut_payload_0_12880 <= _zz_dataOut_payload_0_12512;
    _zz_dataOut_payload_0_12881 <= _zz_dataOut_payload_0_12513;
    _zz_dataOut_payload_0_12882 <= _zz_dataOut_payload_0_12514;
    _zz_dataOut_payload_0_12883 <= _zz_dataOut_payload_0_12515;
    _zz_dataOut_payload_0_12884 <= _zz_dataOut_payload_0_12516;
    _zz_dataOut_payload_0_12885 <= _zz_dataOut_payload_0_12517;
    _zz_dataOut_payload_0_12886 <= _zz_dataOut_payload_0_12518;
    _zz_dataOut_payload_0_12887 <= _zz_dataOut_payload_0_12519;
    _zz_dataOut_payload_0_12888 <= _zz_dataOut_payload_0_12520;
    _zz_dataOut_payload_0_12889 <= _zz_dataOut_payload_0_12521;
    _zz_dataOut_payload_0_12890 <= _zz_dataOut_payload_0_12522;
    _zz_dataOut_payload_0_12891 <= _zz_dataOut_payload_0_12523;
    _zz_dataOut_payload_0_12892 <= _zz_dataOut_payload_0_12524;
    _zz_dataOut_payload_0_12893 <= _zz_dataOut_payload_0_12525;
    _zz_dataOut_payload_0_12894 <= _zz_dataOut_payload_0_12526;
    _zz_dataOut_payload_0_12895 <= _zz_dataOut_payload_0_12527;
    _zz_dataOut_payload_0_12896 <= _zz_dataOut_payload_0_12832;
    _zz_dataOut_payload_0_12897 <= _zz_dataOut_payload_0_12833;
    _zz_dataOut_payload_0_12898 <= _zz_dataOut_payload_0_12834;
    _zz_dataOut_payload_0_12899 <= _zz_dataOut_payload_0_12835;
    _zz_dataOut_payload_0_12900 <= _zz_dataOut_payload_0_12836;
    _zz_dataOut_payload_0_12901 <= _zz_dataOut_payload_0_12837;
    _zz_dataOut_payload_0_12902 <= _zz_dataOut_payload_0_12838;
    _zz_dataOut_payload_0_12903 <= _zz_dataOut_payload_0_12839;
    _zz_dataOut_payload_0_12904 <= _zz_dataOut_payload_0_12840;
    _zz_dataOut_payload_0_12905 <= _zz_dataOut_payload_0_12841;
    _zz_dataOut_payload_0_12906 <= _zz_dataOut_payload_0_12842;
    _zz_dataOut_payload_0_12907 <= _zz_dataOut_payload_0_12843;
    _zz_dataOut_payload_0_12908 <= _zz_dataOut_payload_0_12844;
    _zz_dataOut_payload_0_12909 <= _zz_dataOut_payload_0_12845;
    _zz_dataOut_payload_0_12910 <= _zz_dataOut_payload_0_12846;
    _zz_dataOut_payload_0_12911 <= _zz_dataOut_payload_0_12847;
    _zz_dataOut_payload_0_12912 <= _zz_dataOut_payload_0_12848;
    _zz_dataOut_payload_0_12913 <= _zz_dataOut_payload_0_12849;
    _zz_dataOut_payload_0_12914 <= _zz_dataOut_payload_0_12850;
    _zz_dataOut_payload_0_12915 <= _zz_dataOut_payload_0_12851;
    _zz_dataOut_payload_0_12916 <= _zz_dataOut_payload_0_12852;
    _zz_dataOut_payload_0_12917 <= _zz_dataOut_payload_0_12853;
    _zz_dataOut_payload_0_12918 <= _zz_dataOut_payload_0_12854;
    _zz_dataOut_payload_0_12919 <= _zz_dataOut_payload_0_12855;
    _zz_dataOut_payload_0_12920 <= _zz_dataOut_payload_0_12856;
    _zz_dataOut_payload_0_12921 <= _zz_dataOut_payload_0_12857;
    _zz_dataOut_payload_0_12922 <= _zz_dataOut_payload_0_12858;
    _zz_dataOut_payload_0_12923 <= _zz_dataOut_payload_0_12859;
    _zz_dataOut_payload_0_12924 <= _zz_dataOut_payload_0_12860;
    _zz_dataOut_payload_0_12925 <= _zz_dataOut_payload_0_12861;
    _zz_dataOut_payload_0_12926 <= _zz_dataOut_payload_0_12862;
    _zz_dataOut_payload_0_12927 <= _zz_dataOut_payload_0_12863;
    _zz_dataOut_payload_0_13116 <= (_zz_dataOut_payload_0_13114 ? _zz_dataOut_payload_0_13109 : _zz_dataOut_payload_0_13112);
    _zz_dataOut_payload_0_13117 <= (_zz_dataOut_payload_0_13114 ? _zz_dataOut_payload_0_13112 : _zz_dataOut_payload_0_13109);
    _zz_dataOut_payload_0_13118 <= (_zz_dataOut_payload_0_13115 ? _zz_dataOut_payload_0_13110 : _zz_dataOut_payload_0_13113);
    _zz_dataOut_payload_0_13119 <= (_zz_dataOut_payload_0_13115 ? _zz_dataOut_payload_0_13113 : _zz_dataOut_payload_0_13110);
    _zz_dataOut_payload_0_13128 <= (_zz_dataOut_payload_0_13126 ? _zz_dataOut_payload_0_13121 : _zz_dataOut_payload_0_13124);
    _zz_dataOut_payload_0_13129 <= (_zz_dataOut_payload_0_13126 ? _zz_dataOut_payload_0_13124 : _zz_dataOut_payload_0_13121);
    _zz_dataOut_payload_0_13130 <= (_zz_dataOut_payload_0_13127 ? _zz_dataOut_payload_0_13122 : _zz_dataOut_payload_0_13125);
    _zz_dataOut_payload_0_13131 <= (_zz_dataOut_payload_0_13127 ? _zz_dataOut_payload_0_13125 : _zz_dataOut_payload_0_13122);
    _zz_dataOut_payload_0_13132 <= _zz_dataOut_payload_0_13116;
    _zz_dataOut_payload_0_13133 <= _zz_dataOut_payload_0_13117;
    _zz_dataOut_payload_0_13134 <= _zz_dataOut_payload_0_13118;
    _zz_dataOut_payload_0_13135 <= _zz_dataOut_payload_0_13119;
    _zz_dataOut_payload_0_13136 <= _zz_dataOut_payload_0_13128;
    _zz_dataOut_payload_0_13137 <= _zz_dataOut_payload_0_13129;
    _zz_dataOut_payload_0_13138 <= _zz_dataOut_payload_0_13130;
    _zz_dataOut_payload_0_13139 <= _zz_dataOut_payload_0_13131;
    _zz_dataOut_payload_0_13160 <= (_zz_dataOut_payload_0_13158 ? _zz_dataOut_payload_0_13153 : _zz_dataOut_payload_0_13156);
    _zz_dataOut_payload_0_13161 <= (_zz_dataOut_payload_0_13158 ? _zz_dataOut_payload_0_13156 : _zz_dataOut_payload_0_13153);
    _zz_dataOut_payload_0_13162 <= (_zz_dataOut_payload_0_13159 ? _zz_dataOut_payload_0_13154 : _zz_dataOut_payload_0_13157);
    _zz_dataOut_payload_0_13163 <= (_zz_dataOut_payload_0_13159 ? _zz_dataOut_payload_0_13157 : _zz_dataOut_payload_0_13154);
    _zz_dataOut_payload_0_13172 <= (_zz_dataOut_payload_0_13170 ? _zz_dataOut_payload_0_13165 : _zz_dataOut_payload_0_13168);
    _zz_dataOut_payload_0_13173 <= (_zz_dataOut_payload_0_13170 ? _zz_dataOut_payload_0_13168 : _zz_dataOut_payload_0_13165);
    _zz_dataOut_payload_0_13174 <= (_zz_dataOut_payload_0_13171 ? _zz_dataOut_payload_0_13166 : _zz_dataOut_payload_0_13169);
    _zz_dataOut_payload_0_13175 <= (_zz_dataOut_payload_0_13171 ? _zz_dataOut_payload_0_13169 : _zz_dataOut_payload_0_13166);
    _zz_dataOut_payload_0_13176 <= _zz_dataOut_payload_0_13160;
    _zz_dataOut_payload_0_13177 <= _zz_dataOut_payload_0_13161;
    _zz_dataOut_payload_0_13178 <= _zz_dataOut_payload_0_13162;
    _zz_dataOut_payload_0_13179 <= _zz_dataOut_payload_0_13163;
    _zz_dataOut_payload_0_13180 <= _zz_dataOut_payload_0_13172;
    _zz_dataOut_payload_0_13181 <= _zz_dataOut_payload_0_13173;
    _zz_dataOut_payload_0_13182 <= _zz_dataOut_payload_0_13174;
    _zz_dataOut_payload_0_13183 <= _zz_dataOut_payload_0_13175;
    _zz_dataOut_payload_0_13184 <= _zz_dataOut_payload_0_13132;
    _zz_dataOut_payload_0_13185 <= _zz_dataOut_payload_0_13133;
    _zz_dataOut_payload_0_13186 <= _zz_dataOut_payload_0_13134;
    _zz_dataOut_payload_0_13187 <= _zz_dataOut_payload_0_13135;
    _zz_dataOut_payload_0_13188 <= _zz_dataOut_payload_0_13136;
    _zz_dataOut_payload_0_13189 <= _zz_dataOut_payload_0_13137;
    _zz_dataOut_payload_0_13190 <= _zz_dataOut_payload_0_13138;
    _zz_dataOut_payload_0_13191 <= _zz_dataOut_payload_0_13139;
    _zz_dataOut_payload_0_13192 <= _zz_dataOut_payload_0_13176;
    _zz_dataOut_payload_0_13193 <= _zz_dataOut_payload_0_13177;
    _zz_dataOut_payload_0_13194 <= _zz_dataOut_payload_0_13178;
    _zz_dataOut_payload_0_13195 <= _zz_dataOut_payload_0_13179;
    _zz_dataOut_payload_0_13196 <= _zz_dataOut_payload_0_13180;
    _zz_dataOut_payload_0_13197 <= _zz_dataOut_payload_0_13181;
    _zz_dataOut_payload_0_13198 <= _zz_dataOut_payload_0_13182;
    _zz_dataOut_payload_0_13199 <= _zz_dataOut_payload_0_13183;
    _zz_dataOut_payload_0_13244 <= (_zz_dataOut_payload_0_13242 ? _zz_dataOut_payload_0_13237 : _zz_dataOut_payload_0_13240);
    _zz_dataOut_payload_0_13245 <= (_zz_dataOut_payload_0_13242 ? _zz_dataOut_payload_0_13240 : _zz_dataOut_payload_0_13237);
    _zz_dataOut_payload_0_13246 <= (_zz_dataOut_payload_0_13243 ? _zz_dataOut_payload_0_13238 : _zz_dataOut_payload_0_13241);
    _zz_dataOut_payload_0_13247 <= (_zz_dataOut_payload_0_13243 ? _zz_dataOut_payload_0_13241 : _zz_dataOut_payload_0_13238);
    _zz_dataOut_payload_0_13256 <= (_zz_dataOut_payload_0_13254 ? _zz_dataOut_payload_0_13249 : _zz_dataOut_payload_0_13252);
    _zz_dataOut_payload_0_13257 <= (_zz_dataOut_payload_0_13254 ? _zz_dataOut_payload_0_13252 : _zz_dataOut_payload_0_13249);
    _zz_dataOut_payload_0_13258 <= (_zz_dataOut_payload_0_13255 ? _zz_dataOut_payload_0_13250 : _zz_dataOut_payload_0_13253);
    _zz_dataOut_payload_0_13259 <= (_zz_dataOut_payload_0_13255 ? _zz_dataOut_payload_0_13253 : _zz_dataOut_payload_0_13250);
    _zz_dataOut_payload_0_13260 <= _zz_dataOut_payload_0_13244;
    _zz_dataOut_payload_0_13261 <= _zz_dataOut_payload_0_13245;
    _zz_dataOut_payload_0_13262 <= _zz_dataOut_payload_0_13246;
    _zz_dataOut_payload_0_13263 <= _zz_dataOut_payload_0_13247;
    _zz_dataOut_payload_0_13264 <= _zz_dataOut_payload_0_13256;
    _zz_dataOut_payload_0_13265 <= _zz_dataOut_payload_0_13257;
    _zz_dataOut_payload_0_13266 <= _zz_dataOut_payload_0_13258;
    _zz_dataOut_payload_0_13267 <= _zz_dataOut_payload_0_13259;
    _zz_dataOut_payload_0_13288 <= (_zz_dataOut_payload_0_13286 ? _zz_dataOut_payload_0_13281 : _zz_dataOut_payload_0_13284);
    _zz_dataOut_payload_0_13289 <= (_zz_dataOut_payload_0_13286 ? _zz_dataOut_payload_0_13284 : _zz_dataOut_payload_0_13281);
    _zz_dataOut_payload_0_13290 <= (_zz_dataOut_payload_0_13287 ? _zz_dataOut_payload_0_13282 : _zz_dataOut_payload_0_13285);
    _zz_dataOut_payload_0_13291 <= (_zz_dataOut_payload_0_13287 ? _zz_dataOut_payload_0_13285 : _zz_dataOut_payload_0_13282);
    _zz_dataOut_payload_0_13300 <= (_zz_dataOut_payload_0_13298 ? _zz_dataOut_payload_0_13293 : _zz_dataOut_payload_0_13296);
    _zz_dataOut_payload_0_13301 <= (_zz_dataOut_payload_0_13298 ? _zz_dataOut_payload_0_13296 : _zz_dataOut_payload_0_13293);
    _zz_dataOut_payload_0_13302 <= (_zz_dataOut_payload_0_13299 ? _zz_dataOut_payload_0_13294 : _zz_dataOut_payload_0_13297);
    _zz_dataOut_payload_0_13303 <= (_zz_dataOut_payload_0_13299 ? _zz_dataOut_payload_0_13297 : _zz_dataOut_payload_0_13294);
    _zz_dataOut_payload_0_13304 <= _zz_dataOut_payload_0_13288;
    _zz_dataOut_payload_0_13305 <= _zz_dataOut_payload_0_13289;
    _zz_dataOut_payload_0_13306 <= _zz_dataOut_payload_0_13290;
    _zz_dataOut_payload_0_13307 <= _zz_dataOut_payload_0_13291;
    _zz_dataOut_payload_0_13308 <= _zz_dataOut_payload_0_13300;
    _zz_dataOut_payload_0_13309 <= _zz_dataOut_payload_0_13301;
    _zz_dataOut_payload_0_13310 <= _zz_dataOut_payload_0_13302;
    _zz_dataOut_payload_0_13311 <= _zz_dataOut_payload_0_13303;
    _zz_dataOut_payload_0_13312 <= _zz_dataOut_payload_0_13260;
    _zz_dataOut_payload_0_13313 <= _zz_dataOut_payload_0_13261;
    _zz_dataOut_payload_0_13314 <= _zz_dataOut_payload_0_13262;
    _zz_dataOut_payload_0_13315 <= _zz_dataOut_payload_0_13263;
    _zz_dataOut_payload_0_13316 <= _zz_dataOut_payload_0_13264;
    _zz_dataOut_payload_0_13317 <= _zz_dataOut_payload_0_13265;
    _zz_dataOut_payload_0_13318 <= _zz_dataOut_payload_0_13266;
    _zz_dataOut_payload_0_13319 <= _zz_dataOut_payload_0_13267;
    _zz_dataOut_payload_0_13320 <= _zz_dataOut_payload_0_13304;
    _zz_dataOut_payload_0_13321 <= _zz_dataOut_payload_0_13305;
    _zz_dataOut_payload_0_13322 <= _zz_dataOut_payload_0_13306;
    _zz_dataOut_payload_0_13323 <= _zz_dataOut_payload_0_13307;
    _zz_dataOut_payload_0_13324 <= _zz_dataOut_payload_0_13308;
    _zz_dataOut_payload_0_13325 <= _zz_dataOut_payload_0_13309;
    _zz_dataOut_payload_0_13326 <= _zz_dataOut_payload_0_13310;
    _zz_dataOut_payload_0_13327 <= _zz_dataOut_payload_0_13311;
    _zz_dataOut_payload_0_13328 <= _zz_dataOut_payload_0_13184;
    _zz_dataOut_payload_0_13329 <= _zz_dataOut_payload_0_13185;
    _zz_dataOut_payload_0_13330 <= _zz_dataOut_payload_0_13186;
    _zz_dataOut_payload_0_13331 <= _zz_dataOut_payload_0_13187;
    _zz_dataOut_payload_0_13332 <= _zz_dataOut_payload_0_13188;
    _zz_dataOut_payload_0_13333 <= _zz_dataOut_payload_0_13189;
    _zz_dataOut_payload_0_13334 <= _zz_dataOut_payload_0_13190;
    _zz_dataOut_payload_0_13335 <= _zz_dataOut_payload_0_13191;
    _zz_dataOut_payload_0_13336 <= _zz_dataOut_payload_0_13192;
    _zz_dataOut_payload_0_13337 <= _zz_dataOut_payload_0_13193;
    _zz_dataOut_payload_0_13338 <= _zz_dataOut_payload_0_13194;
    _zz_dataOut_payload_0_13339 <= _zz_dataOut_payload_0_13195;
    _zz_dataOut_payload_0_13340 <= _zz_dataOut_payload_0_13196;
    _zz_dataOut_payload_0_13341 <= _zz_dataOut_payload_0_13197;
    _zz_dataOut_payload_0_13342 <= _zz_dataOut_payload_0_13198;
    _zz_dataOut_payload_0_13343 <= _zz_dataOut_payload_0_13199;
    _zz_dataOut_payload_0_13344 <= _zz_dataOut_payload_0_13312;
    _zz_dataOut_payload_0_13345 <= _zz_dataOut_payload_0_13313;
    _zz_dataOut_payload_0_13346 <= _zz_dataOut_payload_0_13314;
    _zz_dataOut_payload_0_13347 <= _zz_dataOut_payload_0_13315;
    _zz_dataOut_payload_0_13348 <= _zz_dataOut_payload_0_13316;
    _zz_dataOut_payload_0_13349 <= _zz_dataOut_payload_0_13317;
    _zz_dataOut_payload_0_13350 <= _zz_dataOut_payload_0_13318;
    _zz_dataOut_payload_0_13351 <= _zz_dataOut_payload_0_13319;
    _zz_dataOut_payload_0_13352 <= _zz_dataOut_payload_0_13320;
    _zz_dataOut_payload_0_13353 <= _zz_dataOut_payload_0_13321;
    _zz_dataOut_payload_0_13354 <= _zz_dataOut_payload_0_13322;
    _zz_dataOut_payload_0_13355 <= _zz_dataOut_payload_0_13323;
    _zz_dataOut_payload_0_13356 <= _zz_dataOut_payload_0_13324;
    _zz_dataOut_payload_0_13357 <= _zz_dataOut_payload_0_13325;
    _zz_dataOut_payload_0_13358 <= _zz_dataOut_payload_0_13326;
    _zz_dataOut_payload_0_13359 <= _zz_dataOut_payload_0_13327;
    _zz_dataOut_payload_0_13452 <= (_zz_dataOut_payload_0_13450 ? _zz_dataOut_payload_0_13445 : _zz_dataOut_payload_0_13448);
    _zz_dataOut_payload_0_13453 <= (_zz_dataOut_payload_0_13450 ? _zz_dataOut_payload_0_13448 : _zz_dataOut_payload_0_13445);
    _zz_dataOut_payload_0_13454 <= (_zz_dataOut_payload_0_13451 ? _zz_dataOut_payload_0_13446 : _zz_dataOut_payload_0_13449);
    _zz_dataOut_payload_0_13455 <= (_zz_dataOut_payload_0_13451 ? _zz_dataOut_payload_0_13449 : _zz_dataOut_payload_0_13446);
    _zz_dataOut_payload_0_13464 <= (_zz_dataOut_payload_0_13462 ? _zz_dataOut_payload_0_13457 : _zz_dataOut_payload_0_13460);
    _zz_dataOut_payload_0_13465 <= (_zz_dataOut_payload_0_13462 ? _zz_dataOut_payload_0_13460 : _zz_dataOut_payload_0_13457);
    _zz_dataOut_payload_0_13466 <= (_zz_dataOut_payload_0_13463 ? _zz_dataOut_payload_0_13458 : _zz_dataOut_payload_0_13461);
    _zz_dataOut_payload_0_13467 <= (_zz_dataOut_payload_0_13463 ? _zz_dataOut_payload_0_13461 : _zz_dataOut_payload_0_13458);
    _zz_dataOut_payload_0_13468 <= _zz_dataOut_payload_0_13452;
    _zz_dataOut_payload_0_13469 <= _zz_dataOut_payload_0_13453;
    _zz_dataOut_payload_0_13470 <= _zz_dataOut_payload_0_13454;
    _zz_dataOut_payload_0_13471 <= _zz_dataOut_payload_0_13455;
    _zz_dataOut_payload_0_13472 <= _zz_dataOut_payload_0_13464;
    _zz_dataOut_payload_0_13473 <= _zz_dataOut_payload_0_13465;
    _zz_dataOut_payload_0_13474 <= _zz_dataOut_payload_0_13466;
    _zz_dataOut_payload_0_13475 <= _zz_dataOut_payload_0_13467;
    _zz_dataOut_payload_0_13496 <= (_zz_dataOut_payload_0_13494 ? _zz_dataOut_payload_0_13489 : _zz_dataOut_payload_0_13492);
    _zz_dataOut_payload_0_13497 <= (_zz_dataOut_payload_0_13494 ? _zz_dataOut_payload_0_13492 : _zz_dataOut_payload_0_13489);
    _zz_dataOut_payload_0_13498 <= (_zz_dataOut_payload_0_13495 ? _zz_dataOut_payload_0_13490 : _zz_dataOut_payload_0_13493);
    _zz_dataOut_payload_0_13499 <= (_zz_dataOut_payload_0_13495 ? _zz_dataOut_payload_0_13493 : _zz_dataOut_payload_0_13490);
    _zz_dataOut_payload_0_13508 <= (_zz_dataOut_payload_0_13506 ? _zz_dataOut_payload_0_13501 : _zz_dataOut_payload_0_13504);
    _zz_dataOut_payload_0_13509 <= (_zz_dataOut_payload_0_13506 ? _zz_dataOut_payload_0_13504 : _zz_dataOut_payload_0_13501);
    _zz_dataOut_payload_0_13510 <= (_zz_dataOut_payload_0_13507 ? _zz_dataOut_payload_0_13502 : _zz_dataOut_payload_0_13505);
    _zz_dataOut_payload_0_13511 <= (_zz_dataOut_payload_0_13507 ? _zz_dataOut_payload_0_13505 : _zz_dataOut_payload_0_13502);
    _zz_dataOut_payload_0_13512 <= _zz_dataOut_payload_0_13496;
    _zz_dataOut_payload_0_13513 <= _zz_dataOut_payload_0_13497;
    _zz_dataOut_payload_0_13514 <= _zz_dataOut_payload_0_13498;
    _zz_dataOut_payload_0_13515 <= _zz_dataOut_payload_0_13499;
    _zz_dataOut_payload_0_13516 <= _zz_dataOut_payload_0_13508;
    _zz_dataOut_payload_0_13517 <= _zz_dataOut_payload_0_13509;
    _zz_dataOut_payload_0_13518 <= _zz_dataOut_payload_0_13510;
    _zz_dataOut_payload_0_13519 <= _zz_dataOut_payload_0_13511;
    _zz_dataOut_payload_0_13520 <= _zz_dataOut_payload_0_13468;
    _zz_dataOut_payload_0_13521 <= _zz_dataOut_payload_0_13469;
    _zz_dataOut_payload_0_13522 <= _zz_dataOut_payload_0_13470;
    _zz_dataOut_payload_0_13523 <= _zz_dataOut_payload_0_13471;
    _zz_dataOut_payload_0_13524 <= _zz_dataOut_payload_0_13472;
    _zz_dataOut_payload_0_13525 <= _zz_dataOut_payload_0_13473;
    _zz_dataOut_payload_0_13526 <= _zz_dataOut_payload_0_13474;
    _zz_dataOut_payload_0_13527 <= _zz_dataOut_payload_0_13475;
    _zz_dataOut_payload_0_13528 <= _zz_dataOut_payload_0_13512;
    _zz_dataOut_payload_0_13529 <= _zz_dataOut_payload_0_13513;
    _zz_dataOut_payload_0_13530 <= _zz_dataOut_payload_0_13514;
    _zz_dataOut_payload_0_13531 <= _zz_dataOut_payload_0_13515;
    _zz_dataOut_payload_0_13532 <= _zz_dataOut_payload_0_13516;
    _zz_dataOut_payload_0_13533 <= _zz_dataOut_payload_0_13517;
    _zz_dataOut_payload_0_13534 <= _zz_dataOut_payload_0_13518;
    _zz_dataOut_payload_0_13535 <= _zz_dataOut_payload_0_13519;
    _zz_dataOut_payload_0_13580 <= (_zz_dataOut_payload_0_13578 ? _zz_dataOut_payload_0_13573 : _zz_dataOut_payload_0_13576);
    _zz_dataOut_payload_0_13581 <= (_zz_dataOut_payload_0_13578 ? _zz_dataOut_payload_0_13576 : _zz_dataOut_payload_0_13573);
    _zz_dataOut_payload_0_13582 <= (_zz_dataOut_payload_0_13579 ? _zz_dataOut_payload_0_13574 : _zz_dataOut_payload_0_13577);
    _zz_dataOut_payload_0_13583 <= (_zz_dataOut_payload_0_13579 ? _zz_dataOut_payload_0_13577 : _zz_dataOut_payload_0_13574);
    _zz_dataOut_payload_0_13592 <= (_zz_dataOut_payload_0_13590 ? _zz_dataOut_payload_0_13585 : _zz_dataOut_payload_0_13588);
    _zz_dataOut_payload_0_13593 <= (_zz_dataOut_payload_0_13590 ? _zz_dataOut_payload_0_13588 : _zz_dataOut_payload_0_13585);
    _zz_dataOut_payload_0_13594 <= (_zz_dataOut_payload_0_13591 ? _zz_dataOut_payload_0_13586 : _zz_dataOut_payload_0_13589);
    _zz_dataOut_payload_0_13595 <= (_zz_dataOut_payload_0_13591 ? _zz_dataOut_payload_0_13589 : _zz_dataOut_payload_0_13586);
    _zz_dataOut_payload_0_13596 <= _zz_dataOut_payload_0_13580;
    _zz_dataOut_payload_0_13597 <= _zz_dataOut_payload_0_13581;
    _zz_dataOut_payload_0_13598 <= _zz_dataOut_payload_0_13582;
    _zz_dataOut_payload_0_13599 <= _zz_dataOut_payload_0_13583;
    _zz_dataOut_payload_0_13600 <= _zz_dataOut_payload_0_13592;
    _zz_dataOut_payload_0_13601 <= _zz_dataOut_payload_0_13593;
    _zz_dataOut_payload_0_13602 <= _zz_dataOut_payload_0_13594;
    _zz_dataOut_payload_0_13603 <= _zz_dataOut_payload_0_13595;
    _zz_dataOut_payload_0_13624 <= (_zz_dataOut_payload_0_13622 ? _zz_dataOut_payload_0_13617 : _zz_dataOut_payload_0_13620);
    _zz_dataOut_payload_0_13625 <= (_zz_dataOut_payload_0_13622 ? _zz_dataOut_payload_0_13620 : _zz_dataOut_payload_0_13617);
    _zz_dataOut_payload_0_13626 <= (_zz_dataOut_payload_0_13623 ? _zz_dataOut_payload_0_13618 : _zz_dataOut_payload_0_13621);
    _zz_dataOut_payload_0_13627 <= (_zz_dataOut_payload_0_13623 ? _zz_dataOut_payload_0_13621 : _zz_dataOut_payload_0_13618);
    _zz_dataOut_payload_0_13636 <= (_zz_dataOut_payload_0_13634 ? _zz_dataOut_payload_0_13629 : _zz_dataOut_payload_0_13632);
    _zz_dataOut_payload_0_13637 <= (_zz_dataOut_payload_0_13634 ? _zz_dataOut_payload_0_13632 : _zz_dataOut_payload_0_13629);
    _zz_dataOut_payload_0_13638 <= (_zz_dataOut_payload_0_13635 ? _zz_dataOut_payload_0_13630 : _zz_dataOut_payload_0_13633);
    _zz_dataOut_payload_0_13639 <= (_zz_dataOut_payload_0_13635 ? _zz_dataOut_payload_0_13633 : _zz_dataOut_payload_0_13630);
    _zz_dataOut_payload_0_13640 <= _zz_dataOut_payload_0_13624;
    _zz_dataOut_payload_0_13641 <= _zz_dataOut_payload_0_13625;
    _zz_dataOut_payload_0_13642 <= _zz_dataOut_payload_0_13626;
    _zz_dataOut_payload_0_13643 <= _zz_dataOut_payload_0_13627;
    _zz_dataOut_payload_0_13644 <= _zz_dataOut_payload_0_13636;
    _zz_dataOut_payload_0_13645 <= _zz_dataOut_payload_0_13637;
    _zz_dataOut_payload_0_13646 <= _zz_dataOut_payload_0_13638;
    _zz_dataOut_payload_0_13647 <= _zz_dataOut_payload_0_13639;
    _zz_dataOut_payload_0_13648 <= _zz_dataOut_payload_0_13596;
    _zz_dataOut_payload_0_13649 <= _zz_dataOut_payload_0_13597;
    _zz_dataOut_payload_0_13650 <= _zz_dataOut_payload_0_13598;
    _zz_dataOut_payload_0_13651 <= _zz_dataOut_payload_0_13599;
    _zz_dataOut_payload_0_13652 <= _zz_dataOut_payload_0_13600;
    _zz_dataOut_payload_0_13653 <= _zz_dataOut_payload_0_13601;
    _zz_dataOut_payload_0_13654 <= _zz_dataOut_payload_0_13602;
    _zz_dataOut_payload_0_13655 <= _zz_dataOut_payload_0_13603;
    _zz_dataOut_payload_0_13656 <= _zz_dataOut_payload_0_13640;
    _zz_dataOut_payload_0_13657 <= _zz_dataOut_payload_0_13641;
    _zz_dataOut_payload_0_13658 <= _zz_dataOut_payload_0_13642;
    _zz_dataOut_payload_0_13659 <= _zz_dataOut_payload_0_13643;
    _zz_dataOut_payload_0_13660 <= _zz_dataOut_payload_0_13644;
    _zz_dataOut_payload_0_13661 <= _zz_dataOut_payload_0_13645;
    _zz_dataOut_payload_0_13662 <= _zz_dataOut_payload_0_13646;
    _zz_dataOut_payload_0_13663 <= _zz_dataOut_payload_0_13647;
    _zz_dataOut_payload_0_13664 <= _zz_dataOut_payload_0_13520;
    _zz_dataOut_payload_0_13665 <= _zz_dataOut_payload_0_13521;
    _zz_dataOut_payload_0_13666 <= _zz_dataOut_payload_0_13522;
    _zz_dataOut_payload_0_13667 <= _zz_dataOut_payload_0_13523;
    _zz_dataOut_payload_0_13668 <= _zz_dataOut_payload_0_13524;
    _zz_dataOut_payload_0_13669 <= _zz_dataOut_payload_0_13525;
    _zz_dataOut_payload_0_13670 <= _zz_dataOut_payload_0_13526;
    _zz_dataOut_payload_0_13671 <= _zz_dataOut_payload_0_13527;
    _zz_dataOut_payload_0_13672 <= _zz_dataOut_payload_0_13528;
    _zz_dataOut_payload_0_13673 <= _zz_dataOut_payload_0_13529;
    _zz_dataOut_payload_0_13674 <= _zz_dataOut_payload_0_13530;
    _zz_dataOut_payload_0_13675 <= _zz_dataOut_payload_0_13531;
    _zz_dataOut_payload_0_13676 <= _zz_dataOut_payload_0_13532;
    _zz_dataOut_payload_0_13677 <= _zz_dataOut_payload_0_13533;
    _zz_dataOut_payload_0_13678 <= _zz_dataOut_payload_0_13534;
    _zz_dataOut_payload_0_13679 <= _zz_dataOut_payload_0_13535;
    _zz_dataOut_payload_0_13680 <= _zz_dataOut_payload_0_13648;
    _zz_dataOut_payload_0_13681 <= _zz_dataOut_payload_0_13649;
    _zz_dataOut_payload_0_13682 <= _zz_dataOut_payload_0_13650;
    _zz_dataOut_payload_0_13683 <= _zz_dataOut_payload_0_13651;
    _zz_dataOut_payload_0_13684 <= _zz_dataOut_payload_0_13652;
    _zz_dataOut_payload_0_13685 <= _zz_dataOut_payload_0_13653;
    _zz_dataOut_payload_0_13686 <= _zz_dataOut_payload_0_13654;
    _zz_dataOut_payload_0_13687 <= _zz_dataOut_payload_0_13655;
    _zz_dataOut_payload_0_13688 <= _zz_dataOut_payload_0_13656;
    _zz_dataOut_payload_0_13689 <= _zz_dataOut_payload_0_13657;
    _zz_dataOut_payload_0_13690 <= _zz_dataOut_payload_0_13658;
    _zz_dataOut_payload_0_13691 <= _zz_dataOut_payload_0_13659;
    _zz_dataOut_payload_0_13692 <= _zz_dataOut_payload_0_13660;
    _zz_dataOut_payload_0_13693 <= _zz_dataOut_payload_0_13661;
    _zz_dataOut_payload_0_13694 <= _zz_dataOut_payload_0_13662;
    _zz_dataOut_payload_0_13695 <= _zz_dataOut_payload_0_13663;
    _zz_dataOut_payload_0_13696 <= _zz_dataOut_payload_0_13328;
    _zz_dataOut_payload_0_13697 <= _zz_dataOut_payload_0_13329;
    _zz_dataOut_payload_0_13698 <= _zz_dataOut_payload_0_13330;
    _zz_dataOut_payload_0_13699 <= _zz_dataOut_payload_0_13331;
    _zz_dataOut_payload_0_13700 <= _zz_dataOut_payload_0_13332;
    _zz_dataOut_payload_0_13701 <= _zz_dataOut_payload_0_13333;
    _zz_dataOut_payload_0_13702 <= _zz_dataOut_payload_0_13334;
    _zz_dataOut_payload_0_13703 <= _zz_dataOut_payload_0_13335;
    _zz_dataOut_payload_0_13704 <= _zz_dataOut_payload_0_13336;
    _zz_dataOut_payload_0_13705 <= _zz_dataOut_payload_0_13337;
    _zz_dataOut_payload_0_13706 <= _zz_dataOut_payload_0_13338;
    _zz_dataOut_payload_0_13707 <= _zz_dataOut_payload_0_13339;
    _zz_dataOut_payload_0_13708 <= _zz_dataOut_payload_0_13340;
    _zz_dataOut_payload_0_13709 <= _zz_dataOut_payload_0_13341;
    _zz_dataOut_payload_0_13710 <= _zz_dataOut_payload_0_13342;
    _zz_dataOut_payload_0_13711 <= _zz_dataOut_payload_0_13343;
    _zz_dataOut_payload_0_13712 <= _zz_dataOut_payload_0_13344;
    _zz_dataOut_payload_0_13713 <= _zz_dataOut_payload_0_13345;
    _zz_dataOut_payload_0_13714 <= _zz_dataOut_payload_0_13346;
    _zz_dataOut_payload_0_13715 <= _zz_dataOut_payload_0_13347;
    _zz_dataOut_payload_0_13716 <= _zz_dataOut_payload_0_13348;
    _zz_dataOut_payload_0_13717 <= _zz_dataOut_payload_0_13349;
    _zz_dataOut_payload_0_13718 <= _zz_dataOut_payload_0_13350;
    _zz_dataOut_payload_0_13719 <= _zz_dataOut_payload_0_13351;
    _zz_dataOut_payload_0_13720 <= _zz_dataOut_payload_0_13352;
    _zz_dataOut_payload_0_13721 <= _zz_dataOut_payload_0_13353;
    _zz_dataOut_payload_0_13722 <= _zz_dataOut_payload_0_13354;
    _zz_dataOut_payload_0_13723 <= _zz_dataOut_payload_0_13355;
    _zz_dataOut_payload_0_13724 <= _zz_dataOut_payload_0_13356;
    _zz_dataOut_payload_0_13725 <= _zz_dataOut_payload_0_13357;
    _zz_dataOut_payload_0_13726 <= _zz_dataOut_payload_0_13358;
    _zz_dataOut_payload_0_13727 <= _zz_dataOut_payload_0_13359;
    _zz_dataOut_payload_0_13728 <= _zz_dataOut_payload_0_13664;
    _zz_dataOut_payload_0_13729 <= _zz_dataOut_payload_0_13665;
    _zz_dataOut_payload_0_13730 <= _zz_dataOut_payload_0_13666;
    _zz_dataOut_payload_0_13731 <= _zz_dataOut_payload_0_13667;
    _zz_dataOut_payload_0_13732 <= _zz_dataOut_payload_0_13668;
    _zz_dataOut_payload_0_13733 <= _zz_dataOut_payload_0_13669;
    _zz_dataOut_payload_0_13734 <= _zz_dataOut_payload_0_13670;
    _zz_dataOut_payload_0_13735 <= _zz_dataOut_payload_0_13671;
    _zz_dataOut_payload_0_13736 <= _zz_dataOut_payload_0_13672;
    _zz_dataOut_payload_0_13737 <= _zz_dataOut_payload_0_13673;
    _zz_dataOut_payload_0_13738 <= _zz_dataOut_payload_0_13674;
    _zz_dataOut_payload_0_13739 <= _zz_dataOut_payload_0_13675;
    _zz_dataOut_payload_0_13740 <= _zz_dataOut_payload_0_13676;
    _zz_dataOut_payload_0_13741 <= _zz_dataOut_payload_0_13677;
    _zz_dataOut_payload_0_13742 <= _zz_dataOut_payload_0_13678;
    _zz_dataOut_payload_0_13743 <= _zz_dataOut_payload_0_13679;
    _zz_dataOut_payload_0_13744 <= _zz_dataOut_payload_0_13680;
    _zz_dataOut_payload_0_13745 <= _zz_dataOut_payload_0_13681;
    _zz_dataOut_payload_0_13746 <= _zz_dataOut_payload_0_13682;
    _zz_dataOut_payload_0_13747 <= _zz_dataOut_payload_0_13683;
    _zz_dataOut_payload_0_13748 <= _zz_dataOut_payload_0_13684;
    _zz_dataOut_payload_0_13749 <= _zz_dataOut_payload_0_13685;
    _zz_dataOut_payload_0_13750 <= _zz_dataOut_payload_0_13686;
    _zz_dataOut_payload_0_13751 <= _zz_dataOut_payload_0_13687;
    _zz_dataOut_payload_0_13752 <= _zz_dataOut_payload_0_13688;
    _zz_dataOut_payload_0_13753 <= _zz_dataOut_payload_0_13689;
    _zz_dataOut_payload_0_13754 <= _zz_dataOut_payload_0_13690;
    _zz_dataOut_payload_0_13755 <= _zz_dataOut_payload_0_13691;
    _zz_dataOut_payload_0_13756 <= _zz_dataOut_payload_0_13692;
    _zz_dataOut_payload_0_13757 <= _zz_dataOut_payload_0_13693;
    _zz_dataOut_payload_0_13758 <= _zz_dataOut_payload_0_13694;
    _zz_dataOut_payload_0_13759 <= _zz_dataOut_payload_0_13695;
    _zz_dataOut_payload_0_13760 <= _zz_dataOut_payload_0_12864;
    _zz_dataOut_payload_0_13761 <= _zz_dataOut_payload_0_12865;
    _zz_dataOut_payload_0_13762 <= _zz_dataOut_payload_0_12866;
    _zz_dataOut_payload_0_13763 <= _zz_dataOut_payload_0_12867;
    _zz_dataOut_payload_0_13764 <= _zz_dataOut_payload_0_12868;
    _zz_dataOut_payload_0_13765 <= _zz_dataOut_payload_0_12869;
    _zz_dataOut_payload_0_13766 <= _zz_dataOut_payload_0_12870;
    _zz_dataOut_payload_0_13767 <= _zz_dataOut_payload_0_12871;
    _zz_dataOut_payload_0_13768 <= _zz_dataOut_payload_0_12872;
    _zz_dataOut_payload_0_13769 <= _zz_dataOut_payload_0_12873;
    _zz_dataOut_payload_0_13770 <= _zz_dataOut_payload_0_12874;
    _zz_dataOut_payload_0_13771 <= _zz_dataOut_payload_0_12875;
    _zz_dataOut_payload_0_13772 <= _zz_dataOut_payload_0_12876;
    _zz_dataOut_payload_0_13773 <= _zz_dataOut_payload_0_12877;
    _zz_dataOut_payload_0_13774 <= _zz_dataOut_payload_0_12878;
    _zz_dataOut_payload_0_13775 <= _zz_dataOut_payload_0_12879;
    _zz_dataOut_payload_0_13776 <= _zz_dataOut_payload_0_12880;
    _zz_dataOut_payload_0_13777 <= _zz_dataOut_payload_0_12881;
    _zz_dataOut_payload_0_13778 <= _zz_dataOut_payload_0_12882;
    _zz_dataOut_payload_0_13779 <= _zz_dataOut_payload_0_12883;
    _zz_dataOut_payload_0_13780 <= _zz_dataOut_payload_0_12884;
    _zz_dataOut_payload_0_13781 <= _zz_dataOut_payload_0_12885;
    _zz_dataOut_payload_0_13782 <= _zz_dataOut_payload_0_12886;
    _zz_dataOut_payload_0_13783 <= _zz_dataOut_payload_0_12887;
    _zz_dataOut_payload_0_13784 <= _zz_dataOut_payload_0_12888;
    _zz_dataOut_payload_0_13785 <= _zz_dataOut_payload_0_12889;
    _zz_dataOut_payload_0_13786 <= _zz_dataOut_payload_0_12890;
    _zz_dataOut_payload_0_13787 <= _zz_dataOut_payload_0_12891;
    _zz_dataOut_payload_0_13788 <= _zz_dataOut_payload_0_12892;
    _zz_dataOut_payload_0_13789 <= _zz_dataOut_payload_0_12893;
    _zz_dataOut_payload_0_13790 <= _zz_dataOut_payload_0_12894;
    _zz_dataOut_payload_0_13791 <= _zz_dataOut_payload_0_12895;
    _zz_dataOut_payload_0_13792 <= _zz_dataOut_payload_0_12896;
    _zz_dataOut_payload_0_13793 <= _zz_dataOut_payload_0_12897;
    _zz_dataOut_payload_0_13794 <= _zz_dataOut_payload_0_12898;
    _zz_dataOut_payload_0_13795 <= _zz_dataOut_payload_0_12899;
    _zz_dataOut_payload_0_13796 <= _zz_dataOut_payload_0_12900;
    _zz_dataOut_payload_0_13797 <= _zz_dataOut_payload_0_12901;
    _zz_dataOut_payload_0_13798 <= _zz_dataOut_payload_0_12902;
    _zz_dataOut_payload_0_13799 <= _zz_dataOut_payload_0_12903;
    _zz_dataOut_payload_0_13800 <= _zz_dataOut_payload_0_12904;
    _zz_dataOut_payload_0_13801 <= _zz_dataOut_payload_0_12905;
    _zz_dataOut_payload_0_13802 <= _zz_dataOut_payload_0_12906;
    _zz_dataOut_payload_0_13803 <= _zz_dataOut_payload_0_12907;
    _zz_dataOut_payload_0_13804 <= _zz_dataOut_payload_0_12908;
    _zz_dataOut_payload_0_13805 <= _zz_dataOut_payload_0_12909;
    _zz_dataOut_payload_0_13806 <= _zz_dataOut_payload_0_12910;
    _zz_dataOut_payload_0_13807 <= _zz_dataOut_payload_0_12911;
    _zz_dataOut_payload_0_13808 <= _zz_dataOut_payload_0_12912;
    _zz_dataOut_payload_0_13809 <= _zz_dataOut_payload_0_12913;
    _zz_dataOut_payload_0_13810 <= _zz_dataOut_payload_0_12914;
    _zz_dataOut_payload_0_13811 <= _zz_dataOut_payload_0_12915;
    _zz_dataOut_payload_0_13812 <= _zz_dataOut_payload_0_12916;
    _zz_dataOut_payload_0_13813 <= _zz_dataOut_payload_0_12917;
    _zz_dataOut_payload_0_13814 <= _zz_dataOut_payload_0_12918;
    _zz_dataOut_payload_0_13815 <= _zz_dataOut_payload_0_12919;
    _zz_dataOut_payload_0_13816 <= _zz_dataOut_payload_0_12920;
    _zz_dataOut_payload_0_13817 <= _zz_dataOut_payload_0_12921;
    _zz_dataOut_payload_0_13818 <= _zz_dataOut_payload_0_12922;
    _zz_dataOut_payload_0_13819 <= _zz_dataOut_payload_0_12923;
    _zz_dataOut_payload_0_13820 <= _zz_dataOut_payload_0_12924;
    _zz_dataOut_payload_0_13821 <= _zz_dataOut_payload_0_12925;
    _zz_dataOut_payload_0_13822 <= _zz_dataOut_payload_0_12926;
    _zz_dataOut_payload_0_13823 <= _zz_dataOut_payload_0_12927;
    _zz_dataOut_payload_0_13824 <= _zz_dataOut_payload_0_13696;
    _zz_dataOut_payload_0_13825 <= _zz_dataOut_payload_0_13697;
    _zz_dataOut_payload_0_13826 <= _zz_dataOut_payload_0_13698;
    _zz_dataOut_payload_0_13827 <= _zz_dataOut_payload_0_13699;
    _zz_dataOut_payload_0_13828 <= _zz_dataOut_payload_0_13700;
    _zz_dataOut_payload_0_13829 <= _zz_dataOut_payload_0_13701;
    _zz_dataOut_payload_0_13830 <= _zz_dataOut_payload_0_13702;
    _zz_dataOut_payload_0_13831 <= _zz_dataOut_payload_0_13703;
    _zz_dataOut_payload_0_13832 <= _zz_dataOut_payload_0_13704;
    _zz_dataOut_payload_0_13833 <= _zz_dataOut_payload_0_13705;
    _zz_dataOut_payload_0_13834 <= _zz_dataOut_payload_0_13706;
    _zz_dataOut_payload_0_13835 <= _zz_dataOut_payload_0_13707;
    _zz_dataOut_payload_0_13836 <= _zz_dataOut_payload_0_13708;
    _zz_dataOut_payload_0_13837 <= _zz_dataOut_payload_0_13709;
    _zz_dataOut_payload_0_13838 <= _zz_dataOut_payload_0_13710;
    _zz_dataOut_payload_0_13839 <= _zz_dataOut_payload_0_13711;
    _zz_dataOut_payload_0_13840 <= _zz_dataOut_payload_0_13712;
    _zz_dataOut_payload_0_13841 <= _zz_dataOut_payload_0_13713;
    _zz_dataOut_payload_0_13842 <= _zz_dataOut_payload_0_13714;
    _zz_dataOut_payload_0_13843 <= _zz_dataOut_payload_0_13715;
    _zz_dataOut_payload_0_13844 <= _zz_dataOut_payload_0_13716;
    _zz_dataOut_payload_0_13845 <= _zz_dataOut_payload_0_13717;
    _zz_dataOut_payload_0_13846 <= _zz_dataOut_payload_0_13718;
    _zz_dataOut_payload_0_13847 <= _zz_dataOut_payload_0_13719;
    _zz_dataOut_payload_0_13848 <= _zz_dataOut_payload_0_13720;
    _zz_dataOut_payload_0_13849 <= _zz_dataOut_payload_0_13721;
    _zz_dataOut_payload_0_13850 <= _zz_dataOut_payload_0_13722;
    _zz_dataOut_payload_0_13851 <= _zz_dataOut_payload_0_13723;
    _zz_dataOut_payload_0_13852 <= _zz_dataOut_payload_0_13724;
    _zz_dataOut_payload_0_13853 <= _zz_dataOut_payload_0_13725;
    _zz_dataOut_payload_0_13854 <= _zz_dataOut_payload_0_13726;
    _zz_dataOut_payload_0_13855 <= _zz_dataOut_payload_0_13727;
    _zz_dataOut_payload_0_13856 <= _zz_dataOut_payload_0_13728;
    _zz_dataOut_payload_0_13857 <= _zz_dataOut_payload_0_13729;
    _zz_dataOut_payload_0_13858 <= _zz_dataOut_payload_0_13730;
    _zz_dataOut_payload_0_13859 <= _zz_dataOut_payload_0_13731;
    _zz_dataOut_payload_0_13860 <= _zz_dataOut_payload_0_13732;
    _zz_dataOut_payload_0_13861 <= _zz_dataOut_payload_0_13733;
    _zz_dataOut_payload_0_13862 <= _zz_dataOut_payload_0_13734;
    _zz_dataOut_payload_0_13863 <= _zz_dataOut_payload_0_13735;
    _zz_dataOut_payload_0_13864 <= _zz_dataOut_payload_0_13736;
    _zz_dataOut_payload_0_13865 <= _zz_dataOut_payload_0_13737;
    _zz_dataOut_payload_0_13866 <= _zz_dataOut_payload_0_13738;
    _zz_dataOut_payload_0_13867 <= _zz_dataOut_payload_0_13739;
    _zz_dataOut_payload_0_13868 <= _zz_dataOut_payload_0_13740;
    _zz_dataOut_payload_0_13869 <= _zz_dataOut_payload_0_13741;
    _zz_dataOut_payload_0_13870 <= _zz_dataOut_payload_0_13742;
    _zz_dataOut_payload_0_13871 <= _zz_dataOut_payload_0_13743;
    _zz_dataOut_payload_0_13872 <= _zz_dataOut_payload_0_13744;
    _zz_dataOut_payload_0_13873 <= _zz_dataOut_payload_0_13745;
    _zz_dataOut_payload_0_13874 <= _zz_dataOut_payload_0_13746;
    _zz_dataOut_payload_0_13875 <= _zz_dataOut_payload_0_13747;
    _zz_dataOut_payload_0_13876 <= _zz_dataOut_payload_0_13748;
    _zz_dataOut_payload_0_13877 <= _zz_dataOut_payload_0_13749;
    _zz_dataOut_payload_0_13878 <= _zz_dataOut_payload_0_13750;
    _zz_dataOut_payload_0_13879 <= _zz_dataOut_payload_0_13751;
    _zz_dataOut_payload_0_13880 <= _zz_dataOut_payload_0_13752;
    _zz_dataOut_payload_0_13881 <= _zz_dataOut_payload_0_13753;
    _zz_dataOut_payload_0_13882 <= _zz_dataOut_payload_0_13754;
    _zz_dataOut_payload_0_13883 <= _zz_dataOut_payload_0_13755;
    _zz_dataOut_payload_0_13884 <= _zz_dataOut_payload_0_13756;
    _zz_dataOut_payload_0_13885 <= _zz_dataOut_payload_0_13757;
    _zz_dataOut_payload_0_13886 <= _zz_dataOut_payload_0_13758;
    _zz_dataOut_payload_0_13887 <= _zz_dataOut_payload_0_13759;
    _zz_dataOut_payload_0_14268 <= (_zz_dataOut_payload_0_14266 ? _zz_dataOut_payload_0_14261 : _zz_dataOut_payload_0_14264);
    _zz_dataOut_payload_0_14269 <= (_zz_dataOut_payload_0_14266 ? _zz_dataOut_payload_0_14264 : _zz_dataOut_payload_0_14261);
    _zz_dataOut_payload_0_14270 <= (_zz_dataOut_payload_0_14267 ? _zz_dataOut_payload_0_14262 : _zz_dataOut_payload_0_14265);
    _zz_dataOut_payload_0_14271 <= (_zz_dataOut_payload_0_14267 ? _zz_dataOut_payload_0_14265 : _zz_dataOut_payload_0_14262);
    _zz_dataOut_payload_0_14280 <= (_zz_dataOut_payload_0_14278 ? _zz_dataOut_payload_0_14273 : _zz_dataOut_payload_0_14276);
    _zz_dataOut_payload_0_14281 <= (_zz_dataOut_payload_0_14278 ? _zz_dataOut_payload_0_14276 : _zz_dataOut_payload_0_14273);
    _zz_dataOut_payload_0_14282 <= (_zz_dataOut_payload_0_14279 ? _zz_dataOut_payload_0_14274 : _zz_dataOut_payload_0_14277);
    _zz_dataOut_payload_0_14283 <= (_zz_dataOut_payload_0_14279 ? _zz_dataOut_payload_0_14277 : _zz_dataOut_payload_0_14274);
    _zz_dataOut_payload_0_14284 <= _zz_dataOut_payload_0_14268;
    _zz_dataOut_payload_0_14285 <= _zz_dataOut_payload_0_14269;
    _zz_dataOut_payload_0_14286 <= _zz_dataOut_payload_0_14270;
    _zz_dataOut_payload_0_14287 <= _zz_dataOut_payload_0_14271;
    _zz_dataOut_payload_0_14288 <= _zz_dataOut_payload_0_14280;
    _zz_dataOut_payload_0_14289 <= _zz_dataOut_payload_0_14281;
    _zz_dataOut_payload_0_14290 <= _zz_dataOut_payload_0_14282;
    _zz_dataOut_payload_0_14291 <= _zz_dataOut_payload_0_14283;
    _zz_dataOut_payload_0_14312 <= (_zz_dataOut_payload_0_14310 ? _zz_dataOut_payload_0_14305 : _zz_dataOut_payload_0_14308);
    _zz_dataOut_payload_0_14313 <= (_zz_dataOut_payload_0_14310 ? _zz_dataOut_payload_0_14308 : _zz_dataOut_payload_0_14305);
    _zz_dataOut_payload_0_14314 <= (_zz_dataOut_payload_0_14311 ? _zz_dataOut_payload_0_14306 : _zz_dataOut_payload_0_14309);
    _zz_dataOut_payload_0_14315 <= (_zz_dataOut_payload_0_14311 ? _zz_dataOut_payload_0_14309 : _zz_dataOut_payload_0_14306);
    _zz_dataOut_payload_0_14324 <= (_zz_dataOut_payload_0_14322 ? _zz_dataOut_payload_0_14317 : _zz_dataOut_payload_0_14320);
    _zz_dataOut_payload_0_14325 <= (_zz_dataOut_payload_0_14322 ? _zz_dataOut_payload_0_14320 : _zz_dataOut_payload_0_14317);
    _zz_dataOut_payload_0_14326 <= (_zz_dataOut_payload_0_14323 ? _zz_dataOut_payload_0_14318 : _zz_dataOut_payload_0_14321);
    _zz_dataOut_payload_0_14327 <= (_zz_dataOut_payload_0_14323 ? _zz_dataOut_payload_0_14321 : _zz_dataOut_payload_0_14318);
    _zz_dataOut_payload_0_14328 <= _zz_dataOut_payload_0_14312;
    _zz_dataOut_payload_0_14329 <= _zz_dataOut_payload_0_14313;
    _zz_dataOut_payload_0_14330 <= _zz_dataOut_payload_0_14314;
    _zz_dataOut_payload_0_14331 <= _zz_dataOut_payload_0_14315;
    _zz_dataOut_payload_0_14332 <= _zz_dataOut_payload_0_14324;
    _zz_dataOut_payload_0_14333 <= _zz_dataOut_payload_0_14325;
    _zz_dataOut_payload_0_14334 <= _zz_dataOut_payload_0_14326;
    _zz_dataOut_payload_0_14335 <= _zz_dataOut_payload_0_14327;
    _zz_dataOut_payload_0_14336 <= _zz_dataOut_payload_0_14284;
    _zz_dataOut_payload_0_14337 <= _zz_dataOut_payload_0_14285;
    _zz_dataOut_payload_0_14338 <= _zz_dataOut_payload_0_14286;
    _zz_dataOut_payload_0_14339 <= _zz_dataOut_payload_0_14287;
    _zz_dataOut_payload_0_14340 <= _zz_dataOut_payload_0_14288;
    _zz_dataOut_payload_0_14341 <= _zz_dataOut_payload_0_14289;
    _zz_dataOut_payload_0_14342 <= _zz_dataOut_payload_0_14290;
    _zz_dataOut_payload_0_14343 <= _zz_dataOut_payload_0_14291;
    _zz_dataOut_payload_0_14344 <= _zz_dataOut_payload_0_14328;
    _zz_dataOut_payload_0_14345 <= _zz_dataOut_payload_0_14329;
    _zz_dataOut_payload_0_14346 <= _zz_dataOut_payload_0_14330;
    _zz_dataOut_payload_0_14347 <= _zz_dataOut_payload_0_14331;
    _zz_dataOut_payload_0_14348 <= _zz_dataOut_payload_0_14332;
    _zz_dataOut_payload_0_14349 <= _zz_dataOut_payload_0_14333;
    _zz_dataOut_payload_0_14350 <= _zz_dataOut_payload_0_14334;
    _zz_dataOut_payload_0_14351 <= _zz_dataOut_payload_0_14335;
    _zz_dataOut_payload_0_14396 <= (_zz_dataOut_payload_0_14394 ? _zz_dataOut_payload_0_14389 : _zz_dataOut_payload_0_14392);
    _zz_dataOut_payload_0_14397 <= (_zz_dataOut_payload_0_14394 ? _zz_dataOut_payload_0_14392 : _zz_dataOut_payload_0_14389);
    _zz_dataOut_payload_0_14398 <= (_zz_dataOut_payload_0_14395 ? _zz_dataOut_payload_0_14390 : _zz_dataOut_payload_0_14393);
    _zz_dataOut_payload_0_14399 <= (_zz_dataOut_payload_0_14395 ? _zz_dataOut_payload_0_14393 : _zz_dataOut_payload_0_14390);
    _zz_dataOut_payload_0_14408 <= (_zz_dataOut_payload_0_14406 ? _zz_dataOut_payload_0_14401 : _zz_dataOut_payload_0_14404);
    _zz_dataOut_payload_0_14409 <= (_zz_dataOut_payload_0_14406 ? _zz_dataOut_payload_0_14404 : _zz_dataOut_payload_0_14401);
    _zz_dataOut_payload_0_14410 <= (_zz_dataOut_payload_0_14407 ? _zz_dataOut_payload_0_14402 : _zz_dataOut_payload_0_14405);
    _zz_dataOut_payload_0_14411 <= (_zz_dataOut_payload_0_14407 ? _zz_dataOut_payload_0_14405 : _zz_dataOut_payload_0_14402);
    _zz_dataOut_payload_0_14412 <= _zz_dataOut_payload_0_14396;
    _zz_dataOut_payload_0_14413 <= _zz_dataOut_payload_0_14397;
    _zz_dataOut_payload_0_14414 <= _zz_dataOut_payload_0_14398;
    _zz_dataOut_payload_0_14415 <= _zz_dataOut_payload_0_14399;
    _zz_dataOut_payload_0_14416 <= _zz_dataOut_payload_0_14408;
    _zz_dataOut_payload_0_14417 <= _zz_dataOut_payload_0_14409;
    _zz_dataOut_payload_0_14418 <= _zz_dataOut_payload_0_14410;
    _zz_dataOut_payload_0_14419 <= _zz_dataOut_payload_0_14411;
    _zz_dataOut_payload_0_14440 <= (_zz_dataOut_payload_0_14438 ? _zz_dataOut_payload_0_14433 : _zz_dataOut_payload_0_14436);
    _zz_dataOut_payload_0_14441 <= (_zz_dataOut_payload_0_14438 ? _zz_dataOut_payload_0_14436 : _zz_dataOut_payload_0_14433);
    _zz_dataOut_payload_0_14442 <= (_zz_dataOut_payload_0_14439 ? _zz_dataOut_payload_0_14434 : _zz_dataOut_payload_0_14437);
    _zz_dataOut_payload_0_14443 <= (_zz_dataOut_payload_0_14439 ? _zz_dataOut_payload_0_14437 : _zz_dataOut_payload_0_14434);
    _zz_dataOut_payload_0_14452 <= (_zz_dataOut_payload_0_14450 ? _zz_dataOut_payload_0_14445 : _zz_dataOut_payload_0_14448);
    _zz_dataOut_payload_0_14453 <= (_zz_dataOut_payload_0_14450 ? _zz_dataOut_payload_0_14448 : _zz_dataOut_payload_0_14445);
    _zz_dataOut_payload_0_14454 <= (_zz_dataOut_payload_0_14451 ? _zz_dataOut_payload_0_14446 : _zz_dataOut_payload_0_14449);
    _zz_dataOut_payload_0_14455 <= (_zz_dataOut_payload_0_14451 ? _zz_dataOut_payload_0_14449 : _zz_dataOut_payload_0_14446);
    _zz_dataOut_payload_0_14456 <= _zz_dataOut_payload_0_14440;
    _zz_dataOut_payload_0_14457 <= _zz_dataOut_payload_0_14441;
    _zz_dataOut_payload_0_14458 <= _zz_dataOut_payload_0_14442;
    _zz_dataOut_payload_0_14459 <= _zz_dataOut_payload_0_14443;
    _zz_dataOut_payload_0_14460 <= _zz_dataOut_payload_0_14452;
    _zz_dataOut_payload_0_14461 <= _zz_dataOut_payload_0_14453;
    _zz_dataOut_payload_0_14462 <= _zz_dataOut_payload_0_14454;
    _zz_dataOut_payload_0_14463 <= _zz_dataOut_payload_0_14455;
    _zz_dataOut_payload_0_14464 <= _zz_dataOut_payload_0_14412;
    _zz_dataOut_payload_0_14465 <= _zz_dataOut_payload_0_14413;
    _zz_dataOut_payload_0_14466 <= _zz_dataOut_payload_0_14414;
    _zz_dataOut_payload_0_14467 <= _zz_dataOut_payload_0_14415;
    _zz_dataOut_payload_0_14468 <= _zz_dataOut_payload_0_14416;
    _zz_dataOut_payload_0_14469 <= _zz_dataOut_payload_0_14417;
    _zz_dataOut_payload_0_14470 <= _zz_dataOut_payload_0_14418;
    _zz_dataOut_payload_0_14471 <= _zz_dataOut_payload_0_14419;
    _zz_dataOut_payload_0_14472 <= _zz_dataOut_payload_0_14456;
    _zz_dataOut_payload_0_14473 <= _zz_dataOut_payload_0_14457;
    _zz_dataOut_payload_0_14474 <= _zz_dataOut_payload_0_14458;
    _zz_dataOut_payload_0_14475 <= _zz_dataOut_payload_0_14459;
    _zz_dataOut_payload_0_14476 <= _zz_dataOut_payload_0_14460;
    _zz_dataOut_payload_0_14477 <= _zz_dataOut_payload_0_14461;
    _zz_dataOut_payload_0_14478 <= _zz_dataOut_payload_0_14462;
    _zz_dataOut_payload_0_14479 <= _zz_dataOut_payload_0_14463;
    _zz_dataOut_payload_0_14480 <= _zz_dataOut_payload_0_14336;
    _zz_dataOut_payload_0_14481 <= _zz_dataOut_payload_0_14337;
    _zz_dataOut_payload_0_14482 <= _zz_dataOut_payload_0_14338;
    _zz_dataOut_payload_0_14483 <= _zz_dataOut_payload_0_14339;
    _zz_dataOut_payload_0_14484 <= _zz_dataOut_payload_0_14340;
    _zz_dataOut_payload_0_14485 <= _zz_dataOut_payload_0_14341;
    _zz_dataOut_payload_0_14486 <= _zz_dataOut_payload_0_14342;
    _zz_dataOut_payload_0_14487 <= _zz_dataOut_payload_0_14343;
    _zz_dataOut_payload_0_14488 <= _zz_dataOut_payload_0_14344;
    _zz_dataOut_payload_0_14489 <= _zz_dataOut_payload_0_14345;
    _zz_dataOut_payload_0_14490 <= _zz_dataOut_payload_0_14346;
    _zz_dataOut_payload_0_14491 <= _zz_dataOut_payload_0_14347;
    _zz_dataOut_payload_0_14492 <= _zz_dataOut_payload_0_14348;
    _zz_dataOut_payload_0_14493 <= _zz_dataOut_payload_0_14349;
    _zz_dataOut_payload_0_14494 <= _zz_dataOut_payload_0_14350;
    _zz_dataOut_payload_0_14495 <= _zz_dataOut_payload_0_14351;
    _zz_dataOut_payload_0_14496 <= _zz_dataOut_payload_0_14464;
    _zz_dataOut_payload_0_14497 <= _zz_dataOut_payload_0_14465;
    _zz_dataOut_payload_0_14498 <= _zz_dataOut_payload_0_14466;
    _zz_dataOut_payload_0_14499 <= _zz_dataOut_payload_0_14467;
    _zz_dataOut_payload_0_14500 <= _zz_dataOut_payload_0_14468;
    _zz_dataOut_payload_0_14501 <= _zz_dataOut_payload_0_14469;
    _zz_dataOut_payload_0_14502 <= _zz_dataOut_payload_0_14470;
    _zz_dataOut_payload_0_14503 <= _zz_dataOut_payload_0_14471;
    _zz_dataOut_payload_0_14504 <= _zz_dataOut_payload_0_14472;
    _zz_dataOut_payload_0_14505 <= _zz_dataOut_payload_0_14473;
    _zz_dataOut_payload_0_14506 <= _zz_dataOut_payload_0_14474;
    _zz_dataOut_payload_0_14507 <= _zz_dataOut_payload_0_14475;
    _zz_dataOut_payload_0_14508 <= _zz_dataOut_payload_0_14476;
    _zz_dataOut_payload_0_14509 <= _zz_dataOut_payload_0_14477;
    _zz_dataOut_payload_0_14510 <= _zz_dataOut_payload_0_14478;
    _zz_dataOut_payload_0_14511 <= _zz_dataOut_payload_0_14479;
    _zz_dataOut_payload_0_14604 <= (_zz_dataOut_payload_0_14602 ? _zz_dataOut_payload_0_14597 : _zz_dataOut_payload_0_14600);
    _zz_dataOut_payload_0_14605 <= (_zz_dataOut_payload_0_14602 ? _zz_dataOut_payload_0_14600 : _zz_dataOut_payload_0_14597);
    _zz_dataOut_payload_0_14606 <= (_zz_dataOut_payload_0_14603 ? _zz_dataOut_payload_0_14598 : _zz_dataOut_payload_0_14601);
    _zz_dataOut_payload_0_14607 <= (_zz_dataOut_payload_0_14603 ? _zz_dataOut_payload_0_14601 : _zz_dataOut_payload_0_14598);
    _zz_dataOut_payload_0_14616 <= (_zz_dataOut_payload_0_14614 ? _zz_dataOut_payload_0_14609 : _zz_dataOut_payload_0_14612);
    _zz_dataOut_payload_0_14617 <= (_zz_dataOut_payload_0_14614 ? _zz_dataOut_payload_0_14612 : _zz_dataOut_payload_0_14609);
    _zz_dataOut_payload_0_14618 <= (_zz_dataOut_payload_0_14615 ? _zz_dataOut_payload_0_14610 : _zz_dataOut_payload_0_14613);
    _zz_dataOut_payload_0_14619 <= (_zz_dataOut_payload_0_14615 ? _zz_dataOut_payload_0_14613 : _zz_dataOut_payload_0_14610);
    _zz_dataOut_payload_0_14620 <= _zz_dataOut_payload_0_14604;
    _zz_dataOut_payload_0_14621 <= _zz_dataOut_payload_0_14605;
    _zz_dataOut_payload_0_14622 <= _zz_dataOut_payload_0_14606;
    _zz_dataOut_payload_0_14623 <= _zz_dataOut_payload_0_14607;
    _zz_dataOut_payload_0_14624 <= _zz_dataOut_payload_0_14616;
    _zz_dataOut_payload_0_14625 <= _zz_dataOut_payload_0_14617;
    _zz_dataOut_payload_0_14626 <= _zz_dataOut_payload_0_14618;
    _zz_dataOut_payload_0_14627 <= _zz_dataOut_payload_0_14619;
    _zz_dataOut_payload_0_14648 <= (_zz_dataOut_payload_0_14646 ? _zz_dataOut_payload_0_14641 : _zz_dataOut_payload_0_14644);
    _zz_dataOut_payload_0_14649 <= (_zz_dataOut_payload_0_14646 ? _zz_dataOut_payload_0_14644 : _zz_dataOut_payload_0_14641);
    _zz_dataOut_payload_0_14650 <= (_zz_dataOut_payload_0_14647 ? _zz_dataOut_payload_0_14642 : _zz_dataOut_payload_0_14645);
    _zz_dataOut_payload_0_14651 <= (_zz_dataOut_payload_0_14647 ? _zz_dataOut_payload_0_14645 : _zz_dataOut_payload_0_14642);
    _zz_dataOut_payload_0_14660 <= (_zz_dataOut_payload_0_14658 ? _zz_dataOut_payload_0_14653 : _zz_dataOut_payload_0_14656);
    _zz_dataOut_payload_0_14661 <= (_zz_dataOut_payload_0_14658 ? _zz_dataOut_payload_0_14656 : _zz_dataOut_payload_0_14653);
    _zz_dataOut_payload_0_14662 <= (_zz_dataOut_payload_0_14659 ? _zz_dataOut_payload_0_14654 : _zz_dataOut_payload_0_14657);
    _zz_dataOut_payload_0_14663 <= (_zz_dataOut_payload_0_14659 ? _zz_dataOut_payload_0_14657 : _zz_dataOut_payload_0_14654);
    _zz_dataOut_payload_0_14664 <= _zz_dataOut_payload_0_14648;
    _zz_dataOut_payload_0_14665 <= _zz_dataOut_payload_0_14649;
    _zz_dataOut_payload_0_14666 <= _zz_dataOut_payload_0_14650;
    _zz_dataOut_payload_0_14667 <= _zz_dataOut_payload_0_14651;
    _zz_dataOut_payload_0_14668 <= _zz_dataOut_payload_0_14660;
    _zz_dataOut_payload_0_14669 <= _zz_dataOut_payload_0_14661;
    _zz_dataOut_payload_0_14670 <= _zz_dataOut_payload_0_14662;
    _zz_dataOut_payload_0_14671 <= _zz_dataOut_payload_0_14663;
    _zz_dataOut_payload_0_14672 <= _zz_dataOut_payload_0_14620;
    _zz_dataOut_payload_0_14673 <= _zz_dataOut_payload_0_14621;
    _zz_dataOut_payload_0_14674 <= _zz_dataOut_payload_0_14622;
    _zz_dataOut_payload_0_14675 <= _zz_dataOut_payload_0_14623;
    _zz_dataOut_payload_0_14676 <= _zz_dataOut_payload_0_14624;
    _zz_dataOut_payload_0_14677 <= _zz_dataOut_payload_0_14625;
    _zz_dataOut_payload_0_14678 <= _zz_dataOut_payload_0_14626;
    _zz_dataOut_payload_0_14679 <= _zz_dataOut_payload_0_14627;
    _zz_dataOut_payload_0_14680 <= _zz_dataOut_payload_0_14664;
    _zz_dataOut_payload_0_14681 <= _zz_dataOut_payload_0_14665;
    _zz_dataOut_payload_0_14682 <= _zz_dataOut_payload_0_14666;
    _zz_dataOut_payload_0_14683 <= _zz_dataOut_payload_0_14667;
    _zz_dataOut_payload_0_14684 <= _zz_dataOut_payload_0_14668;
    _zz_dataOut_payload_0_14685 <= _zz_dataOut_payload_0_14669;
    _zz_dataOut_payload_0_14686 <= _zz_dataOut_payload_0_14670;
    _zz_dataOut_payload_0_14687 <= _zz_dataOut_payload_0_14671;
    _zz_dataOut_payload_0_14732 <= (_zz_dataOut_payload_0_14730 ? _zz_dataOut_payload_0_14725 : _zz_dataOut_payload_0_14728);
    _zz_dataOut_payload_0_14733 <= (_zz_dataOut_payload_0_14730 ? _zz_dataOut_payload_0_14728 : _zz_dataOut_payload_0_14725);
    _zz_dataOut_payload_0_14734 <= (_zz_dataOut_payload_0_14731 ? _zz_dataOut_payload_0_14726 : _zz_dataOut_payload_0_14729);
    _zz_dataOut_payload_0_14735 <= (_zz_dataOut_payload_0_14731 ? _zz_dataOut_payload_0_14729 : _zz_dataOut_payload_0_14726);
    _zz_dataOut_payload_0_14744 <= (_zz_dataOut_payload_0_14742 ? _zz_dataOut_payload_0_14737 : _zz_dataOut_payload_0_14740);
    _zz_dataOut_payload_0_14745 <= (_zz_dataOut_payload_0_14742 ? _zz_dataOut_payload_0_14740 : _zz_dataOut_payload_0_14737);
    _zz_dataOut_payload_0_14746 <= (_zz_dataOut_payload_0_14743 ? _zz_dataOut_payload_0_14738 : _zz_dataOut_payload_0_14741);
    _zz_dataOut_payload_0_14747 <= (_zz_dataOut_payload_0_14743 ? _zz_dataOut_payload_0_14741 : _zz_dataOut_payload_0_14738);
    _zz_dataOut_payload_0_14748 <= _zz_dataOut_payload_0_14732;
    _zz_dataOut_payload_0_14749 <= _zz_dataOut_payload_0_14733;
    _zz_dataOut_payload_0_14750 <= _zz_dataOut_payload_0_14734;
    _zz_dataOut_payload_0_14751 <= _zz_dataOut_payload_0_14735;
    _zz_dataOut_payload_0_14752 <= _zz_dataOut_payload_0_14744;
    _zz_dataOut_payload_0_14753 <= _zz_dataOut_payload_0_14745;
    _zz_dataOut_payload_0_14754 <= _zz_dataOut_payload_0_14746;
    _zz_dataOut_payload_0_14755 <= _zz_dataOut_payload_0_14747;
    _zz_dataOut_payload_0_14776 <= (_zz_dataOut_payload_0_14774 ? _zz_dataOut_payload_0_14769 : _zz_dataOut_payload_0_14772);
    _zz_dataOut_payload_0_14777 <= (_zz_dataOut_payload_0_14774 ? _zz_dataOut_payload_0_14772 : _zz_dataOut_payload_0_14769);
    _zz_dataOut_payload_0_14778 <= (_zz_dataOut_payload_0_14775 ? _zz_dataOut_payload_0_14770 : _zz_dataOut_payload_0_14773);
    _zz_dataOut_payload_0_14779 <= (_zz_dataOut_payload_0_14775 ? _zz_dataOut_payload_0_14773 : _zz_dataOut_payload_0_14770);
    _zz_dataOut_payload_0_14788 <= (_zz_dataOut_payload_0_14786 ? _zz_dataOut_payload_0_14781 : _zz_dataOut_payload_0_14784);
    _zz_dataOut_payload_0_14789 <= (_zz_dataOut_payload_0_14786 ? _zz_dataOut_payload_0_14784 : _zz_dataOut_payload_0_14781);
    _zz_dataOut_payload_0_14790 <= (_zz_dataOut_payload_0_14787 ? _zz_dataOut_payload_0_14782 : _zz_dataOut_payload_0_14785);
    _zz_dataOut_payload_0_14791 <= (_zz_dataOut_payload_0_14787 ? _zz_dataOut_payload_0_14785 : _zz_dataOut_payload_0_14782);
    _zz_dataOut_payload_0_14792 <= _zz_dataOut_payload_0_14776;
    _zz_dataOut_payload_0_14793 <= _zz_dataOut_payload_0_14777;
    _zz_dataOut_payload_0_14794 <= _zz_dataOut_payload_0_14778;
    _zz_dataOut_payload_0_14795 <= _zz_dataOut_payload_0_14779;
    _zz_dataOut_payload_0_14796 <= _zz_dataOut_payload_0_14788;
    _zz_dataOut_payload_0_14797 <= _zz_dataOut_payload_0_14789;
    _zz_dataOut_payload_0_14798 <= _zz_dataOut_payload_0_14790;
    _zz_dataOut_payload_0_14799 <= _zz_dataOut_payload_0_14791;
    _zz_dataOut_payload_0_14800 <= _zz_dataOut_payload_0_14748;
    _zz_dataOut_payload_0_14801 <= _zz_dataOut_payload_0_14749;
    _zz_dataOut_payload_0_14802 <= _zz_dataOut_payload_0_14750;
    _zz_dataOut_payload_0_14803 <= _zz_dataOut_payload_0_14751;
    _zz_dataOut_payload_0_14804 <= _zz_dataOut_payload_0_14752;
    _zz_dataOut_payload_0_14805 <= _zz_dataOut_payload_0_14753;
    _zz_dataOut_payload_0_14806 <= _zz_dataOut_payload_0_14754;
    _zz_dataOut_payload_0_14807 <= _zz_dataOut_payload_0_14755;
    _zz_dataOut_payload_0_14808 <= _zz_dataOut_payload_0_14792;
    _zz_dataOut_payload_0_14809 <= _zz_dataOut_payload_0_14793;
    _zz_dataOut_payload_0_14810 <= _zz_dataOut_payload_0_14794;
    _zz_dataOut_payload_0_14811 <= _zz_dataOut_payload_0_14795;
    _zz_dataOut_payload_0_14812 <= _zz_dataOut_payload_0_14796;
    _zz_dataOut_payload_0_14813 <= _zz_dataOut_payload_0_14797;
    _zz_dataOut_payload_0_14814 <= _zz_dataOut_payload_0_14798;
    _zz_dataOut_payload_0_14815 <= _zz_dataOut_payload_0_14799;
    _zz_dataOut_payload_0_14816 <= _zz_dataOut_payload_0_14672;
    _zz_dataOut_payload_0_14817 <= _zz_dataOut_payload_0_14673;
    _zz_dataOut_payload_0_14818 <= _zz_dataOut_payload_0_14674;
    _zz_dataOut_payload_0_14819 <= _zz_dataOut_payload_0_14675;
    _zz_dataOut_payload_0_14820 <= _zz_dataOut_payload_0_14676;
    _zz_dataOut_payload_0_14821 <= _zz_dataOut_payload_0_14677;
    _zz_dataOut_payload_0_14822 <= _zz_dataOut_payload_0_14678;
    _zz_dataOut_payload_0_14823 <= _zz_dataOut_payload_0_14679;
    _zz_dataOut_payload_0_14824 <= _zz_dataOut_payload_0_14680;
    _zz_dataOut_payload_0_14825 <= _zz_dataOut_payload_0_14681;
    _zz_dataOut_payload_0_14826 <= _zz_dataOut_payload_0_14682;
    _zz_dataOut_payload_0_14827 <= _zz_dataOut_payload_0_14683;
    _zz_dataOut_payload_0_14828 <= _zz_dataOut_payload_0_14684;
    _zz_dataOut_payload_0_14829 <= _zz_dataOut_payload_0_14685;
    _zz_dataOut_payload_0_14830 <= _zz_dataOut_payload_0_14686;
    _zz_dataOut_payload_0_14831 <= _zz_dataOut_payload_0_14687;
    _zz_dataOut_payload_0_14832 <= _zz_dataOut_payload_0_14800;
    _zz_dataOut_payload_0_14833 <= _zz_dataOut_payload_0_14801;
    _zz_dataOut_payload_0_14834 <= _zz_dataOut_payload_0_14802;
    _zz_dataOut_payload_0_14835 <= _zz_dataOut_payload_0_14803;
    _zz_dataOut_payload_0_14836 <= _zz_dataOut_payload_0_14804;
    _zz_dataOut_payload_0_14837 <= _zz_dataOut_payload_0_14805;
    _zz_dataOut_payload_0_14838 <= _zz_dataOut_payload_0_14806;
    _zz_dataOut_payload_0_14839 <= _zz_dataOut_payload_0_14807;
    _zz_dataOut_payload_0_14840 <= _zz_dataOut_payload_0_14808;
    _zz_dataOut_payload_0_14841 <= _zz_dataOut_payload_0_14809;
    _zz_dataOut_payload_0_14842 <= _zz_dataOut_payload_0_14810;
    _zz_dataOut_payload_0_14843 <= _zz_dataOut_payload_0_14811;
    _zz_dataOut_payload_0_14844 <= _zz_dataOut_payload_0_14812;
    _zz_dataOut_payload_0_14845 <= _zz_dataOut_payload_0_14813;
    _zz_dataOut_payload_0_14846 <= _zz_dataOut_payload_0_14814;
    _zz_dataOut_payload_0_14847 <= _zz_dataOut_payload_0_14815;
    _zz_dataOut_payload_0_14848 <= _zz_dataOut_payload_0_14480;
    _zz_dataOut_payload_0_14849 <= _zz_dataOut_payload_0_14481;
    _zz_dataOut_payload_0_14850 <= _zz_dataOut_payload_0_14482;
    _zz_dataOut_payload_0_14851 <= _zz_dataOut_payload_0_14483;
    _zz_dataOut_payload_0_14852 <= _zz_dataOut_payload_0_14484;
    _zz_dataOut_payload_0_14853 <= _zz_dataOut_payload_0_14485;
    _zz_dataOut_payload_0_14854 <= _zz_dataOut_payload_0_14486;
    _zz_dataOut_payload_0_14855 <= _zz_dataOut_payload_0_14487;
    _zz_dataOut_payload_0_14856 <= _zz_dataOut_payload_0_14488;
    _zz_dataOut_payload_0_14857 <= _zz_dataOut_payload_0_14489;
    _zz_dataOut_payload_0_14858 <= _zz_dataOut_payload_0_14490;
    _zz_dataOut_payload_0_14859 <= _zz_dataOut_payload_0_14491;
    _zz_dataOut_payload_0_14860 <= _zz_dataOut_payload_0_14492;
    _zz_dataOut_payload_0_14861 <= _zz_dataOut_payload_0_14493;
    _zz_dataOut_payload_0_14862 <= _zz_dataOut_payload_0_14494;
    _zz_dataOut_payload_0_14863 <= _zz_dataOut_payload_0_14495;
    _zz_dataOut_payload_0_14864 <= _zz_dataOut_payload_0_14496;
    _zz_dataOut_payload_0_14865 <= _zz_dataOut_payload_0_14497;
    _zz_dataOut_payload_0_14866 <= _zz_dataOut_payload_0_14498;
    _zz_dataOut_payload_0_14867 <= _zz_dataOut_payload_0_14499;
    _zz_dataOut_payload_0_14868 <= _zz_dataOut_payload_0_14500;
    _zz_dataOut_payload_0_14869 <= _zz_dataOut_payload_0_14501;
    _zz_dataOut_payload_0_14870 <= _zz_dataOut_payload_0_14502;
    _zz_dataOut_payload_0_14871 <= _zz_dataOut_payload_0_14503;
    _zz_dataOut_payload_0_14872 <= _zz_dataOut_payload_0_14504;
    _zz_dataOut_payload_0_14873 <= _zz_dataOut_payload_0_14505;
    _zz_dataOut_payload_0_14874 <= _zz_dataOut_payload_0_14506;
    _zz_dataOut_payload_0_14875 <= _zz_dataOut_payload_0_14507;
    _zz_dataOut_payload_0_14876 <= _zz_dataOut_payload_0_14508;
    _zz_dataOut_payload_0_14877 <= _zz_dataOut_payload_0_14509;
    _zz_dataOut_payload_0_14878 <= _zz_dataOut_payload_0_14510;
    _zz_dataOut_payload_0_14879 <= _zz_dataOut_payload_0_14511;
    _zz_dataOut_payload_0_14880 <= _zz_dataOut_payload_0_14816;
    _zz_dataOut_payload_0_14881 <= _zz_dataOut_payload_0_14817;
    _zz_dataOut_payload_0_14882 <= _zz_dataOut_payload_0_14818;
    _zz_dataOut_payload_0_14883 <= _zz_dataOut_payload_0_14819;
    _zz_dataOut_payload_0_14884 <= _zz_dataOut_payload_0_14820;
    _zz_dataOut_payload_0_14885 <= _zz_dataOut_payload_0_14821;
    _zz_dataOut_payload_0_14886 <= _zz_dataOut_payload_0_14822;
    _zz_dataOut_payload_0_14887 <= _zz_dataOut_payload_0_14823;
    _zz_dataOut_payload_0_14888 <= _zz_dataOut_payload_0_14824;
    _zz_dataOut_payload_0_14889 <= _zz_dataOut_payload_0_14825;
    _zz_dataOut_payload_0_14890 <= _zz_dataOut_payload_0_14826;
    _zz_dataOut_payload_0_14891 <= _zz_dataOut_payload_0_14827;
    _zz_dataOut_payload_0_14892 <= _zz_dataOut_payload_0_14828;
    _zz_dataOut_payload_0_14893 <= _zz_dataOut_payload_0_14829;
    _zz_dataOut_payload_0_14894 <= _zz_dataOut_payload_0_14830;
    _zz_dataOut_payload_0_14895 <= _zz_dataOut_payload_0_14831;
    _zz_dataOut_payload_0_14896 <= _zz_dataOut_payload_0_14832;
    _zz_dataOut_payload_0_14897 <= _zz_dataOut_payload_0_14833;
    _zz_dataOut_payload_0_14898 <= _zz_dataOut_payload_0_14834;
    _zz_dataOut_payload_0_14899 <= _zz_dataOut_payload_0_14835;
    _zz_dataOut_payload_0_14900 <= _zz_dataOut_payload_0_14836;
    _zz_dataOut_payload_0_14901 <= _zz_dataOut_payload_0_14837;
    _zz_dataOut_payload_0_14902 <= _zz_dataOut_payload_0_14838;
    _zz_dataOut_payload_0_14903 <= _zz_dataOut_payload_0_14839;
    _zz_dataOut_payload_0_14904 <= _zz_dataOut_payload_0_14840;
    _zz_dataOut_payload_0_14905 <= _zz_dataOut_payload_0_14841;
    _zz_dataOut_payload_0_14906 <= _zz_dataOut_payload_0_14842;
    _zz_dataOut_payload_0_14907 <= _zz_dataOut_payload_0_14843;
    _zz_dataOut_payload_0_14908 <= _zz_dataOut_payload_0_14844;
    _zz_dataOut_payload_0_14909 <= _zz_dataOut_payload_0_14845;
    _zz_dataOut_payload_0_14910 <= _zz_dataOut_payload_0_14846;
    _zz_dataOut_payload_0_14911 <= _zz_dataOut_payload_0_14847;
    _zz_dataOut_payload_0_15100 <= (_zz_dataOut_payload_0_15098 ? _zz_dataOut_payload_0_15093 : _zz_dataOut_payload_0_15096);
    _zz_dataOut_payload_0_15101 <= (_zz_dataOut_payload_0_15098 ? _zz_dataOut_payload_0_15096 : _zz_dataOut_payload_0_15093);
    _zz_dataOut_payload_0_15102 <= (_zz_dataOut_payload_0_15099 ? _zz_dataOut_payload_0_15094 : _zz_dataOut_payload_0_15097);
    _zz_dataOut_payload_0_15103 <= (_zz_dataOut_payload_0_15099 ? _zz_dataOut_payload_0_15097 : _zz_dataOut_payload_0_15094);
    _zz_dataOut_payload_0_15112 <= (_zz_dataOut_payload_0_15110 ? _zz_dataOut_payload_0_15105 : _zz_dataOut_payload_0_15108);
    _zz_dataOut_payload_0_15113 <= (_zz_dataOut_payload_0_15110 ? _zz_dataOut_payload_0_15108 : _zz_dataOut_payload_0_15105);
    _zz_dataOut_payload_0_15114 <= (_zz_dataOut_payload_0_15111 ? _zz_dataOut_payload_0_15106 : _zz_dataOut_payload_0_15109);
    _zz_dataOut_payload_0_15115 <= (_zz_dataOut_payload_0_15111 ? _zz_dataOut_payload_0_15109 : _zz_dataOut_payload_0_15106);
    _zz_dataOut_payload_0_15116 <= _zz_dataOut_payload_0_15100;
    _zz_dataOut_payload_0_15117 <= _zz_dataOut_payload_0_15101;
    _zz_dataOut_payload_0_15118 <= _zz_dataOut_payload_0_15102;
    _zz_dataOut_payload_0_15119 <= _zz_dataOut_payload_0_15103;
    _zz_dataOut_payload_0_15120 <= _zz_dataOut_payload_0_15112;
    _zz_dataOut_payload_0_15121 <= _zz_dataOut_payload_0_15113;
    _zz_dataOut_payload_0_15122 <= _zz_dataOut_payload_0_15114;
    _zz_dataOut_payload_0_15123 <= _zz_dataOut_payload_0_15115;
    _zz_dataOut_payload_0_15144 <= (_zz_dataOut_payload_0_15142 ? _zz_dataOut_payload_0_15137 : _zz_dataOut_payload_0_15140);
    _zz_dataOut_payload_0_15145 <= (_zz_dataOut_payload_0_15142 ? _zz_dataOut_payload_0_15140 : _zz_dataOut_payload_0_15137);
    _zz_dataOut_payload_0_15146 <= (_zz_dataOut_payload_0_15143 ? _zz_dataOut_payload_0_15138 : _zz_dataOut_payload_0_15141);
    _zz_dataOut_payload_0_15147 <= (_zz_dataOut_payload_0_15143 ? _zz_dataOut_payload_0_15141 : _zz_dataOut_payload_0_15138);
    _zz_dataOut_payload_0_15156 <= (_zz_dataOut_payload_0_15154 ? _zz_dataOut_payload_0_15149 : _zz_dataOut_payload_0_15152);
    _zz_dataOut_payload_0_15157 <= (_zz_dataOut_payload_0_15154 ? _zz_dataOut_payload_0_15152 : _zz_dataOut_payload_0_15149);
    _zz_dataOut_payload_0_15158 <= (_zz_dataOut_payload_0_15155 ? _zz_dataOut_payload_0_15150 : _zz_dataOut_payload_0_15153);
    _zz_dataOut_payload_0_15159 <= (_zz_dataOut_payload_0_15155 ? _zz_dataOut_payload_0_15153 : _zz_dataOut_payload_0_15150);
    _zz_dataOut_payload_0_15160 <= _zz_dataOut_payload_0_15144;
    _zz_dataOut_payload_0_15161 <= _zz_dataOut_payload_0_15145;
    _zz_dataOut_payload_0_15162 <= _zz_dataOut_payload_0_15146;
    _zz_dataOut_payload_0_15163 <= _zz_dataOut_payload_0_15147;
    _zz_dataOut_payload_0_15164 <= _zz_dataOut_payload_0_15156;
    _zz_dataOut_payload_0_15165 <= _zz_dataOut_payload_0_15157;
    _zz_dataOut_payload_0_15166 <= _zz_dataOut_payload_0_15158;
    _zz_dataOut_payload_0_15167 <= _zz_dataOut_payload_0_15159;
    _zz_dataOut_payload_0_15168 <= _zz_dataOut_payload_0_15116;
    _zz_dataOut_payload_0_15169 <= _zz_dataOut_payload_0_15117;
    _zz_dataOut_payload_0_15170 <= _zz_dataOut_payload_0_15118;
    _zz_dataOut_payload_0_15171 <= _zz_dataOut_payload_0_15119;
    _zz_dataOut_payload_0_15172 <= _zz_dataOut_payload_0_15120;
    _zz_dataOut_payload_0_15173 <= _zz_dataOut_payload_0_15121;
    _zz_dataOut_payload_0_15174 <= _zz_dataOut_payload_0_15122;
    _zz_dataOut_payload_0_15175 <= _zz_dataOut_payload_0_15123;
    _zz_dataOut_payload_0_15176 <= _zz_dataOut_payload_0_15160;
    _zz_dataOut_payload_0_15177 <= _zz_dataOut_payload_0_15161;
    _zz_dataOut_payload_0_15178 <= _zz_dataOut_payload_0_15162;
    _zz_dataOut_payload_0_15179 <= _zz_dataOut_payload_0_15163;
    _zz_dataOut_payload_0_15180 <= _zz_dataOut_payload_0_15164;
    _zz_dataOut_payload_0_15181 <= _zz_dataOut_payload_0_15165;
    _zz_dataOut_payload_0_15182 <= _zz_dataOut_payload_0_15166;
    _zz_dataOut_payload_0_15183 <= _zz_dataOut_payload_0_15167;
    _zz_dataOut_payload_0_15228 <= (_zz_dataOut_payload_0_15226 ? _zz_dataOut_payload_0_15221 : _zz_dataOut_payload_0_15224);
    _zz_dataOut_payload_0_15229 <= (_zz_dataOut_payload_0_15226 ? _zz_dataOut_payload_0_15224 : _zz_dataOut_payload_0_15221);
    _zz_dataOut_payload_0_15230 <= (_zz_dataOut_payload_0_15227 ? _zz_dataOut_payload_0_15222 : _zz_dataOut_payload_0_15225);
    _zz_dataOut_payload_0_15231 <= (_zz_dataOut_payload_0_15227 ? _zz_dataOut_payload_0_15225 : _zz_dataOut_payload_0_15222);
    _zz_dataOut_payload_0_15240 <= (_zz_dataOut_payload_0_15238 ? _zz_dataOut_payload_0_15233 : _zz_dataOut_payload_0_15236);
    _zz_dataOut_payload_0_15241 <= (_zz_dataOut_payload_0_15238 ? _zz_dataOut_payload_0_15236 : _zz_dataOut_payload_0_15233);
    _zz_dataOut_payload_0_15242 <= (_zz_dataOut_payload_0_15239 ? _zz_dataOut_payload_0_15234 : _zz_dataOut_payload_0_15237);
    _zz_dataOut_payload_0_15243 <= (_zz_dataOut_payload_0_15239 ? _zz_dataOut_payload_0_15237 : _zz_dataOut_payload_0_15234);
    _zz_dataOut_payload_0_15244 <= _zz_dataOut_payload_0_15228;
    _zz_dataOut_payload_0_15245 <= _zz_dataOut_payload_0_15229;
    _zz_dataOut_payload_0_15246 <= _zz_dataOut_payload_0_15230;
    _zz_dataOut_payload_0_15247 <= _zz_dataOut_payload_0_15231;
    _zz_dataOut_payload_0_15248 <= _zz_dataOut_payload_0_15240;
    _zz_dataOut_payload_0_15249 <= _zz_dataOut_payload_0_15241;
    _zz_dataOut_payload_0_15250 <= _zz_dataOut_payload_0_15242;
    _zz_dataOut_payload_0_15251 <= _zz_dataOut_payload_0_15243;
    _zz_dataOut_payload_0_15272 <= (_zz_dataOut_payload_0_15270 ? _zz_dataOut_payload_0_15265 : _zz_dataOut_payload_0_15268);
    _zz_dataOut_payload_0_15273 <= (_zz_dataOut_payload_0_15270 ? _zz_dataOut_payload_0_15268 : _zz_dataOut_payload_0_15265);
    _zz_dataOut_payload_0_15274 <= (_zz_dataOut_payload_0_15271 ? _zz_dataOut_payload_0_15266 : _zz_dataOut_payload_0_15269);
    _zz_dataOut_payload_0_15275 <= (_zz_dataOut_payload_0_15271 ? _zz_dataOut_payload_0_15269 : _zz_dataOut_payload_0_15266);
    _zz_dataOut_payload_0_15284 <= (_zz_dataOut_payload_0_15282 ? _zz_dataOut_payload_0_15277 : _zz_dataOut_payload_0_15280);
    _zz_dataOut_payload_0_15285 <= (_zz_dataOut_payload_0_15282 ? _zz_dataOut_payload_0_15280 : _zz_dataOut_payload_0_15277);
    _zz_dataOut_payload_0_15286 <= (_zz_dataOut_payload_0_15283 ? _zz_dataOut_payload_0_15278 : _zz_dataOut_payload_0_15281);
    _zz_dataOut_payload_0_15287 <= (_zz_dataOut_payload_0_15283 ? _zz_dataOut_payload_0_15281 : _zz_dataOut_payload_0_15278);
    _zz_dataOut_payload_0_15288 <= _zz_dataOut_payload_0_15272;
    _zz_dataOut_payload_0_15289 <= _zz_dataOut_payload_0_15273;
    _zz_dataOut_payload_0_15290 <= _zz_dataOut_payload_0_15274;
    _zz_dataOut_payload_0_15291 <= _zz_dataOut_payload_0_15275;
    _zz_dataOut_payload_0_15292 <= _zz_dataOut_payload_0_15284;
    _zz_dataOut_payload_0_15293 <= _zz_dataOut_payload_0_15285;
    _zz_dataOut_payload_0_15294 <= _zz_dataOut_payload_0_15286;
    _zz_dataOut_payload_0_15295 <= _zz_dataOut_payload_0_15287;
    _zz_dataOut_payload_0_15296 <= _zz_dataOut_payload_0_15244;
    _zz_dataOut_payload_0_15297 <= _zz_dataOut_payload_0_15245;
    _zz_dataOut_payload_0_15298 <= _zz_dataOut_payload_0_15246;
    _zz_dataOut_payload_0_15299 <= _zz_dataOut_payload_0_15247;
    _zz_dataOut_payload_0_15300 <= _zz_dataOut_payload_0_15248;
    _zz_dataOut_payload_0_15301 <= _zz_dataOut_payload_0_15249;
    _zz_dataOut_payload_0_15302 <= _zz_dataOut_payload_0_15250;
    _zz_dataOut_payload_0_15303 <= _zz_dataOut_payload_0_15251;
    _zz_dataOut_payload_0_15304 <= _zz_dataOut_payload_0_15288;
    _zz_dataOut_payload_0_15305 <= _zz_dataOut_payload_0_15289;
    _zz_dataOut_payload_0_15306 <= _zz_dataOut_payload_0_15290;
    _zz_dataOut_payload_0_15307 <= _zz_dataOut_payload_0_15291;
    _zz_dataOut_payload_0_15308 <= _zz_dataOut_payload_0_15292;
    _zz_dataOut_payload_0_15309 <= _zz_dataOut_payload_0_15293;
    _zz_dataOut_payload_0_15310 <= _zz_dataOut_payload_0_15294;
    _zz_dataOut_payload_0_15311 <= _zz_dataOut_payload_0_15295;
    _zz_dataOut_payload_0_15312 <= _zz_dataOut_payload_0_15168;
    _zz_dataOut_payload_0_15313 <= _zz_dataOut_payload_0_15169;
    _zz_dataOut_payload_0_15314 <= _zz_dataOut_payload_0_15170;
    _zz_dataOut_payload_0_15315 <= _zz_dataOut_payload_0_15171;
    _zz_dataOut_payload_0_15316 <= _zz_dataOut_payload_0_15172;
    _zz_dataOut_payload_0_15317 <= _zz_dataOut_payload_0_15173;
    _zz_dataOut_payload_0_15318 <= _zz_dataOut_payload_0_15174;
    _zz_dataOut_payload_0_15319 <= _zz_dataOut_payload_0_15175;
    _zz_dataOut_payload_0_15320 <= _zz_dataOut_payload_0_15176;
    _zz_dataOut_payload_0_15321 <= _zz_dataOut_payload_0_15177;
    _zz_dataOut_payload_0_15322 <= _zz_dataOut_payload_0_15178;
    _zz_dataOut_payload_0_15323 <= _zz_dataOut_payload_0_15179;
    _zz_dataOut_payload_0_15324 <= _zz_dataOut_payload_0_15180;
    _zz_dataOut_payload_0_15325 <= _zz_dataOut_payload_0_15181;
    _zz_dataOut_payload_0_15326 <= _zz_dataOut_payload_0_15182;
    _zz_dataOut_payload_0_15327 <= _zz_dataOut_payload_0_15183;
    _zz_dataOut_payload_0_15328 <= _zz_dataOut_payload_0_15296;
    _zz_dataOut_payload_0_15329 <= _zz_dataOut_payload_0_15297;
    _zz_dataOut_payload_0_15330 <= _zz_dataOut_payload_0_15298;
    _zz_dataOut_payload_0_15331 <= _zz_dataOut_payload_0_15299;
    _zz_dataOut_payload_0_15332 <= _zz_dataOut_payload_0_15300;
    _zz_dataOut_payload_0_15333 <= _zz_dataOut_payload_0_15301;
    _zz_dataOut_payload_0_15334 <= _zz_dataOut_payload_0_15302;
    _zz_dataOut_payload_0_15335 <= _zz_dataOut_payload_0_15303;
    _zz_dataOut_payload_0_15336 <= _zz_dataOut_payload_0_15304;
    _zz_dataOut_payload_0_15337 <= _zz_dataOut_payload_0_15305;
    _zz_dataOut_payload_0_15338 <= _zz_dataOut_payload_0_15306;
    _zz_dataOut_payload_0_15339 <= _zz_dataOut_payload_0_15307;
    _zz_dataOut_payload_0_15340 <= _zz_dataOut_payload_0_15308;
    _zz_dataOut_payload_0_15341 <= _zz_dataOut_payload_0_15309;
    _zz_dataOut_payload_0_15342 <= _zz_dataOut_payload_0_15310;
    _zz_dataOut_payload_0_15343 <= _zz_dataOut_payload_0_15311;
    _zz_dataOut_payload_0_15436 <= (_zz_dataOut_payload_0_15434 ? _zz_dataOut_payload_0_15429 : _zz_dataOut_payload_0_15432);
    _zz_dataOut_payload_0_15437 <= (_zz_dataOut_payload_0_15434 ? _zz_dataOut_payload_0_15432 : _zz_dataOut_payload_0_15429);
    _zz_dataOut_payload_0_15438 <= (_zz_dataOut_payload_0_15435 ? _zz_dataOut_payload_0_15430 : _zz_dataOut_payload_0_15433);
    _zz_dataOut_payload_0_15439 <= (_zz_dataOut_payload_0_15435 ? _zz_dataOut_payload_0_15433 : _zz_dataOut_payload_0_15430);
    _zz_dataOut_payload_0_15448 <= (_zz_dataOut_payload_0_15446 ? _zz_dataOut_payload_0_15441 : _zz_dataOut_payload_0_15444);
    _zz_dataOut_payload_0_15449 <= (_zz_dataOut_payload_0_15446 ? _zz_dataOut_payload_0_15444 : _zz_dataOut_payload_0_15441);
    _zz_dataOut_payload_0_15450 <= (_zz_dataOut_payload_0_15447 ? _zz_dataOut_payload_0_15442 : _zz_dataOut_payload_0_15445);
    _zz_dataOut_payload_0_15451 <= (_zz_dataOut_payload_0_15447 ? _zz_dataOut_payload_0_15445 : _zz_dataOut_payload_0_15442);
    _zz_dataOut_payload_0_15452 <= _zz_dataOut_payload_0_15436;
    _zz_dataOut_payload_0_15453 <= _zz_dataOut_payload_0_15437;
    _zz_dataOut_payload_0_15454 <= _zz_dataOut_payload_0_15438;
    _zz_dataOut_payload_0_15455 <= _zz_dataOut_payload_0_15439;
    _zz_dataOut_payload_0_15456 <= _zz_dataOut_payload_0_15448;
    _zz_dataOut_payload_0_15457 <= _zz_dataOut_payload_0_15449;
    _zz_dataOut_payload_0_15458 <= _zz_dataOut_payload_0_15450;
    _zz_dataOut_payload_0_15459 <= _zz_dataOut_payload_0_15451;
    _zz_dataOut_payload_0_15480 <= (_zz_dataOut_payload_0_15478 ? _zz_dataOut_payload_0_15473 : _zz_dataOut_payload_0_15476);
    _zz_dataOut_payload_0_15481 <= (_zz_dataOut_payload_0_15478 ? _zz_dataOut_payload_0_15476 : _zz_dataOut_payload_0_15473);
    _zz_dataOut_payload_0_15482 <= (_zz_dataOut_payload_0_15479 ? _zz_dataOut_payload_0_15474 : _zz_dataOut_payload_0_15477);
    _zz_dataOut_payload_0_15483 <= (_zz_dataOut_payload_0_15479 ? _zz_dataOut_payload_0_15477 : _zz_dataOut_payload_0_15474);
    _zz_dataOut_payload_0_15492 <= (_zz_dataOut_payload_0_15490 ? _zz_dataOut_payload_0_15485 : _zz_dataOut_payload_0_15488);
    _zz_dataOut_payload_0_15493 <= (_zz_dataOut_payload_0_15490 ? _zz_dataOut_payload_0_15488 : _zz_dataOut_payload_0_15485);
    _zz_dataOut_payload_0_15494 <= (_zz_dataOut_payload_0_15491 ? _zz_dataOut_payload_0_15486 : _zz_dataOut_payload_0_15489);
    _zz_dataOut_payload_0_15495 <= (_zz_dataOut_payload_0_15491 ? _zz_dataOut_payload_0_15489 : _zz_dataOut_payload_0_15486);
    _zz_dataOut_payload_0_15496 <= _zz_dataOut_payload_0_15480;
    _zz_dataOut_payload_0_15497 <= _zz_dataOut_payload_0_15481;
    _zz_dataOut_payload_0_15498 <= _zz_dataOut_payload_0_15482;
    _zz_dataOut_payload_0_15499 <= _zz_dataOut_payload_0_15483;
    _zz_dataOut_payload_0_15500 <= _zz_dataOut_payload_0_15492;
    _zz_dataOut_payload_0_15501 <= _zz_dataOut_payload_0_15493;
    _zz_dataOut_payload_0_15502 <= _zz_dataOut_payload_0_15494;
    _zz_dataOut_payload_0_15503 <= _zz_dataOut_payload_0_15495;
    _zz_dataOut_payload_0_15504 <= _zz_dataOut_payload_0_15452;
    _zz_dataOut_payload_0_15505 <= _zz_dataOut_payload_0_15453;
    _zz_dataOut_payload_0_15506 <= _zz_dataOut_payload_0_15454;
    _zz_dataOut_payload_0_15507 <= _zz_dataOut_payload_0_15455;
    _zz_dataOut_payload_0_15508 <= _zz_dataOut_payload_0_15456;
    _zz_dataOut_payload_0_15509 <= _zz_dataOut_payload_0_15457;
    _zz_dataOut_payload_0_15510 <= _zz_dataOut_payload_0_15458;
    _zz_dataOut_payload_0_15511 <= _zz_dataOut_payload_0_15459;
    _zz_dataOut_payload_0_15512 <= _zz_dataOut_payload_0_15496;
    _zz_dataOut_payload_0_15513 <= _zz_dataOut_payload_0_15497;
    _zz_dataOut_payload_0_15514 <= _zz_dataOut_payload_0_15498;
    _zz_dataOut_payload_0_15515 <= _zz_dataOut_payload_0_15499;
    _zz_dataOut_payload_0_15516 <= _zz_dataOut_payload_0_15500;
    _zz_dataOut_payload_0_15517 <= _zz_dataOut_payload_0_15501;
    _zz_dataOut_payload_0_15518 <= _zz_dataOut_payload_0_15502;
    _zz_dataOut_payload_0_15519 <= _zz_dataOut_payload_0_15503;
    _zz_dataOut_payload_0_15564 <= (_zz_dataOut_payload_0_15562 ? _zz_dataOut_payload_0_15557 : _zz_dataOut_payload_0_15560);
    _zz_dataOut_payload_0_15565 <= (_zz_dataOut_payload_0_15562 ? _zz_dataOut_payload_0_15560 : _zz_dataOut_payload_0_15557);
    _zz_dataOut_payload_0_15566 <= (_zz_dataOut_payload_0_15563 ? _zz_dataOut_payload_0_15558 : _zz_dataOut_payload_0_15561);
    _zz_dataOut_payload_0_15567 <= (_zz_dataOut_payload_0_15563 ? _zz_dataOut_payload_0_15561 : _zz_dataOut_payload_0_15558);
    _zz_dataOut_payload_0_15576 <= (_zz_dataOut_payload_0_15574 ? _zz_dataOut_payload_0_15569 : _zz_dataOut_payload_0_15572);
    _zz_dataOut_payload_0_15577 <= (_zz_dataOut_payload_0_15574 ? _zz_dataOut_payload_0_15572 : _zz_dataOut_payload_0_15569);
    _zz_dataOut_payload_0_15578 <= (_zz_dataOut_payload_0_15575 ? _zz_dataOut_payload_0_15570 : _zz_dataOut_payload_0_15573);
    _zz_dataOut_payload_0_15579 <= (_zz_dataOut_payload_0_15575 ? _zz_dataOut_payload_0_15573 : _zz_dataOut_payload_0_15570);
    _zz_dataOut_payload_0_15580 <= _zz_dataOut_payload_0_15564;
    _zz_dataOut_payload_0_15581 <= _zz_dataOut_payload_0_15565;
    _zz_dataOut_payload_0_15582 <= _zz_dataOut_payload_0_15566;
    _zz_dataOut_payload_0_15583 <= _zz_dataOut_payload_0_15567;
    _zz_dataOut_payload_0_15584 <= _zz_dataOut_payload_0_15576;
    _zz_dataOut_payload_0_15585 <= _zz_dataOut_payload_0_15577;
    _zz_dataOut_payload_0_15586 <= _zz_dataOut_payload_0_15578;
    _zz_dataOut_payload_0_15587 <= _zz_dataOut_payload_0_15579;
    _zz_dataOut_payload_0_15608 <= (_zz_dataOut_payload_0_15606 ? _zz_dataOut_payload_0_15601 : _zz_dataOut_payload_0_15604);
    _zz_dataOut_payload_0_15609 <= (_zz_dataOut_payload_0_15606 ? _zz_dataOut_payload_0_15604 : _zz_dataOut_payload_0_15601);
    _zz_dataOut_payload_0_15610 <= (_zz_dataOut_payload_0_15607 ? _zz_dataOut_payload_0_15602 : _zz_dataOut_payload_0_15605);
    _zz_dataOut_payload_0_15611 <= (_zz_dataOut_payload_0_15607 ? _zz_dataOut_payload_0_15605 : _zz_dataOut_payload_0_15602);
    _zz_dataOut_payload_0_15620 <= (_zz_dataOut_payload_0_15618 ? _zz_dataOut_payload_0_15613 : _zz_dataOut_payload_0_15616);
    _zz_dataOut_payload_0_15621 <= (_zz_dataOut_payload_0_15618 ? _zz_dataOut_payload_0_15616 : _zz_dataOut_payload_0_15613);
    _zz_dataOut_payload_0_15622 <= (_zz_dataOut_payload_0_15619 ? _zz_dataOut_payload_0_15614 : _zz_dataOut_payload_0_15617);
    _zz_dataOut_payload_0_15623 <= (_zz_dataOut_payload_0_15619 ? _zz_dataOut_payload_0_15617 : _zz_dataOut_payload_0_15614);
    _zz_dataOut_payload_0_15624 <= _zz_dataOut_payload_0_15608;
    _zz_dataOut_payload_0_15625 <= _zz_dataOut_payload_0_15609;
    _zz_dataOut_payload_0_15626 <= _zz_dataOut_payload_0_15610;
    _zz_dataOut_payload_0_15627 <= _zz_dataOut_payload_0_15611;
    _zz_dataOut_payload_0_15628 <= _zz_dataOut_payload_0_15620;
    _zz_dataOut_payload_0_15629 <= _zz_dataOut_payload_0_15621;
    _zz_dataOut_payload_0_15630 <= _zz_dataOut_payload_0_15622;
    _zz_dataOut_payload_0_15631 <= _zz_dataOut_payload_0_15623;
    _zz_dataOut_payload_0_15632 <= _zz_dataOut_payload_0_15580;
    _zz_dataOut_payload_0_15633 <= _zz_dataOut_payload_0_15581;
    _zz_dataOut_payload_0_15634 <= _zz_dataOut_payload_0_15582;
    _zz_dataOut_payload_0_15635 <= _zz_dataOut_payload_0_15583;
    _zz_dataOut_payload_0_15636 <= _zz_dataOut_payload_0_15584;
    _zz_dataOut_payload_0_15637 <= _zz_dataOut_payload_0_15585;
    _zz_dataOut_payload_0_15638 <= _zz_dataOut_payload_0_15586;
    _zz_dataOut_payload_0_15639 <= _zz_dataOut_payload_0_15587;
    _zz_dataOut_payload_0_15640 <= _zz_dataOut_payload_0_15624;
    _zz_dataOut_payload_0_15641 <= _zz_dataOut_payload_0_15625;
    _zz_dataOut_payload_0_15642 <= _zz_dataOut_payload_0_15626;
    _zz_dataOut_payload_0_15643 <= _zz_dataOut_payload_0_15627;
    _zz_dataOut_payload_0_15644 <= _zz_dataOut_payload_0_15628;
    _zz_dataOut_payload_0_15645 <= _zz_dataOut_payload_0_15629;
    _zz_dataOut_payload_0_15646 <= _zz_dataOut_payload_0_15630;
    _zz_dataOut_payload_0_15647 <= _zz_dataOut_payload_0_15631;
    _zz_dataOut_payload_0_15648 <= _zz_dataOut_payload_0_15504;
    _zz_dataOut_payload_0_15649 <= _zz_dataOut_payload_0_15505;
    _zz_dataOut_payload_0_15650 <= _zz_dataOut_payload_0_15506;
    _zz_dataOut_payload_0_15651 <= _zz_dataOut_payload_0_15507;
    _zz_dataOut_payload_0_15652 <= _zz_dataOut_payload_0_15508;
    _zz_dataOut_payload_0_15653 <= _zz_dataOut_payload_0_15509;
    _zz_dataOut_payload_0_15654 <= _zz_dataOut_payload_0_15510;
    _zz_dataOut_payload_0_15655 <= _zz_dataOut_payload_0_15511;
    _zz_dataOut_payload_0_15656 <= _zz_dataOut_payload_0_15512;
    _zz_dataOut_payload_0_15657 <= _zz_dataOut_payload_0_15513;
    _zz_dataOut_payload_0_15658 <= _zz_dataOut_payload_0_15514;
    _zz_dataOut_payload_0_15659 <= _zz_dataOut_payload_0_15515;
    _zz_dataOut_payload_0_15660 <= _zz_dataOut_payload_0_15516;
    _zz_dataOut_payload_0_15661 <= _zz_dataOut_payload_0_15517;
    _zz_dataOut_payload_0_15662 <= _zz_dataOut_payload_0_15518;
    _zz_dataOut_payload_0_15663 <= _zz_dataOut_payload_0_15519;
    _zz_dataOut_payload_0_15664 <= _zz_dataOut_payload_0_15632;
    _zz_dataOut_payload_0_15665 <= _zz_dataOut_payload_0_15633;
    _zz_dataOut_payload_0_15666 <= _zz_dataOut_payload_0_15634;
    _zz_dataOut_payload_0_15667 <= _zz_dataOut_payload_0_15635;
    _zz_dataOut_payload_0_15668 <= _zz_dataOut_payload_0_15636;
    _zz_dataOut_payload_0_15669 <= _zz_dataOut_payload_0_15637;
    _zz_dataOut_payload_0_15670 <= _zz_dataOut_payload_0_15638;
    _zz_dataOut_payload_0_15671 <= _zz_dataOut_payload_0_15639;
    _zz_dataOut_payload_0_15672 <= _zz_dataOut_payload_0_15640;
    _zz_dataOut_payload_0_15673 <= _zz_dataOut_payload_0_15641;
    _zz_dataOut_payload_0_15674 <= _zz_dataOut_payload_0_15642;
    _zz_dataOut_payload_0_15675 <= _zz_dataOut_payload_0_15643;
    _zz_dataOut_payload_0_15676 <= _zz_dataOut_payload_0_15644;
    _zz_dataOut_payload_0_15677 <= _zz_dataOut_payload_0_15645;
    _zz_dataOut_payload_0_15678 <= _zz_dataOut_payload_0_15646;
    _zz_dataOut_payload_0_15679 <= _zz_dataOut_payload_0_15647;
    _zz_dataOut_payload_0_15680 <= _zz_dataOut_payload_0_15312;
    _zz_dataOut_payload_0_15681 <= _zz_dataOut_payload_0_15313;
    _zz_dataOut_payload_0_15682 <= _zz_dataOut_payload_0_15314;
    _zz_dataOut_payload_0_15683 <= _zz_dataOut_payload_0_15315;
    _zz_dataOut_payload_0_15684 <= _zz_dataOut_payload_0_15316;
    _zz_dataOut_payload_0_15685 <= _zz_dataOut_payload_0_15317;
    _zz_dataOut_payload_0_15686 <= _zz_dataOut_payload_0_15318;
    _zz_dataOut_payload_0_15687 <= _zz_dataOut_payload_0_15319;
    _zz_dataOut_payload_0_15688 <= _zz_dataOut_payload_0_15320;
    _zz_dataOut_payload_0_15689 <= _zz_dataOut_payload_0_15321;
    _zz_dataOut_payload_0_15690 <= _zz_dataOut_payload_0_15322;
    _zz_dataOut_payload_0_15691 <= _zz_dataOut_payload_0_15323;
    _zz_dataOut_payload_0_15692 <= _zz_dataOut_payload_0_15324;
    _zz_dataOut_payload_0_15693 <= _zz_dataOut_payload_0_15325;
    _zz_dataOut_payload_0_15694 <= _zz_dataOut_payload_0_15326;
    _zz_dataOut_payload_0_15695 <= _zz_dataOut_payload_0_15327;
    _zz_dataOut_payload_0_15696 <= _zz_dataOut_payload_0_15328;
    _zz_dataOut_payload_0_15697 <= _zz_dataOut_payload_0_15329;
    _zz_dataOut_payload_0_15698 <= _zz_dataOut_payload_0_15330;
    _zz_dataOut_payload_0_15699 <= _zz_dataOut_payload_0_15331;
    _zz_dataOut_payload_0_15700 <= _zz_dataOut_payload_0_15332;
    _zz_dataOut_payload_0_15701 <= _zz_dataOut_payload_0_15333;
    _zz_dataOut_payload_0_15702 <= _zz_dataOut_payload_0_15334;
    _zz_dataOut_payload_0_15703 <= _zz_dataOut_payload_0_15335;
    _zz_dataOut_payload_0_15704 <= _zz_dataOut_payload_0_15336;
    _zz_dataOut_payload_0_15705 <= _zz_dataOut_payload_0_15337;
    _zz_dataOut_payload_0_15706 <= _zz_dataOut_payload_0_15338;
    _zz_dataOut_payload_0_15707 <= _zz_dataOut_payload_0_15339;
    _zz_dataOut_payload_0_15708 <= _zz_dataOut_payload_0_15340;
    _zz_dataOut_payload_0_15709 <= _zz_dataOut_payload_0_15341;
    _zz_dataOut_payload_0_15710 <= _zz_dataOut_payload_0_15342;
    _zz_dataOut_payload_0_15711 <= _zz_dataOut_payload_0_15343;
    _zz_dataOut_payload_0_15712 <= _zz_dataOut_payload_0_15648;
    _zz_dataOut_payload_0_15713 <= _zz_dataOut_payload_0_15649;
    _zz_dataOut_payload_0_15714 <= _zz_dataOut_payload_0_15650;
    _zz_dataOut_payload_0_15715 <= _zz_dataOut_payload_0_15651;
    _zz_dataOut_payload_0_15716 <= _zz_dataOut_payload_0_15652;
    _zz_dataOut_payload_0_15717 <= _zz_dataOut_payload_0_15653;
    _zz_dataOut_payload_0_15718 <= _zz_dataOut_payload_0_15654;
    _zz_dataOut_payload_0_15719 <= _zz_dataOut_payload_0_15655;
    _zz_dataOut_payload_0_15720 <= _zz_dataOut_payload_0_15656;
    _zz_dataOut_payload_0_15721 <= _zz_dataOut_payload_0_15657;
    _zz_dataOut_payload_0_15722 <= _zz_dataOut_payload_0_15658;
    _zz_dataOut_payload_0_15723 <= _zz_dataOut_payload_0_15659;
    _zz_dataOut_payload_0_15724 <= _zz_dataOut_payload_0_15660;
    _zz_dataOut_payload_0_15725 <= _zz_dataOut_payload_0_15661;
    _zz_dataOut_payload_0_15726 <= _zz_dataOut_payload_0_15662;
    _zz_dataOut_payload_0_15727 <= _zz_dataOut_payload_0_15663;
    _zz_dataOut_payload_0_15728 <= _zz_dataOut_payload_0_15664;
    _zz_dataOut_payload_0_15729 <= _zz_dataOut_payload_0_15665;
    _zz_dataOut_payload_0_15730 <= _zz_dataOut_payload_0_15666;
    _zz_dataOut_payload_0_15731 <= _zz_dataOut_payload_0_15667;
    _zz_dataOut_payload_0_15732 <= _zz_dataOut_payload_0_15668;
    _zz_dataOut_payload_0_15733 <= _zz_dataOut_payload_0_15669;
    _zz_dataOut_payload_0_15734 <= _zz_dataOut_payload_0_15670;
    _zz_dataOut_payload_0_15735 <= _zz_dataOut_payload_0_15671;
    _zz_dataOut_payload_0_15736 <= _zz_dataOut_payload_0_15672;
    _zz_dataOut_payload_0_15737 <= _zz_dataOut_payload_0_15673;
    _zz_dataOut_payload_0_15738 <= _zz_dataOut_payload_0_15674;
    _zz_dataOut_payload_0_15739 <= _zz_dataOut_payload_0_15675;
    _zz_dataOut_payload_0_15740 <= _zz_dataOut_payload_0_15676;
    _zz_dataOut_payload_0_15741 <= _zz_dataOut_payload_0_15677;
    _zz_dataOut_payload_0_15742 <= _zz_dataOut_payload_0_15678;
    _zz_dataOut_payload_0_15743 <= _zz_dataOut_payload_0_15679;
    _zz_dataOut_payload_0_15744 <= _zz_dataOut_payload_0_14848;
    _zz_dataOut_payload_0_15745 <= _zz_dataOut_payload_0_14849;
    _zz_dataOut_payload_0_15746 <= _zz_dataOut_payload_0_14850;
    _zz_dataOut_payload_0_15747 <= _zz_dataOut_payload_0_14851;
    _zz_dataOut_payload_0_15748 <= _zz_dataOut_payload_0_14852;
    _zz_dataOut_payload_0_15749 <= _zz_dataOut_payload_0_14853;
    _zz_dataOut_payload_0_15750 <= _zz_dataOut_payload_0_14854;
    _zz_dataOut_payload_0_15751 <= _zz_dataOut_payload_0_14855;
    _zz_dataOut_payload_0_15752 <= _zz_dataOut_payload_0_14856;
    _zz_dataOut_payload_0_15753 <= _zz_dataOut_payload_0_14857;
    _zz_dataOut_payload_0_15754 <= _zz_dataOut_payload_0_14858;
    _zz_dataOut_payload_0_15755 <= _zz_dataOut_payload_0_14859;
    _zz_dataOut_payload_0_15756 <= _zz_dataOut_payload_0_14860;
    _zz_dataOut_payload_0_15757 <= _zz_dataOut_payload_0_14861;
    _zz_dataOut_payload_0_15758 <= _zz_dataOut_payload_0_14862;
    _zz_dataOut_payload_0_15759 <= _zz_dataOut_payload_0_14863;
    _zz_dataOut_payload_0_15760 <= _zz_dataOut_payload_0_14864;
    _zz_dataOut_payload_0_15761 <= _zz_dataOut_payload_0_14865;
    _zz_dataOut_payload_0_15762 <= _zz_dataOut_payload_0_14866;
    _zz_dataOut_payload_0_15763 <= _zz_dataOut_payload_0_14867;
    _zz_dataOut_payload_0_15764 <= _zz_dataOut_payload_0_14868;
    _zz_dataOut_payload_0_15765 <= _zz_dataOut_payload_0_14869;
    _zz_dataOut_payload_0_15766 <= _zz_dataOut_payload_0_14870;
    _zz_dataOut_payload_0_15767 <= _zz_dataOut_payload_0_14871;
    _zz_dataOut_payload_0_15768 <= _zz_dataOut_payload_0_14872;
    _zz_dataOut_payload_0_15769 <= _zz_dataOut_payload_0_14873;
    _zz_dataOut_payload_0_15770 <= _zz_dataOut_payload_0_14874;
    _zz_dataOut_payload_0_15771 <= _zz_dataOut_payload_0_14875;
    _zz_dataOut_payload_0_15772 <= _zz_dataOut_payload_0_14876;
    _zz_dataOut_payload_0_15773 <= _zz_dataOut_payload_0_14877;
    _zz_dataOut_payload_0_15774 <= _zz_dataOut_payload_0_14878;
    _zz_dataOut_payload_0_15775 <= _zz_dataOut_payload_0_14879;
    _zz_dataOut_payload_0_15776 <= _zz_dataOut_payload_0_14880;
    _zz_dataOut_payload_0_15777 <= _zz_dataOut_payload_0_14881;
    _zz_dataOut_payload_0_15778 <= _zz_dataOut_payload_0_14882;
    _zz_dataOut_payload_0_15779 <= _zz_dataOut_payload_0_14883;
    _zz_dataOut_payload_0_15780 <= _zz_dataOut_payload_0_14884;
    _zz_dataOut_payload_0_15781 <= _zz_dataOut_payload_0_14885;
    _zz_dataOut_payload_0_15782 <= _zz_dataOut_payload_0_14886;
    _zz_dataOut_payload_0_15783 <= _zz_dataOut_payload_0_14887;
    _zz_dataOut_payload_0_15784 <= _zz_dataOut_payload_0_14888;
    _zz_dataOut_payload_0_15785 <= _zz_dataOut_payload_0_14889;
    _zz_dataOut_payload_0_15786 <= _zz_dataOut_payload_0_14890;
    _zz_dataOut_payload_0_15787 <= _zz_dataOut_payload_0_14891;
    _zz_dataOut_payload_0_15788 <= _zz_dataOut_payload_0_14892;
    _zz_dataOut_payload_0_15789 <= _zz_dataOut_payload_0_14893;
    _zz_dataOut_payload_0_15790 <= _zz_dataOut_payload_0_14894;
    _zz_dataOut_payload_0_15791 <= _zz_dataOut_payload_0_14895;
    _zz_dataOut_payload_0_15792 <= _zz_dataOut_payload_0_14896;
    _zz_dataOut_payload_0_15793 <= _zz_dataOut_payload_0_14897;
    _zz_dataOut_payload_0_15794 <= _zz_dataOut_payload_0_14898;
    _zz_dataOut_payload_0_15795 <= _zz_dataOut_payload_0_14899;
    _zz_dataOut_payload_0_15796 <= _zz_dataOut_payload_0_14900;
    _zz_dataOut_payload_0_15797 <= _zz_dataOut_payload_0_14901;
    _zz_dataOut_payload_0_15798 <= _zz_dataOut_payload_0_14902;
    _zz_dataOut_payload_0_15799 <= _zz_dataOut_payload_0_14903;
    _zz_dataOut_payload_0_15800 <= _zz_dataOut_payload_0_14904;
    _zz_dataOut_payload_0_15801 <= _zz_dataOut_payload_0_14905;
    _zz_dataOut_payload_0_15802 <= _zz_dataOut_payload_0_14906;
    _zz_dataOut_payload_0_15803 <= _zz_dataOut_payload_0_14907;
    _zz_dataOut_payload_0_15804 <= _zz_dataOut_payload_0_14908;
    _zz_dataOut_payload_0_15805 <= _zz_dataOut_payload_0_14909;
    _zz_dataOut_payload_0_15806 <= _zz_dataOut_payload_0_14910;
    _zz_dataOut_payload_0_15807 <= _zz_dataOut_payload_0_14911;
    _zz_dataOut_payload_0_15808 <= _zz_dataOut_payload_0_15680;
    _zz_dataOut_payload_0_15809 <= _zz_dataOut_payload_0_15681;
    _zz_dataOut_payload_0_15810 <= _zz_dataOut_payload_0_15682;
    _zz_dataOut_payload_0_15811 <= _zz_dataOut_payload_0_15683;
    _zz_dataOut_payload_0_15812 <= _zz_dataOut_payload_0_15684;
    _zz_dataOut_payload_0_15813 <= _zz_dataOut_payload_0_15685;
    _zz_dataOut_payload_0_15814 <= _zz_dataOut_payload_0_15686;
    _zz_dataOut_payload_0_15815 <= _zz_dataOut_payload_0_15687;
    _zz_dataOut_payload_0_15816 <= _zz_dataOut_payload_0_15688;
    _zz_dataOut_payload_0_15817 <= _zz_dataOut_payload_0_15689;
    _zz_dataOut_payload_0_15818 <= _zz_dataOut_payload_0_15690;
    _zz_dataOut_payload_0_15819 <= _zz_dataOut_payload_0_15691;
    _zz_dataOut_payload_0_15820 <= _zz_dataOut_payload_0_15692;
    _zz_dataOut_payload_0_15821 <= _zz_dataOut_payload_0_15693;
    _zz_dataOut_payload_0_15822 <= _zz_dataOut_payload_0_15694;
    _zz_dataOut_payload_0_15823 <= _zz_dataOut_payload_0_15695;
    _zz_dataOut_payload_0_15824 <= _zz_dataOut_payload_0_15696;
    _zz_dataOut_payload_0_15825 <= _zz_dataOut_payload_0_15697;
    _zz_dataOut_payload_0_15826 <= _zz_dataOut_payload_0_15698;
    _zz_dataOut_payload_0_15827 <= _zz_dataOut_payload_0_15699;
    _zz_dataOut_payload_0_15828 <= _zz_dataOut_payload_0_15700;
    _zz_dataOut_payload_0_15829 <= _zz_dataOut_payload_0_15701;
    _zz_dataOut_payload_0_15830 <= _zz_dataOut_payload_0_15702;
    _zz_dataOut_payload_0_15831 <= _zz_dataOut_payload_0_15703;
    _zz_dataOut_payload_0_15832 <= _zz_dataOut_payload_0_15704;
    _zz_dataOut_payload_0_15833 <= _zz_dataOut_payload_0_15705;
    _zz_dataOut_payload_0_15834 <= _zz_dataOut_payload_0_15706;
    _zz_dataOut_payload_0_15835 <= _zz_dataOut_payload_0_15707;
    _zz_dataOut_payload_0_15836 <= _zz_dataOut_payload_0_15708;
    _zz_dataOut_payload_0_15837 <= _zz_dataOut_payload_0_15709;
    _zz_dataOut_payload_0_15838 <= _zz_dataOut_payload_0_15710;
    _zz_dataOut_payload_0_15839 <= _zz_dataOut_payload_0_15711;
    _zz_dataOut_payload_0_15840 <= _zz_dataOut_payload_0_15712;
    _zz_dataOut_payload_0_15841 <= _zz_dataOut_payload_0_15713;
    _zz_dataOut_payload_0_15842 <= _zz_dataOut_payload_0_15714;
    _zz_dataOut_payload_0_15843 <= _zz_dataOut_payload_0_15715;
    _zz_dataOut_payload_0_15844 <= _zz_dataOut_payload_0_15716;
    _zz_dataOut_payload_0_15845 <= _zz_dataOut_payload_0_15717;
    _zz_dataOut_payload_0_15846 <= _zz_dataOut_payload_0_15718;
    _zz_dataOut_payload_0_15847 <= _zz_dataOut_payload_0_15719;
    _zz_dataOut_payload_0_15848 <= _zz_dataOut_payload_0_15720;
    _zz_dataOut_payload_0_15849 <= _zz_dataOut_payload_0_15721;
    _zz_dataOut_payload_0_15850 <= _zz_dataOut_payload_0_15722;
    _zz_dataOut_payload_0_15851 <= _zz_dataOut_payload_0_15723;
    _zz_dataOut_payload_0_15852 <= _zz_dataOut_payload_0_15724;
    _zz_dataOut_payload_0_15853 <= _zz_dataOut_payload_0_15725;
    _zz_dataOut_payload_0_15854 <= _zz_dataOut_payload_0_15726;
    _zz_dataOut_payload_0_15855 <= _zz_dataOut_payload_0_15727;
    _zz_dataOut_payload_0_15856 <= _zz_dataOut_payload_0_15728;
    _zz_dataOut_payload_0_15857 <= _zz_dataOut_payload_0_15729;
    _zz_dataOut_payload_0_15858 <= _zz_dataOut_payload_0_15730;
    _zz_dataOut_payload_0_15859 <= _zz_dataOut_payload_0_15731;
    _zz_dataOut_payload_0_15860 <= _zz_dataOut_payload_0_15732;
    _zz_dataOut_payload_0_15861 <= _zz_dataOut_payload_0_15733;
    _zz_dataOut_payload_0_15862 <= _zz_dataOut_payload_0_15734;
    _zz_dataOut_payload_0_15863 <= _zz_dataOut_payload_0_15735;
    _zz_dataOut_payload_0_15864 <= _zz_dataOut_payload_0_15736;
    _zz_dataOut_payload_0_15865 <= _zz_dataOut_payload_0_15737;
    _zz_dataOut_payload_0_15866 <= _zz_dataOut_payload_0_15738;
    _zz_dataOut_payload_0_15867 <= _zz_dataOut_payload_0_15739;
    _zz_dataOut_payload_0_15868 <= _zz_dataOut_payload_0_15740;
    _zz_dataOut_payload_0_15869 <= _zz_dataOut_payload_0_15741;
    _zz_dataOut_payload_0_15870 <= _zz_dataOut_payload_0_15742;
    _zz_dataOut_payload_0_15871 <= _zz_dataOut_payload_0_15743;
    _zz_dataOut_payload_0_15872 <= _zz_dataOut_payload_0_13760;
    _zz_dataOut_payload_0_15873 <= _zz_dataOut_payload_0_13761;
    _zz_dataOut_payload_0_15874 <= _zz_dataOut_payload_0_13762;
    _zz_dataOut_payload_0_15875 <= _zz_dataOut_payload_0_13763;
    _zz_dataOut_payload_0_15876 <= _zz_dataOut_payload_0_13764;
    _zz_dataOut_payload_0_15877 <= _zz_dataOut_payload_0_13765;
    _zz_dataOut_payload_0_15878 <= _zz_dataOut_payload_0_13766;
    _zz_dataOut_payload_0_15879 <= _zz_dataOut_payload_0_13767;
    _zz_dataOut_payload_0_15880 <= _zz_dataOut_payload_0_13768;
    _zz_dataOut_payload_0_15881 <= _zz_dataOut_payload_0_13769;
    _zz_dataOut_payload_0_15882 <= _zz_dataOut_payload_0_13770;
    _zz_dataOut_payload_0_15883 <= _zz_dataOut_payload_0_13771;
    _zz_dataOut_payload_0_15884 <= _zz_dataOut_payload_0_13772;
    _zz_dataOut_payload_0_15885 <= _zz_dataOut_payload_0_13773;
    _zz_dataOut_payload_0_15886 <= _zz_dataOut_payload_0_13774;
    _zz_dataOut_payload_0_15887 <= _zz_dataOut_payload_0_13775;
    _zz_dataOut_payload_0_15888 <= _zz_dataOut_payload_0_13776;
    _zz_dataOut_payload_0_15889 <= _zz_dataOut_payload_0_13777;
    _zz_dataOut_payload_0_15890 <= _zz_dataOut_payload_0_13778;
    _zz_dataOut_payload_0_15891 <= _zz_dataOut_payload_0_13779;
    _zz_dataOut_payload_0_15892 <= _zz_dataOut_payload_0_13780;
    _zz_dataOut_payload_0_15893 <= _zz_dataOut_payload_0_13781;
    _zz_dataOut_payload_0_15894 <= _zz_dataOut_payload_0_13782;
    _zz_dataOut_payload_0_15895 <= _zz_dataOut_payload_0_13783;
    _zz_dataOut_payload_0_15896 <= _zz_dataOut_payload_0_13784;
    _zz_dataOut_payload_0_15897 <= _zz_dataOut_payload_0_13785;
    _zz_dataOut_payload_0_15898 <= _zz_dataOut_payload_0_13786;
    _zz_dataOut_payload_0_15899 <= _zz_dataOut_payload_0_13787;
    _zz_dataOut_payload_0_15900 <= _zz_dataOut_payload_0_13788;
    _zz_dataOut_payload_0_15901 <= _zz_dataOut_payload_0_13789;
    _zz_dataOut_payload_0_15902 <= _zz_dataOut_payload_0_13790;
    _zz_dataOut_payload_0_15903 <= _zz_dataOut_payload_0_13791;
    _zz_dataOut_payload_0_15904 <= _zz_dataOut_payload_0_13792;
    _zz_dataOut_payload_0_15905 <= _zz_dataOut_payload_0_13793;
    _zz_dataOut_payload_0_15906 <= _zz_dataOut_payload_0_13794;
    _zz_dataOut_payload_0_15907 <= _zz_dataOut_payload_0_13795;
    _zz_dataOut_payload_0_15908 <= _zz_dataOut_payload_0_13796;
    _zz_dataOut_payload_0_15909 <= _zz_dataOut_payload_0_13797;
    _zz_dataOut_payload_0_15910 <= _zz_dataOut_payload_0_13798;
    _zz_dataOut_payload_0_15911 <= _zz_dataOut_payload_0_13799;
    _zz_dataOut_payload_0_15912 <= _zz_dataOut_payload_0_13800;
    _zz_dataOut_payload_0_15913 <= _zz_dataOut_payload_0_13801;
    _zz_dataOut_payload_0_15914 <= _zz_dataOut_payload_0_13802;
    _zz_dataOut_payload_0_15915 <= _zz_dataOut_payload_0_13803;
    _zz_dataOut_payload_0_15916 <= _zz_dataOut_payload_0_13804;
    _zz_dataOut_payload_0_15917 <= _zz_dataOut_payload_0_13805;
    _zz_dataOut_payload_0_15918 <= _zz_dataOut_payload_0_13806;
    _zz_dataOut_payload_0_15919 <= _zz_dataOut_payload_0_13807;
    _zz_dataOut_payload_0_15920 <= _zz_dataOut_payload_0_13808;
    _zz_dataOut_payload_0_15921 <= _zz_dataOut_payload_0_13809;
    _zz_dataOut_payload_0_15922 <= _zz_dataOut_payload_0_13810;
    _zz_dataOut_payload_0_15923 <= _zz_dataOut_payload_0_13811;
    _zz_dataOut_payload_0_15924 <= _zz_dataOut_payload_0_13812;
    _zz_dataOut_payload_0_15925 <= _zz_dataOut_payload_0_13813;
    _zz_dataOut_payload_0_15926 <= _zz_dataOut_payload_0_13814;
    _zz_dataOut_payload_0_15927 <= _zz_dataOut_payload_0_13815;
    _zz_dataOut_payload_0_15928 <= _zz_dataOut_payload_0_13816;
    _zz_dataOut_payload_0_15929 <= _zz_dataOut_payload_0_13817;
    _zz_dataOut_payload_0_15930 <= _zz_dataOut_payload_0_13818;
    _zz_dataOut_payload_0_15931 <= _zz_dataOut_payload_0_13819;
    _zz_dataOut_payload_0_15932 <= _zz_dataOut_payload_0_13820;
    _zz_dataOut_payload_0_15933 <= _zz_dataOut_payload_0_13821;
    _zz_dataOut_payload_0_15934 <= _zz_dataOut_payload_0_13822;
    _zz_dataOut_payload_0_15935 <= _zz_dataOut_payload_0_13823;
    _zz_dataOut_payload_0_15936 <= _zz_dataOut_payload_0_13824;
    _zz_dataOut_payload_0_15937 <= _zz_dataOut_payload_0_13825;
    _zz_dataOut_payload_0_15938 <= _zz_dataOut_payload_0_13826;
    _zz_dataOut_payload_0_15939 <= _zz_dataOut_payload_0_13827;
    _zz_dataOut_payload_0_15940 <= _zz_dataOut_payload_0_13828;
    _zz_dataOut_payload_0_15941 <= _zz_dataOut_payload_0_13829;
    _zz_dataOut_payload_0_15942 <= _zz_dataOut_payload_0_13830;
    _zz_dataOut_payload_0_15943 <= _zz_dataOut_payload_0_13831;
    _zz_dataOut_payload_0_15944 <= _zz_dataOut_payload_0_13832;
    _zz_dataOut_payload_0_15945 <= _zz_dataOut_payload_0_13833;
    _zz_dataOut_payload_0_15946 <= _zz_dataOut_payload_0_13834;
    _zz_dataOut_payload_0_15947 <= _zz_dataOut_payload_0_13835;
    _zz_dataOut_payload_0_15948 <= _zz_dataOut_payload_0_13836;
    _zz_dataOut_payload_0_15949 <= _zz_dataOut_payload_0_13837;
    _zz_dataOut_payload_0_15950 <= _zz_dataOut_payload_0_13838;
    _zz_dataOut_payload_0_15951 <= _zz_dataOut_payload_0_13839;
    _zz_dataOut_payload_0_15952 <= _zz_dataOut_payload_0_13840;
    _zz_dataOut_payload_0_15953 <= _zz_dataOut_payload_0_13841;
    _zz_dataOut_payload_0_15954 <= _zz_dataOut_payload_0_13842;
    _zz_dataOut_payload_0_15955 <= _zz_dataOut_payload_0_13843;
    _zz_dataOut_payload_0_15956 <= _zz_dataOut_payload_0_13844;
    _zz_dataOut_payload_0_15957 <= _zz_dataOut_payload_0_13845;
    _zz_dataOut_payload_0_15958 <= _zz_dataOut_payload_0_13846;
    _zz_dataOut_payload_0_15959 <= _zz_dataOut_payload_0_13847;
    _zz_dataOut_payload_0_15960 <= _zz_dataOut_payload_0_13848;
    _zz_dataOut_payload_0_15961 <= _zz_dataOut_payload_0_13849;
    _zz_dataOut_payload_0_15962 <= _zz_dataOut_payload_0_13850;
    _zz_dataOut_payload_0_15963 <= _zz_dataOut_payload_0_13851;
    _zz_dataOut_payload_0_15964 <= _zz_dataOut_payload_0_13852;
    _zz_dataOut_payload_0_15965 <= _zz_dataOut_payload_0_13853;
    _zz_dataOut_payload_0_15966 <= _zz_dataOut_payload_0_13854;
    _zz_dataOut_payload_0_15967 <= _zz_dataOut_payload_0_13855;
    _zz_dataOut_payload_0_15968 <= _zz_dataOut_payload_0_13856;
    _zz_dataOut_payload_0_15969 <= _zz_dataOut_payload_0_13857;
    _zz_dataOut_payload_0_15970 <= _zz_dataOut_payload_0_13858;
    _zz_dataOut_payload_0_15971 <= _zz_dataOut_payload_0_13859;
    _zz_dataOut_payload_0_15972 <= _zz_dataOut_payload_0_13860;
    _zz_dataOut_payload_0_15973 <= _zz_dataOut_payload_0_13861;
    _zz_dataOut_payload_0_15974 <= _zz_dataOut_payload_0_13862;
    _zz_dataOut_payload_0_15975 <= _zz_dataOut_payload_0_13863;
    _zz_dataOut_payload_0_15976 <= _zz_dataOut_payload_0_13864;
    _zz_dataOut_payload_0_15977 <= _zz_dataOut_payload_0_13865;
    _zz_dataOut_payload_0_15978 <= _zz_dataOut_payload_0_13866;
    _zz_dataOut_payload_0_15979 <= _zz_dataOut_payload_0_13867;
    _zz_dataOut_payload_0_15980 <= _zz_dataOut_payload_0_13868;
    _zz_dataOut_payload_0_15981 <= _zz_dataOut_payload_0_13869;
    _zz_dataOut_payload_0_15982 <= _zz_dataOut_payload_0_13870;
    _zz_dataOut_payload_0_15983 <= _zz_dataOut_payload_0_13871;
    _zz_dataOut_payload_0_15984 <= _zz_dataOut_payload_0_13872;
    _zz_dataOut_payload_0_15985 <= _zz_dataOut_payload_0_13873;
    _zz_dataOut_payload_0_15986 <= _zz_dataOut_payload_0_13874;
    _zz_dataOut_payload_0_15987 <= _zz_dataOut_payload_0_13875;
    _zz_dataOut_payload_0_15988 <= _zz_dataOut_payload_0_13876;
    _zz_dataOut_payload_0_15989 <= _zz_dataOut_payload_0_13877;
    _zz_dataOut_payload_0_15990 <= _zz_dataOut_payload_0_13878;
    _zz_dataOut_payload_0_15991 <= _zz_dataOut_payload_0_13879;
    _zz_dataOut_payload_0_15992 <= _zz_dataOut_payload_0_13880;
    _zz_dataOut_payload_0_15993 <= _zz_dataOut_payload_0_13881;
    _zz_dataOut_payload_0_15994 <= _zz_dataOut_payload_0_13882;
    _zz_dataOut_payload_0_15995 <= _zz_dataOut_payload_0_13883;
    _zz_dataOut_payload_0_15996 <= _zz_dataOut_payload_0_13884;
    _zz_dataOut_payload_0_15997 <= _zz_dataOut_payload_0_13885;
    _zz_dataOut_payload_0_15998 <= _zz_dataOut_payload_0_13886;
    _zz_dataOut_payload_0_15999 <= _zz_dataOut_payload_0_13887;
    _zz_dataOut_payload_0_16000 <= _zz_dataOut_payload_0_15744;
    _zz_dataOut_payload_0_16001 <= _zz_dataOut_payload_0_15745;
    _zz_dataOut_payload_0_16002 <= _zz_dataOut_payload_0_15746;
    _zz_dataOut_payload_0_16003 <= _zz_dataOut_payload_0_15747;
    _zz_dataOut_payload_0_16004 <= _zz_dataOut_payload_0_15748;
    _zz_dataOut_payload_0_16005 <= _zz_dataOut_payload_0_15749;
    _zz_dataOut_payload_0_16006 <= _zz_dataOut_payload_0_15750;
    _zz_dataOut_payload_0_16007 <= _zz_dataOut_payload_0_15751;
    _zz_dataOut_payload_0_16008 <= _zz_dataOut_payload_0_15752;
    _zz_dataOut_payload_0_16009 <= _zz_dataOut_payload_0_15753;
    _zz_dataOut_payload_0_16010 <= _zz_dataOut_payload_0_15754;
    _zz_dataOut_payload_0_16011 <= _zz_dataOut_payload_0_15755;
    _zz_dataOut_payload_0_16012 <= _zz_dataOut_payload_0_15756;
    _zz_dataOut_payload_0_16013 <= _zz_dataOut_payload_0_15757;
    _zz_dataOut_payload_0_16014 <= _zz_dataOut_payload_0_15758;
    _zz_dataOut_payload_0_16015 <= _zz_dataOut_payload_0_15759;
    _zz_dataOut_payload_0_16016 <= _zz_dataOut_payload_0_15760;
    _zz_dataOut_payload_0_16017 <= _zz_dataOut_payload_0_15761;
    _zz_dataOut_payload_0_16018 <= _zz_dataOut_payload_0_15762;
    _zz_dataOut_payload_0_16019 <= _zz_dataOut_payload_0_15763;
    _zz_dataOut_payload_0_16020 <= _zz_dataOut_payload_0_15764;
    _zz_dataOut_payload_0_16021 <= _zz_dataOut_payload_0_15765;
    _zz_dataOut_payload_0_16022 <= _zz_dataOut_payload_0_15766;
    _zz_dataOut_payload_0_16023 <= _zz_dataOut_payload_0_15767;
    _zz_dataOut_payload_0_16024 <= _zz_dataOut_payload_0_15768;
    _zz_dataOut_payload_0_16025 <= _zz_dataOut_payload_0_15769;
    _zz_dataOut_payload_0_16026 <= _zz_dataOut_payload_0_15770;
    _zz_dataOut_payload_0_16027 <= _zz_dataOut_payload_0_15771;
    _zz_dataOut_payload_0_16028 <= _zz_dataOut_payload_0_15772;
    _zz_dataOut_payload_0_16029 <= _zz_dataOut_payload_0_15773;
    _zz_dataOut_payload_0_16030 <= _zz_dataOut_payload_0_15774;
    _zz_dataOut_payload_0_16031 <= _zz_dataOut_payload_0_15775;
    _zz_dataOut_payload_0_16032 <= _zz_dataOut_payload_0_15776;
    _zz_dataOut_payload_0_16033 <= _zz_dataOut_payload_0_15777;
    _zz_dataOut_payload_0_16034 <= _zz_dataOut_payload_0_15778;
    _zz_dataOut_payload_0_16035 <= _zz_dataOut_payload_0_15779;
    _zz_dataOut_payload_0_16036 <= _zz_dataOut_payload_0_15780;
    _zz_dataOut_payload_0_16037 <= _zz_dataOut_payload_0_15781;
    _zz_dataOut_payload_0_16038 <= _zz_dataOut_payload_0_15782;
    _zz_dataOut_payload_0_16039 <= _zz_dataOut_payload_0_15783;
    _zz_dataOut_payload_0_16040 <= _zz_dataOut_payload_0_15784;
    _zz_dataOut_payload_0_16041 <= _zz_dataOut_payload_0_15785;
    _zz_dataOut_payload_0_16042 <= _zz_dataOut_payload_0_15786;
    _zz_dataOut_payload_0_16043 <= _zz_dataOut_payload_0_15787;
    _zz_dataOut_payload_0_16044 <= _zz_dataOut_payload_0_15788;
    _zz_dataOut_payload_0_16045 <= _zz_dataOut_payload_0_15789;
    _zz_dataOut_payload_0_16046 <= _zz_dataOut_payload_0_15790;
    _zz_dataOut_payload_0_16047 <= _zz_dataOut_payload_0_15791;
    _zz_dataOut_payload_0_16048 <= _zz_dataOut_payload_0_15792;
    _zz_dataOut_payload_0_16049 <= _zz_dataOut_payload_0_15793;
    _zz_dataOut_payload_0_16050 <= _zz_dataOut_payload_0_15794;
    _zz_dataOut_payload_0_16051 <= _zz_dataOut_payload_0_15795;
    _zz_dataOut_payload_0_16052 <= _zz_dataOut_payload_0_15796;
    _zz_dataOut_payload_0_16053 <= _zz_dataOut_payload_0_15797;
    _zz_dataOut_payload_0_16054 <= _zz_dataOut_payload_0_15798;
    _zz_dataOut_payload_0_16055 <= _zz_dataOut_payload_0_15799;
    _zz_dataOut_payload_0_16056 <= _zz_dataOut_payload_0_15800;
    _zz_dataOut_payload_0_16057 <= _zz_dataOut_payload_0_15801;
    _zz_dataOut_payload_0_16058 <= _zz_dataOut_payload_0_15802;
    _zz_dataOut_payload_0_16059 <= _zz_dataOut_payload_0_15803;
    _zz_dataOut_payload_0_16060 <= _zz_dataOut_payload_0_15804;
    _zz_dataOut_payload_0_16061 <= _zz_dataOut_payload_0_15805;
    _zz_dataOut_payload_0_16062 <= _zz_dataOut_payload_0_15806;
    _zz_dataOut_payload_0_16063 <= _zz_dataOut_payload_0_15807;
    _zz_dataOut_payload_0_16064 <= _zz_dataOut_payload_0_15808;
    _zz_dataOut_payload_0_16065 <= _zz_dataOut_payload_0_15809;
    _zz_dataOut_payload_0_16066 <= _zz_dataOut_payload_0_15810;
    _zz_dataOut_payload_0_16067 <= _zz_dataOut_payload_0_15811;
    _zz_dataOut_payload_0_16068 <= _zz_dataOut_payload_0_15812;
    _zz_dataOut_payload_0_16069 <= _zz_dataOut_payload_0_15813;
    _zz_dataOut_payload_0_16070 <= _zz_dataOut_payload_0_15814;
    _zz_dataOut_payload_0_16071 <= _zz_dataOut_payload_0_15815;
    _zz_dataOut_payload_0_16072 <= _zz_dataOut_payload_0_15816;
    _zz_dataOut_payload_0_16073 <= _zz_dataOut_payload_0_15817;
    _zz_dataOut_payload_0_16074 <= _zz_dataOut_payload_0_15818;
    _zz_dataOut_payload_0_16075 <= _zz_dataOut_payload_0_15819;
    _zz_dataOut_payload_0_16076 <= _zz_dataOut_payload_0_15820;
    _zz_dataOut_payload_0_16077 <= _zz_dataOut_payload_0_15821;
    _zz_dataOut_payload_0_16078 <= _zz_dataOut_payload_0_15822;
    _zz_dataOut_payload_0_16079 <= _zz_dataOut_payload_0_15823;
    _zz_dataOut_payload_0_16080 <= _zz_dataOut_payload_0_15824;
    _zz_dataOut_payload_0_16081 <= _zz_dataOut_payload_0_15825;
    _zz_dataOut_payload_0_16082 <= _zz_dataOut_payload_0_15826;
    _zz_dataOut_payload_0_16083 <= _zz_dataOut_payload_0_15827;
    _zz_dataOut_payload_0_16084 <= _zz_dataOut_payload_0_15828;
    _zz_dataOut_payload_0_16085 <= _zz_dataOut_payload_0_15829;
    _zz_dataOut_payload_0_16086 <= _zz_dataOut_payload_0_15830;
    _zz_dataOut_payload_0_16087 <= _zz_dataOut_payload_0_15831;
    _zz_dataOut_payload_0_16088 <= _zz_dataOut_payload_0_15832;
    _zz_dataOut_payload_0_16089 <= _zz_dataOut_payload_0_15833;
    _zz_dataOut_payload_0_16090 <= _zz_dataOut_payload_0_15834;
    _zz_dataOut_payload_0_16091 <= _zz_dataOut_payload_0_15835;
    _zz_dataOut_payload_0_16092 <= _zz_dataOut_payload_0_15836;
    _zz_dataOut_payload_0_16093 <= _zz_dataOut_payload_0_15837;
    _zz_dataOut_payload_0_16094 <= _zz_dataOut_payload_0_15838;
    _zz_dataOut_payload_0_16095 <= _zz_dataOut_payload_0_15839;
    _zz_dataOut_payload_0_16096 <= _zz_dataOut_payload_0_15840;
    _zz_dataOut_payload_0_16097 <= _zz_dataOut_payload_0_15841;
    _zz_dataOut_payload_0_16098 <= _zz_dataOut_payload_0_15842;
    _zz_dataOut_payload_0_16099 <= _zz_dataOut_payload_0_15843;
    _zz_dataOut_payload_0_16100 <= _zz_dataOut_payload_0_15844;
    _zz_dataOut_payload_0_16101 <= _zz_dataOut_payload_0_15845;
    _zz_dataOut_payload_0_16102 <= _zz_dataOut_payload_0_15846;
    _zz_dataOut_payload_0_16103 <= _zz_dataOut_payload_0_15847;
    _zz_dataOut_payload_0_16104 <= _zz_dataOut_payload_0_15848;
    _zz_dataOut_payload_0_16105 <= _zz_dataOut_payload_0_15849;
    _zz_dataOut_payload_0_16106 <= _zz_dataOut_payload_0_15850;
    _zz_dataOut_payload_0_16107 <= _zz_dataOut_payload_0_15851;
    _zz_dataOut_payload_0_16108 <= _zz_dataOut_payload_0_15852;
    _zz_dataOut_payload_0_16109 <= _zz_dataOut_payload_0_15853;
    _zz_dataOut_payload_0_16110 <= _zz_dataOut_payload_0_15854;
    _zz_dataOut_payload_0_16111 <= _zz_dataOut_payload_0_15855;
    _zz_dataOut_payload_0_16112 <= _zz_dataOut_payload_0_15856;
    _zz_dataOut_payload_0_16113 <= _zz_dataOut_payload_0_15857;
    _zz_dataOut_payload_0_16114 <= _zz_dataOut_payload_0_15858;
    _zz_dataOut_payload_0_16115 <= _zz_dataOut_payload_0_15859;
    _zz_dataOut_payload_0_16116 <= _zz_dataOut_payload_0_15860;
    _zz_dataOut_payload_0_16117 <= _zz_dataOut_payload_0_15861;
    _zz_dataOut_payload_0_16118 <= _zz_dataOut_payload_0_15862;
    _zz_dataOut_payload_0_16119 <= _zz_dataOut_payload_0_15863;
    _zz_dataOut_payload_0_16120 <= _zz_dataOut_payload_0_15864;
    _zz_dataOut_payload_0_16121 <= _zz_dataOut_payload_0_15865;
    _zz_dataOut_payload_0_16122 <= _zz_dataOut_payload_0_15866;
    _zz_dataOut_payload_0_16123 <= _zz_dataOut_payload_0_15867;
    _zz_dataOut_payload_0_16124 <= _zz_dataOut_payload_0_15868;
    _zz_dataOut_payload_0_16125 <= _zz_dataOut_payload_0_15869;
    _zz_dataOut_payload_0_16126 <= _zz_dataOut_payload_0_15870;
    _zz_dataOut_payload_0_16127 <= _zz_dataOut_payload_0_15871;
    _zz_dataOut_payload_0_16637 <= (_zz_dataOut_payload_0_16636 ? _zz_dataOut_payload_0_16633 : _zz_dataOut_payload_0_16635);
    _zz_dataOut_payload_1 <= (_zz_dataOut_payload_0_16636 ? _zz_dataOut_payload_0_16635 : _zz_dataOut_payload_0_16633);
    _zz_dataOut_payload_2_3 <= (_zz_dataOut_payload_2_2 ? _zz_dataOut_payload_2 : _zz_dataOut_payload_2_1);
    _zz_dataOut_payload_3 <= (_zz_dataOut_payload_2_2 ? _zz_dataOut_payload_2_1 : _zz_dataOut_payload_2);
    _zz_dataOut_payload_4_9 <= (_zz_dataOut_payload_4_8 ? _zz_dataOut_payload_4_5 : _zz_dataOut_payload_4_7);
    _zz_dataOut_payload_5 <= (_zz_dataOut_payload_4_8 ? _zz_dataOut_payload_4_7 : _zz_dataOut_payload_4_5);
    _zz_dataOut_payload_6_3 <= (_zz_dataOut_payload_6_2 ? _zz_dataOut_payload_6 : _zz_dataOut_payload_6_1);
    _zz_dataOut_payload_7 <= (_zz_dataOut_payload_6_2 ? _zz_dataOut_payload_6_1 : _zz_dataOut_payload_6);
    _zz_dataOut_payload_0_16638 <= _zz_dataOut_payload_0_16637;
    _zz_dataOut_payload_1_1 <= _zz_dataOut_payload_1;
    _zz_dataOut_payload_2_4 <= _zz_dataOut_payload_2_3;
    _zz_dataOut_payload_3_1 <= _zz_dataOut_payload_3;
    _zz_dataOut_payload_4_10 <= _zz_dataOut_payload_4_9;
    _zz_dataOut_payload_5_1 <= _zz_dataOut_payload_5;
    _zz_dataOut_payload_6_4 <= _zz_dataOut_payload_6_3;
    _zz_dataOut_payload_7_1 <= _zz_dataOut_payload_7;
    _zz_dataOut_payload_8_21 <= (_zz_dataOut_payload_8_20 ? _zz_dataOut_payload_8_17 : _zz_dataOut_payload_8_19);
    _zz_dataOut_payload_9 <= (_zz_dataOut_payload_8_20 ? _zz_dataOut_payload_8_19 : _zz_dataOut_payload_8_17);
    _zz_dataOut_payload_10_3 <= (_zz_dataOut_payload_10_2 ? _zz_dataOut_payload_10 : _zz_dataOut_payload_10_1);
    _zz_dataOut_payload_11 <= (_zz_dataOut_payload_10_2 ? _zz_dataOut_payload_10_1 : _zz_dataOut_payload_10);
    _zz_dataOut_payload_12_9 <= (_zz_dataOut_payload_12_8 ? _zz_dataOut_payload_12_5 : _zz_dataOut_payload_12_7);
    _zz_dataOut_payload_13 <= (_zz_dataOut_payload_12_8 ? _zz_dataOut_payload_12_7 : _zz_dataOut_payload_12_5);
    _zz_dataOut_payload_14_3 <= (_zz_dataOut_payload_14_2 ? _zz_dataOut_payload_14 : _zz_dataOut_payload_14_1);
    _zz_dataOut_payload_15 <= (_zz_dataOut_payload_14_2 ? _zz_dataOut_payload_14_1 : _zz_dataOut_payload_14);
    _zz_dataOut_payload_8_22 <= _zz_dataOut_payload_8_21;
    _zz_dataOut_payload_9_1 <= _zz_dataOut_payload_9;
    _zz_dataOut_payload_10_4 <= _zz_dataOut_payload_10_3;
    _zz_dataOut_payload_11_1 <= _zz_dataOut_payload_11;
    _zz_dataOut_payload_12_10 <= _zz_dataOut_payload_12_9;
    _zz_dataOut_payload_13_1 <= _zz_dataOut_payload_13;
    _zz_dataOut_payload_14_4 <= _zz_dataOut_payload_14_3;
    _zz_dataOut_payload_15_1 <= _zz_dataOut_payload_15;
    _zz_dataOut_payload_0_16639 <= _zz_dataOut_payload_0_16638;
    _zz_dataOut_payload_1_2 <= _zz_dataOut_payload_1_1;
    _zz_dataOut_payload_2_5 <= _zz_dataOut_payload_2_4;
    _zz_dataOut_payload_3_2 <= _zz_dataOut_payload_3_1;
    _zz_dataOut_payload_4_11 <= _zz_dataOut_payload_4_10;
    _zz_dataOut_payload_5_2 <= _zz_dataOut_payload_5_1;
    _zz_dataOut_payload_6_5 <= _zz_dataOut_payload_6_4;
    _zz_dataOut_payload_7_2 <= _zz_dataOut_payload_7_1;
    _zz_dataOut_payload_8_23 <= _zz_dataOut_payload_8_22;
    _zz_dataOut_payload_9_2 <= _zz_dataOut_payload_9_1;
    _zz_dataOut_payload_10_5 <= _zz_dataOut_payload_10_4;
    _zz_dataOut_payload_11_2 <= _zz_dataOut_payload_11_1;
    _zz_dataOut_payload_12_11 <= _zz_dataOut_payload_12_10;
    _zz_dataOut_payload_13_2 <= _zz_dataOut_payload_13_1;
    _zz_dataOut_payload_14_5 <= _zz_dataOut_payload_14_4;
    _zz_dataOut_payload_15_2 <= _zz_dataOut_payload_15_1;
    _zz_dataOut_payload_16_45 <= (_zz_dataOut_payload_16_44 ? _zz_dataOut_payload_16_41 : _zz_dataOut_payload_16_43);
    _zz_dataOut_payload_17 <= (_zz_dataOut_payload_16_44 ? _zz_dataOut_payload_16_43 : _zz_dataOut_payload_16_41);
    _zz_dataOut_payload_18_3 <= (_zz_dataOut_payload_18_2 ? _zz_dataOut_payload_18 : _zz_dataOut_payload_18_1);
    _zz_dataOut_payload_19 <= (_zz_dataOut_payload_18_2 ? _zz_dataOut_payload_18_1 : _zz_dataOut_payload_18);
    _zz_dataOut_payload_20_9 <= (_zz_dataOut_payload_20_8 ? _zz_dataOut_payload_20_5 : _zz_dataOut_payload_20_7);
    _zz_dataOut_payload_21 <= (_zz_dataOut_payload_20_8 ? _zz_dataOut_payload_20_7 : _zz_dataOut_payload_20_5);
    _zz_dataOut_payload_22_3 <= (_zz_dataOut_payload_22_2 ? _zz_dataOut_payload_22 : _zz_dataOut_payload_22_1);
    _zz_dataOut_payload_23 <= (_zz_dataOut_payload_22_2 ? _zz_dataOut_payload_22_1 : _zz_dataOut_payload_22);
    _zz_dataOut_payload_16_46 <= _zz_dataOut_payload_16_45;
    _zz_dataOut_payload_17_1 <= _zz_dataOut_payload_17;
    _zz_dataOut_payload_18_4 <= _zz_dataOut_payload_18_3;
    _zz_dataOut_payload_19_1 <= _zz_dataOut_payload_19;
    _zz_dataOut_payload_20_10 <= _zz_dataOut_payload_20_9;
    _zz_dataOut_payload_21_1 <= _zz_dataOut_payload_21;
    _zz_dataOut_payload_22_4 <= _zz_dataOut_payload_22_3;
    _zz_dataOut_payload_23_1 <= _zz_dataOut_payload_23;
    _zz_dataOut_payload_24_21 <= (_zz_dataOut_payload_24_20 ? _zz_dataOut_payload_24_17 : _zz_dataOut_payload_24_19);
    _zz_dataOut_payload_25 <= (_zz_dataOut_payload_24_20 ? _zz_dataOut_payload_24_19 : _zz_dataOut_payload_24_17);
    _zz_dataOut_payload_26_3 <= (_zz_dataOut_payload_26_2 ? _zz_dataOut_payload_26 : _zz_dataOut_payload_26_1);
    _zz_dataOut_payload_27 <= (_zz_dataOut_payload_26_2 ? _zz_dataOut_payload_26_1 : _zz_dataOut_payload_26);
    _zz_dataOut_payload_28_9 <= (_zz_dataOut_payload_28_8 ? _zz_dataOut_payload_28_5 : _zz_dataOut_payload_28_7);
    _zz_dataOut_payload_29 <= (_zz_dataOut_payload_28_8 ? _zz_dataOut_payload_28_7 : _zz_dataOut_payload_28_5);
    _zz_dataOut_payload_30_3 <= (_zz_dataOut_payload_30_2 ? _zz_dataOut_payload_30 : _zz_dataOut_payload_30_1);
    _zz_dataOut_payload_31 <= (_zz_dataOut_payload_30_2 ? _zz_dataOut_payload_30_1 : _zz_dataOut_payload_30);
    _zz_dataOut_payload_24_22 <= _zz_dataOut_payload_24_21;
    _zz_dataOut_payload_25_1 <= _zz_dataOut_payload_25;
    _zz_dataOut_payload_26_4 <= _zz_dataOut_payload_26_3;
    _zz_dataOut_payload_27_1 <= _zz_dataOut_payload_27;
    _zz_dataOut_payload_28_10 <= _zz_dataOut_payload_28_9;
    _zz_dataOut_payload_29_1 <= _zz_dataOut_payload_29;
    _zz_dataOut_payload_30_4 <= _zz_dataOut_payload_30_3;
    _zz_dataOut_payload_31_1 <= _zz_dataOut_payload_31;
    _zz_dataOut_payload_16_47 <= _zz_dataOut_payload_16_46;
    _zz_dataOut_payload_17_2 <= _zz_dataOut_payload_17_1;
    _zz_dataOut_payload_18_5 <= _zz_dataOut_payload_18_4;
    _zz_dataOut_payload_19_2 <= _zz_dataOut_payload_19_1;
    _zz_dataOut_payload_20_11 <= _zz_dataOut_payload_20_10;
    _zz_dataOut_payload_21_2 <= _zz_dataOut_payload_21_1;
    _zz_dataOut_payload_22_5 <= _zz_dataOut_payload_22_4;
    _zz_dataOut_payload_23_2 <= _zz_dataOut_payload_23_1;
    _zz_dataOut_payload_24_23 <= _zz_dataOut_payload_24_22;
    _zz_dataOut_payload_25_2 <= _zz_dataOut_payload_25_1;
    _zz_dataOut_payload_26_5 <= _zz_dataOut_payload_26_4;
    _zz_dataOut_payload_27_2 <= _zz_dataOut_payload_27_1;
    _zz_dataOut_payload_28_11 <= _zz_dataOut_payload_28_10;
    _zz_dataOut_payload_29_2 <= _zz_dataOut_payload_29_1;
    _zz_dataOut_payload_30_5 <= _zz_dataOut_payload_30_4;
    _zz_dataOut_payload_31_2 <= _zz_dataOut_payload_31_1;
    _zz_dataOut_payload_0_16640 <= _zz_dataOut_payload_0_16639;
    _zz_dataOut_payload_1_3 <= _zz_dataOut_payload_1_2;
    _zz_dataOut_payload_2_6 <= _zz_dataOut_payload_2_5;
    _zz_dataOut_payload_3_3 <= _zz_dataOut_payload_3_2;
    _zz_dataOut_payload_4_12 <= _zz_dataOut_payload_4_11;
    _zz_dataOut_payload_5_3 <= _zz_dataOut_payload_5_2;
    _zz_dataOut_payload_6_6 <= _zz_dataOut_payload_6_5;
    _zz_dataOut_payload_7_3 <= _zz_dataOut_payload_7_2;
    _zz_dataOut_payload_8_24 <= _zz_dataOut_payload_8_23;
    _zz_dataOut_payload_9_3 <= _zz_dataOut_payload_9_2;
    _zz_dataOut_payload_10_6 <= _zz_dataOut_payload_10_5;
    _zz_dataOut_payload_11_3 <= _zz_dataOut_payload_11_2;
    _zz_dataOut_payload_12_12 <= _zz_dataOut_payload_12_11;
    _zz_dataOut_payload_13_3 <= _zz_dataOut_payload_13_2;
    _zz_dataOut_payload_14_6 <= _zz_dataOut_payload_14_5;
    _zz_dataOut_payload_15_3 <= _zz_dataOut_payload_15_2;
    _zz_dataOut_payload_16_48 <= _zz_dataOut_payload_16_47;
    _zz_dataOut_payload_17_3 <= _zz_dataOut_payload_17_2;
    _zz_dataOut_payload_18_6 <= _zz_dataOut_payload_18_5;
    _zz_dataOut_payload_19_3 <= _zz_dataOut_payload_19_2;
    _zz_dataOut_payload_20_12 <= _zz_dataOut_payload_20_11;
    _zz_dataOut_payload_21_3 <= _zz_dataOut_payload_21_2;
    _zz_dataOut_payload_22_6 <= _zz_dataOut_payload_22_5;
    _zz_dataOut_payload_23_3 <= _zz_dataOut_payload_23_2;
    _zz_dataOut_payload_24_24 <= _zz_dataOut_payload_24_23;
    _zz_dataOut_payload_25_3 <= _zz_dataOut_payload_25_2;
    _zz_dataOut_payload_26_6 <= _zz_dataOut_payload_26_5;
    _zz_dataOut_payload_27_3 <= _zz_dataOut_payload_27_2;
    _zz_dataOut_payload_28_12 <= _zz_dataOut_payload_28_11;
    _zz_dataOut_payload_29_3 <= _zz_dataOut_payload_29_2;
    _zz_dataOut_payload_30_6 <= _zz_dataOut_payload_30_5;
    _zz_dataOut_payload_31_3 <= _zz_dataOut_payload_31_2;
    _zz_dataOut_payload_32_93 <= (_zz_dataOut_payload_32_92 ? _zz_dataOut_payload_32_89 : _zz_dataOut_payload_32_91);
    _zz_dataOut_payload_33 <= (_zz_dataOut_payload_32_92 ? _zz_dataOut_payload_32_91 : _zz_dataOut_payload_32_89);
    _zz_dataOut_payload_34_3 <= (_zz_dataOut_payload_34_2 ? _zz_dataOut_payload_34 : _zz_dataOut_payload_34_1);
    _zz_dataOut_payload_35 <= (_zz_dataOut_payload_34_2 ? _zz_dataOut_payload_34_1 : _zz_dataOut_payload_34);
    _zz_dataOut_payload_36_9 <= (_zz_dataOut_payload_36_8 ? _zz_dataOut_payload_36_5 : _zz_dataOut_payload_36_7);
    _zz_dataOut_payload_37 <= (_zz_dataOut_payload_36_8 ? _zz_dataOut_payload_36_7 : _zz_dataOut_payload_36_5);
    _zz_dataOut_payload_38_3 <= (_zz_dataOut_payload_38_2 ? _zz_dataOut_payload_38 : _zz_dataOut_payload_38_1);
    _zz_dataOut_payload_39 <= (_zz_dataOut_payload_38_2 ? _zz_dataOut_payload_38_1 : _zz_dataOut_payload_38);
    _zz_dataOut_payload_32_94 <= _zz_dataOut_payload_32_93;
    _zz_dataOut_payload_33_1 <= _zz_dataOut_payload_33;
    _zz_dataOut_payload_34_4 <= _zz_dataOut_payload_34_3;
    _zz_dataOut_payload_35_1 <= _zz_dataOut_payload_35;
    _zz_dataOut_payload_36_10 <= _zz_dataOut_payload_36_9;
    _zz_dataOut_payload_37_1 <= _zz_dataOut_payload_37;
    _zz_dataOut_payload_38_4 <= _zz_dataOut_payload_38_3;
    _zz_dataOut_payload_39_1 <= _zz_dataOut_payload_39;
    _zz_dataOut_payload_40_21 <= (_zz_dataOut_payload_40_20 ? _zz_dataOut_payload_40_17 : _zz_dataOut_payload_40_19);
    _zz_dataOut_payload_41 <= (_zz_dataOut_payload_40_20 ? _zz_dataOut_payload_40_19 : _zz_dataOut_payload_40_17);
    _zz_dataOut_payload_42_3 <= (_zz_dataOut_payload_42_2 ? _zz_dataOut_payload_42 : _zz_dataOut_payload_42_1);
    _zz_dataOut_payload_43 <= (_zz_dataOut_payload_42_2 ? _zz_dataOut_payload_42_1 : _zz_dataOut_payload_42);
    _zz_dataOut_payload_44_9 <= (_zz_dataOut_payload_44_8 ? _zz_dataOut_payload_44_5 : _zz_dataOut_payload_44_7);
    _zz_dataOut_payload_45 <= (_zz_dataOut_payload_44_8 ? _zz_dataOut_payload_44_7 : _zz_dataOut_payload_44_5);
    _zz_dataOut_payload_46_3 <= (_zz_dataOut_payload_46_2 ? _zz_dataOut_payload_46 : _zz_dataOut_payload_46_1);
    _zz_dataOut_payload_47 <= (_zz_dataOut_payload_46_2 ? _zz_dataOut_payload_46_1 : _zz_dataOut_payload_46);
    _zz_dataOut_payload_40_22 <= _zz_dataOut_payload_40_21;
    _zz_dataOut_payload_41_1 <= _zz_dataOut_payload_41;
    _zz_dataOut_payload_42_4 <= _zz_dataOut_payload_42_3;
    _zz_dataOut_payload_43_1 <= _zz_dataOut_payload_43;
    _zz_dataOut_payload_44_10 <= _zz_dataOut_payload_44_9;
    _zz_dataOut_payload_45_1 <= _zz_dataOut_payload_45;
    _zz_dataOut_payload_46_4 <= _zz_dataOut_payload_46_3;
    _zz_dataOut_payload_47_1 <= _zz_dataOut_payload_47;
    _zz_dataOut_payload_32_95 <= _zz_dataOut_payload_32_94;
    _zz_dataOut_payload_33_2 <= _zz_dataOut_payload_33_1;
    _zz_dataOut_payload_34_5 <= _zz_dataOut_payload_34_4;
    _zz_dataOut_payload_35_2 <= _zz_dataOut_payload_35_1;
    _zz_dataOut_payload_36_11 <= _zz_dataOut_payload_36_10;
    _zz_dataOut_payload_37_2 <= _zz_dataOut_payload_37_1;
    _zz_dataOut_payload_38_5 <= _zz_dataOut_payload_38_4;
    _zz_dataOut_payload_39_2 <= _zz_dataOut_payload_39_1;
    _zz_dataOut_payload_40_23 <= _zz_dataOut_payload_40_22;
    _zz_dataOut_payload_41_2 <= _zz_dataOut_payload_41_1;
    _zz_dataOut_payload_42_5 <= _zz_dataOut_payload_42_4;
    _zz_dataOut_payload_43_2 <= _zz_dataOut_payload_43_1;
    _zz_dataOut_payload_44_11 <= _zz_dataOut_payload_44_10;
    _zz_dataOut_payload_45_2 <= _zz_dataOut_payload_45_1;
    _zz_dataOut_payload_46_5 <= _zz_dataOut_payload_46_4;
    _zz_dataOut_payload_47_2 <= _zz_dataOut_payload_47_1;
    _zz_dataOut_payload_48_45 <= (_zz_dataOut_payload_48_44 ? _zz_dataOut_payload_48_41 : _zz_dataOut_payload_48_43);
    _zz_dataOut_payload_49 <= (_zz_dataOut_payload_48_44 ? _zz_dataOut_payload_48_43 : _zz_dataOut_payload_48_41);
    _zz_dataOut_payload_50_3 <= (_zz_dataOut_payload_50_2 ? _zz_dataOut_payload_50 : _zz_dataOut_payload_50_1);
    _zz_dataOut_payload_51 <= (_zz_dataOut_payload_50_2 ? _zz_dataOut_payload_50_1 : _zz_dataOut_payload_50);
    _zz_dataOut_payload_52_9 <= (_zz_dataOut_payload_52_8 ? _zz_dataOut_payload_52_5 : _zz_dataOut_payload_52_7);
    _zz_dataOut_payload_53 <= (_zz_dataOut_payload_52_8 ? _zz_dataOut_payload_52_7 : _zz_dataOut_payload_52_5);
    _zz_dataOut_payload_54_3 <= (_zz_dataOut_payload_54_2 ? _zz_dataOut_payload_54 : _zz_dataOut_payload_54_1);
    _zz_dataOut_payload_55 <= (_zz_dataOut_payload_54_2 ? _zz_dataOut_payload_54_1 : _zz_dataOut_payload_54);
    _zz_dataOut_payload_48_46 <= _zz_dataOut_payload_48_45;
    _zz_dataOut_payload_49_1 <= _zz_dataOut_payload_49;
    _zz_dataOut_payload_50_4 <= _zz_dataOut_payload_50_3;
    _zz_dataOut_payload_51_1 <= _zz_dataOut_payload_51;
    _zz_dataOut_payload_52_10 <= _zz_dataOut_payload_52_9;
    _zz_dataOut_payload_53_1 <= _zz_dataOut_payload_53;
    _zz_dataOut_payload_54_4 <= _zz_dataOut_payload_54_3;
    _zz_dataOut_payload_55_1 <= _zz_dataOut_payload_55;
    _zz_dataOut_payload_56_21 <= (_zz_dataOut_payload_56_20 ? _zz_dataOut_payload_56_17 : _zz_dataOut_payload_56_19);
    _zz_dataOut_payload_57 <= (_zz_dataOut_payload_56_20 ? _zz_dataOut_payload_56_19 : _zz_dataOut_payload_56_17);
    _zz_dataOut_payload_58_3 <= (_zz_dataOut_payload_58_2 ? _zz_dataOut_payload_58 : _zz_dataOut_payload_58_1);
    _zz_dataOut_payload_59 <= (_zz_dataOut_payload_58_2 ? _zz_dataOut_payload_58_1 : _zz_dataOut_payload_58);
    _zz_dataOut_payload_60_9 <= (_zz_dataOut_payload_60_8 ? _zz_dataOut_payload_60_5 : _zz_dataOut_payload_60_7);
    _zz_dataOut_payload_61 <= (_zz_dataOut_payload_60_8 ? _zz_dataOut_payload_60_7 : _zz_dataOut_payload_60_5);
    _zz_dataOut_payload_62_3 <= (_zz_dataOut_payload_62_2 ? _zz_dataOut_payload_62 : _zz_dataOut_payload_62_1);
    _zz_dataOut_payload_63 <= (_zz_dataOut_payload_62_2 ? _zz_dataOut_payload_62_1 : _zz_dataOut_payload_62);
    _zz_dataOut_payload_56_22 <= _zz_dataOut_payload_56_21;
    _zz_dataOut_payload_57_1 <= _zz_dataOut_payload_57;
    _zz_dataOut_payload_58_4 <= _zz_dataOut_payload_58_3;
    _zz_dataOut_payload_59_1 <= _zz_dataOut_payload_59;
    _zz_dataOut_payload_60_10 <= _zz_dataOut_payload_60_9;
    _zz_dataOut_payload_61_1 <= _zz_dataOut_payload_61;
    _zz_dataOut_payload_62_4 <= _zz_dataOut_payload_62_3;
    _zz_dataOut_payload_63_1 <= _zz_dataOut_payload_63;
    _zz_dataOut_payload_48_47 <= _zz_dataOut_payload_48_46;
    _zz_dataOut_payload_49_2 <= _zz_dataOut_payload_49_1;
    _zz_dataOut_payload_50_5 <= _zz_dataOut_payload_50_4;
    _zz_dataOut_payload_51_2 <= _zz_dataOut_payload_51_1;
    _zz_dataOut_payload_52_11 <= _zz_dataOut_payload_52_10;
    _zz_dataOut_payload_53_2 <= _zz_dataOut_payload_53_1;
    _zz_dataOut_payload_54_5 <= _zz_dataOut_payload_54_4;
    _zz_dataOut_payload_55_2 <= _zz_dataOut_payload_55_1;
    _zz_dataOut_payload_56_23 <= _zz_dataOut_payload_56_22;
    _zz_dataOut_payload_57_2 <= _zz_dataOut_payload_57_1;
    _zz_dataOut_payload_58_5 <= _zz_dataOut_payload_58_4;
    _zz_dataOut_payload_59_2 <= _zz_dataOut_payload_59_1;
    _zz_dataOut_payload_60_11 <= _zz_dataOut_payload_60_10;
    _zz_dataOut_payload_61_2 <= _zz_dataOut_payload_61_1;
    _zz_dataOut_payload_62_5 <= _zz_dataOut_payload_62_4;
    _zz_dataOut_payload_63_2 <= _zz_dataOut_payload_63_1;
    _zz_dataOut_payload_32_96 <= _zz_dataOut_payload_32_95;
    _zz_dataOut_payload_33_3 <= _zz_dataOut_payload_33_2;
    _zz_dataOut_payload_34_6 <= _zz_dataOut_payload_34_5;
    _zz_dataOut_payload_35_3 <= _zz_dataOut_payload_35_2;
    _zz_dataOut_payload_36_12 <= _zz_dataOut_payload_36_11;
    _zz_dataOut_payload_37_3 <= _zz_dataOut_payload_37_2;
    _zz_dataOut_payload_38_6 <= _zz_dataOut_payload_38_5;
    _zz_dataOut_payload_39_3 <= _zz_dataOut_payload_39_2;
    _zz_dataOut_payload_40_24 <= _zz_dataOut_payload_40_23;
    _zz_dataOut_payload_41_3 <= _zz_dataOut_payload_41_2;
    _zz_dataOut_payload_42_6 <= _zz_dataOut_payload_42_5;
    _zz_dataOut_payload_43_3 <= _zz_dataOut_payload_43_2;
    _zz_dataOut_payload_44_12 <= _zz_dataOut_payload_44_11;
    _zz_dataOut_payload_45_3 <= _zz_dataOut_payload_45_2;
    _zz_dataOut_payload_46_6 <= _zz_dataOut_payload_46_5;
    _zz_dataOut_payload_47_3 <= _zz_dataOut_payload_47_2;
    _zz_dataOut_payload_48_48 <= _zz_dataOut_payload_48_47;
    _zz_dataOut_payload_49_3 <= _zz_dataOut_payload_49_2;
    _zz_dataOut_payload_50_6 <= _zz_dataOut_payload_50_5;
    _zz_dataOut_payload_51_3 <= _zz_dataOut_payload_51_2;
    _zz_dataOut_payload_52_12 <= _zz_dataOut_payload_52_11;
    _zz_dataOut_payload_53_3 <= _zz_dataOut_payload_53_2;
    _zz_dataOut_payload_54_6 <= _zz_dataOut_payload_54_5;
    _zz_dataOut_payload_55_3 <= _zz_dataOut_payload_55_2;
    _zz_dataOut_payload_56_24 <= _zz_dataOut_payload_56_23;
    _zz_dataOut_payload_57_3 <= _zz_dataOut_payload_57_2;
    _zz_dataOut_payload_58_6 <= _zz_dataOut_payload_58_5;
    _zz_dataOut_payload_59_3 <= _zz_dataOut_payload_59_2;
    _zz_dataOut_payload_60_12 <= _zz_dataOut_payload_60_11;
    _zz_dataOut_payload_61_3 <= _zz_dataOut_payload_61_2;
    _zz_dataOut_payload_62_6 <= _zz_dataOut_payload_62_5;
    _zz_dataOut_payload_63_3 <= _zz_dataOut_payload_63_2;
    _zz_dataOut_payload_0_16641 <= _zz_dataOut_payload_0_16640;
    _zz_dataOut_payload_1_4 <= _zz_dataOut_payload_1_3;
    _zz_dataOut_payload_2_7 <= _zz_dataOut_payload_2_6;
    _zz_dataOut_payload_3_4 <= _zz_dataOut_payload_3_3;
    _zz_dataOut_payload_4_13 <= _zz_dataOut_payload_4_12;
    _zz_dataOut_payload_5_4 <= _zz_dataOut_payload_5_3;
    _zz_dataOut_payload_6_7 <= _zz_dataOut_payload_6_6;
    _zz_dataOut_payload_7_4 <= _zz_dataOut_payload_7_3;
    _zz_dataOut_payload_8_25 <= _zz_dataOut_payload_8_24;
    _zz_dataOut_payload_9_4 <= _zz_dataOut_payload_9_3;
    _zz_dataOut_payload_10_7 <= _zz_dataOut_payload_10_6;
    _zz_dataOut_payload_11_4 <= _zz_dataOut_payload_11_3;
    _zz_dataOut_payload_12_13 <= _zz_dataOut_payload_12_12;
    _zz_dataOut_payload_13_4 <= _zz_dataOut_payload_13_3;
    _zz_dataOut_payload_14_7 <= _zz_dataOut_payload_14_6;
    _zz_dataOut_payload_15_4 <= _zz_dataOut_payload_15_3;
    _zz_dataOut_payload_16_49 <= _zz_dataOut_payload_16_48;
    _zz_dataOut_payload_17_4 <= _zz_dataOut_payload_17_3;
    _zz_dataOut_payload_18_7 <= _zz_dataOut_payload_18_6;
    _zz_dataOut_payload_19_4 <= _zz_dataOut_payload_19_3;
    _zz_dataOut_payload_20_13 <= _zz_dataOut_payload_20_12;
    _zz_dataOut_payload_21_4 <= _zz_dataOut_payload_21_3;
    _zz_dataOut_payload_22_7 <= _zz_dataOut_payload_22_6;
    _zz_dataOut_payload_23_4 <= _zz_dataOut_payload_23_3;
    _zz_dataOut_payload_24_25 <= _zz_dataOut_payload_24_24;
    _zz_dataOut_payload_25_4 <= _zz_dataOut_payload_25_3;
    _zz_dataOut_payload_26_7 <= _zz_dataOut_payload_26_6;
    _zz_dataOut_payload_27_4 <= _zz_dataOut_payload_27_3;
    _zz_dataOut_payload_28_13 <= _zz_dataOut_payload_28_12;
    _zz_dataOut_payload_29_4 <= _zz_dataOut_payload_29_3;
    _zz_dataOut_payload_30_7 <= _zz_dataOut_payload_30_6;
    _zz_dataOut_payload_31_4 <= _zz_dataOut_payload_31_3;
    _zz_dataOut_payload_32_97 <= _zz_dataOut_payload_32_96;
    _zz_dataOut_payload_33_4 <= _zz_dataOut_payload_33_3;
    _zz_dataOut_payload_34_7 <= _zz_dataOut_payload_34_6;
    _zz_dataOut_payload_35_4 <= _zz_dataOut_payload_35_3;
    _zz_dataOut_payload_36_13 <= _zz_dataOut_payload_36_12;
    _zz_dataOut_payload_37_4 <= _zz_dataOut_payload_37_3;
    _zz_dataOut_payload_38_7 <= _zz_dataOut_payload_38_6;
    _zz_dataOut_payload_39_4 <= _zz_dataOut_payload_39_3;
    _zz_dataOut_payload_40_25 <= _zz_dataOut_payload_40_24;
    _zz_dataOut_payload_41_4 <= _zz_dataOut_payload_41_3;
    _zz_dataOut_payload_42_7 <= _zz_dataOut_payload_42_6;
    _zz_dataOut_payload_43_4 <= _zz_dataOut_payload_43_3;
    _zz_dataOut_payload_44_13 <= _zz_dataOut_payload_44_12;
    _zz_dataOut_payload_45_4 <= _zz_dataOut_payload_45_3;
    _zz_dataOut_payload_46_7 <= _zz_dataOut_payload_46_6;
    _zz_dataOut_payload_47_4 <= _zz_dataOut_payload_47_3;
    _zz_dataOut_payload_48_49 <= _zz_dataOut_payload_48_48;
    _zz_dataOut_payload_49_4 <= _zz_dataOut_payload_49_3;
    _zz_dataOut_payload_50_7 <= _zz_dataOut_payload_50_6;
    _zz_dataOut_payload_51_4 <= _zz_dataOut_payload_51_3;
    _zz_dataOut_payload_52_13 <= _zz_dataOut_payload_52_12;
    _zz_dataOut_payload_53_4 <= _zz_dataOut_payload_53_3;
    _zz_dataOut_payload_54_7 <= _zz_dataOut_payload_54_6;
    _zz_dataOut_payload_55_4 <= _zz_dataOut_payload_55_3;
    _zz_dataOut_payload_56_25 <= _zz_dataOut_payload_56_24;
    _zz_dataOut_payload_57_4 <= _zz_dataOut_payload_57_3;
    _zz_dataOut_payload_58_7 <= _zz_dataOut_payload_58_6;
    _zz_dataOut_payload_59_4 <= _zz_dataOut_payload_59_3;
    _zz_dataOut_payload_60_13 <= _zz_dataOut_payload_60_12;
    _zz_dataOut_payload_61_4 <= _zz_dataOut_payload_61_3;
    _zz_dataOut_payload_62_7 <= _zz_dataOut_payload_62_6;
    _zz_dataOut_payload_63_4 <= _zz_dataOut_payload_63_3;
    _zz_dataOut_payload_64_189 <= (_zz_dataOut_payload_64_188 ? _zz_dataOut_payload_64_185 : _zz_dataOut_payload_64_187);
    _zz_dataOut_payload_65 <= (_zz_dataOut_payload_64_188 ? _zz_dataOut_payload_64_187 : _zz_dataOut_payload_64_185);
    _zz_dataOut_payload_66_3 <= (_zz_dataOut_payload_66_2 ? _zz_dataOut_payload_66 : _zz_dataOut_payload_66_1);
    _zz_dataOut_payload_67 <= (_zz_dataOut_payload_66_2 ? _zz_dataOut_payload_66_1 : _zz_dataOut_payload_66);
    _zz_dataOut_payload_68_9 <= (_zz_dataOut_payload_68_8 ? _zz_dataOut_payload_68_5 : _zz_dataOut_payload_68_7);
    _zz_dataOut_payload_69 <= (_zz_dataOut_payload_68_8 ? _zz_dataOut_payload_68_7 : _zz_dataOut_payload_68_5);
    _zz_dataOut_payload_70_3 <= (_zz_dataOut_payload_70_2 ? _zz_dataOut_payload_70 : _zz_dataOut_payload_70_1);
    _zz_dataOut_payload_71 <= (_zz_dataOut_payload_70_2 ? _zz_dataOut_payload_70_1 : _zz_dataOut_payload_70);
    _zz_dataOut_payload_64_190 <= _zz_dataOut_payload_64_189;
    _zz_dataOut_payload_65_1 <= _zz_dataOut_payload_65;
    _zz_dataOut_payload_66_4 <= _zz_dataOut_payload_66_3;
    _zz_dataOut_payload_67_1 <= _zz_dataOut_payload_67;
    _zz_dataOut_payload_68_10 <= _zz_dataOut_payload_68_9;
    _zz_dataOut_payload_69_1 <= _zz_dataOut_payload_69;
    _zz_dataOut_payload_70_4 <= _zz_dataOut_payload_70_3;
    _zz_dataOut_payload_71_1 <= _zz_dataOut_payload_71;
    _zz_dataOut_payload_72_21 <= (_zz_dataOut_payload_72_20 ? _zz_dataOut_payload_72_17 : _zz_dataOut_payload_72_19);
    _zz_dataOut_payload_73 <= (_zz_dataOut_payload_72_20 ? _zz_dataOut_payload_72_19 : _zz_dataOut_payload_72_17);
    _zz_dataOut_payload_74_3 <= (_zz_dataOut_payload_74_2 ? _zz_dataOut_payload_74 : _zz_dataOut_payload_74_1);
    _zz_dataOut_payload_75 <= (_zz_dataOut_payload_74_2 ? _zz_dataOut_payload_74_1 : _zz_dataOut_payload_74);
    _zz_dataOut_payload_76_9 <= (_zz_dataOut_payload_76_8 ? _zz_dataOut_payload_76_5 : _zz_dataOut_payload_76_7);
    _zz_dataOut_payload_77 <= (_zz_dataOut_payload_76_8 ? _zz_dataOut_payload_76_7 : _zz_dataOut_payload_76_5);
    _zz_dataOut_payload_78_3 <= (_zz_dataOut_payload_78_2 ? _zz_dataOut_payload_78 : _zz_dataOut_payload_78_1);
    _zz_dataOut_payload_79 <= (_zz_dataOut_payload_78_2 ? _zz_dataOut_payload_78_1 : _zz_dataOut_payload_78);
    _zz_dataOut_payload_72_22 <= _zz_dataOut_payload_72_21;
    _zz_dataOut_payload_73_1 <= _zz_dataOut_payload_73;
    _zz_dataOut_payload_74_4 <= _zz_dataOut_payload_74_3;
    _zz_dataOut_payload_75_1 <= _zz_dataOut_payload_75;
    _zz_dataOut_payload_76_10 <= _zz_dataOut_payload_76_9;
    _zz_dataOut_payload_77_1 <= _zz_dataOut_payload_77;
    _zz_dataOut_payload_78_4 <= _zz_dataOut_payload_78_3;
    _zz_dataOut_payload_79_1 <= _zz_dataOut_payload_79;
    _zz_dataOut_payload_64_191 <= _zz_dataOut_payload_64_190;
    _zz_dataOut_payload_65_2 <= _zz_dataOut_payload_65_1;
    _zz_dataOut_payload_66_5 <= _zz_dataOut_payload_66_4;
    _zz_dataOut_payload_67_2 <= _zz_dataOut_payload_67_1;
    _zz_dataOut_payload_68_11 <= _zz_dataOut_payload_68_10;
    _zz_dataOut_payload_69_2 <= _zz_dataOut_payload_69_1;
    _zz_dataOut_payload_70_5 <= _zz_dataOut_payload_70_4;
    _zz_dataOut_payload_71_2 <= _zz_dataOut_payload_71_1;
    _zz_dataOut_payload_72_23 <= _zz_dataOut_payload_72_22;
    _zz_dataOut_payload_73_2 <= _zz_dataOut_payload_73_1;
    _zz_dataOut_payload_74_5 <= _zz_dataOut_payload_74_4;
    _zz_dataOut_payload_75_2 <= _zz_dataOut_payload_75_1;
    _zz_dataOut_payload_76_11 <= _zz_dataOut_payload_76_10;
    _zz_dataOut_payload_77_2 <= _zz_dataOut_payload_77_1;
    _zz_dataOut_payload_78_5 <= _zz_dataOut_payload_78_4;
    _zz_dataOut_payload_79_2 <= _zz_dataOut_payload_79_1;
    _zz_dataOut_payload_80_45 <= (_zz_dataOut_payload_80_44 ? _zz_dataOut_payload_80_41 : _zz_dataOut_payload_80_43);
    _zz_dataOut_payload_81 <= (_zz_dataOut_payload_80_44 ? _zz_dataOut_payload_80_43 : _zz_dataOut_payload_80_41);
    _zz_dataOut_payload_82_3 <= (_zz_dataOut_payload_82_2 ? _zz_dataOut_payload_82 : _zz_dataOut_payload_82_1);
    _zz_dataOut_payload_83 <= (_zz_dataOut_payload_82_2 ? _zz_dataOut_payload_82_1 : _zz_dataOut_payload_82);
    _zz_dataOut_payload_84_9 <= (_zz_dataOut_payload_84_8 ? _zz_dataOut_payload_84_5 : _zz_dataOut_payload_84_7);
    _zz_dataOut_payload_85 <= (_zz_dataOut_payload_84_8 ? _zz_dataOut_payload_84_7 : _zz_dataOut_payload_84_5);
    _zz_dataOut_payload_86_3 <= (_zz_dataOut_payload_86_2 ? _zz_dataOut_payload_86 : _zz_dataOut_payload_86_1);
    _zz_dataOut_payload_87 <= (_zz_dataOut_payload_86_2 ? _zz_dataOut_payload_86_1 : _zz_dataOut_payload_86);
    _zz_dataOut_payload_80_46 <= _zz_dataOut_payload_80_45;
    _zz_dataOut_payload_81_1 <= _zz_dataOut_payload_81;
    _zz_dataOut_payload_82_4 <= _zz_dataOut_payload_82_3;
    _zz_dataOut_payload_83_1 <= _zz_dataOut_payload_83;
    _zz_dataOut_payload_84_10 <= _zz_dataOut_payload_84_9;
    _zz_dataOut_payload_85_1 <= _zz_dataOut_payload_85;
    _zz_dataOut_payload_86_4 <= _zz_dataOut_payload_86_3;
    _zz_dataOut_payload_87_1 <= _zz_dataOut_payload_87;
    _zz_dataOut_payload_88_21 <= (_zz_dataOut_payload_88_20 ? _zz_dataOut_payload_88_17 : _zz_dataOut_payload_88_19);
    _zz_dataOut_payload_89 <= (_zz_dataOut_payload_88_20 ? _zz_dataOut_payload_88_19 : _zz_dataOut_payload_88_17);
    _zz_dataOut_payload_90_3 <= (_zz_dataOut_payload_90_2 ? _zz_dataOut_payload_90 : _zz_dataOut_payload_90_1);
    _zz_dataOut_payload_91 <= (_zz_dataOut_payload_90_2 ? _zz_dataOut_payload_90_1 : _zz_dataOut_payload_90);
    _zz_dataOut_payload_92_9 <= (_zz_dataOut_payload_92_8 ? _zz_dataOut_payload_92_5 : _zz_dataOut_payload_92_7);
    _zz_dataOut_payload_93 <= (_zz_dataOut_payload_92_8 ? _zz_dataOut_payload_92_7 : _zz_dataOut_payload_92_5);
    _zz_dataOut_payload_94_3 <= (_zz_dataOut_payload_94_2 ? _zz_dataOut_payload_94 : _zz_dataOut_payload_94_1);
    _zz_dataOut_payload_95 <= (_zz_dataOut_payload_94_2 ? _zz_dataOut_payload_94_1 : _zz_dataOut_payload_94);
    _zz_dataOut_payload_88_22 <= _zz_dataOut_payload_88_21;
    _zz_dataOut_payload_89_1 <= _zz_dataOut_payload_89;
    _zz_dataOut_payload_90_4 <= _zz_dataOut_payload_90_3;
    _zz_dataOut_payload_91_1 <= _zz_dataOut_payload_91;
    _zz_dataOut_payload_92_10 <= _zz_dataOut_payload_92_9;
    _zz_dataOut_payload_93_1 <= _zz_dataOut_payload_93;
    _zz_dataOut_payload_94_4 <= _zz_dataOut_payload_94_3;
    _zz_dataOut_payload_95_1 <= _zz_dataOut_payload_95;
    _zz_dataOut_payload_80_47 <= _zz_dataOut_payload_80_46;
    _zz_dataOut_payload_81_2 <= _zz_dataOut_payload_81_1;
    _zz_dataOut_payload_82_5 <= _zz_dataOut_payload_82_4;
    _zz_dataOut_payload_83_2 <= _zz_dataOut_payload_83_1;
    _zz_dataOut_payload_84_11 <= _zz_dataOut_payload_84_10;
    _zz_dataOut_payload_85_2 <= _zz_dataOut_payload_85_1;
    _zz_dataOut_payload_86_5 <= _zz_dataOut_payload_86_4;
    _zz_dataOut_payload_87_2 <= _zz_dataOut_payload_87_1;
    _zz_dataOut_payload_88_23 <= _zz_dataOut_payload_88_22;
    _zz_dataOut_payload_89_2 <= _zz_dataOut_payload_89_1;
    _zz_dataOut_payload_90_5 <= _zz_dataOut_payload_90_4;
    _zz_dataOut_payload_91_2 <= _zz_dataOut_payload_91_1;
    _zz_dataOut_payload_92_11 <= _zz_dataOut_payload_92_10;
    _zz_dataOut_payload_93_2 <= _zz_dataOut_payload_93_1;
    _zz_dataOut_payload_94_5 <= _zz_dataOut_payload_94_4;
    _zz_dataOut_payload_95_2 <= _zz_dataOut_payload_95_1;
    _zz_dataOut_payload_64_192 <= _zz_dataOut_payload_64_191;
    _zz_dataOut_payload_65_3 <= _zz_dataOut_payload_65_2;
    _zz_dataOut_payload_66_6 <= _zz_dataOut_payload_66_5;
    _zz_dataOut_payload_67_3 <= _zz_dataOut_payload_67_2;
    _zz_dataOut_payload_68_12 <= _zz_dataOut_payload_68_11;
    _zz_dataOut_payload_69_3 <= _zz_dataOut_payload_69_2;
    _zz_dataOut_payload_70_6 <= _zz_dataOut_payload_70_5;
    _zz_dataOut_payload_71_3 <= _zz_dataOut_payload_71_2;
    _zz_dataOut_payload_72_24 <= _zz_dataOut_payload_72_23;
    _zz_dataOut_payload_73_3 <= _zz_dataOut_payload_73_2;
    _zz_dataOut_payload_74_6 <= _zz_dataOut_payload_74_5;
    _zz_dataOut_payload_75_3 <= _zz_dataOut_payload_75_2;
    _zz_dataOut_payload_76_12 <= _zz_dataOut_payload_76_11;
    _zz_dataOut_payload_77_3 <= _zz_dataOut_payload_77_2;
    _zz_dataOut_payload_78_6 <= _zz_dataOut_payload_78_5;
    _zz_dataOut_payload_79_3 <= _zz_dataOut_payload_79_2;
    _zz_dataOut_payload_80_48 <= _zz_dataOut_payload_80_47;
    _zz_dataOut_payload_81_3 <= _zz_dataOut_payload_81_2;
    _zz_dataOut_payload_82_6 <= _zz_dataOut_payload_82_5;
    _zz_dataOut_payload_83_3 <= _zz_dataOut_payload_83_2;
    _zz_dataOut_payload_84_12 <= _zz_dataOut_payload_84_11;
    _zz_dataOut_payload_85_3 <= _zz_dataOut_payload_85_2;
    _zz_dataOut_payload_86_6 <= _zz_dataOut_payload_86_5;
    _zz_dataOut_payload_87_3 <= _zz_dataOut_payload_87_2;
    _zz_dataOut_payload_88_24 <= _zz_dataOut_payload_88_23;
    _zz_dataOut_payload_89_3 <= _zz_dataOut_payload_89_2;
    _zz_dataOut_payload_90_6 <= _zz_dataOut_payload_90_5;
    _zz_dataOut_payload_91_3 <= _zz_dataOut_payload_91_2;
    _zz_dataOut_payload_92_12 <= _zz_dataOut_payload_92_11;
    _zz_dataOut_payload_93_3 <= _zz_dataOut_payload_93_2;
    _zz_dataOut_payload_94_6 <= _zz_dataOut_payload_94_5;
    _zz_dataOut_payload_95_3 <= _zz_dataOut_payload_95_2;
    _zz_dataOut_payload_96_93 <= (_zz_dataOut_payload_96_92 ? _zz_dataOut_payload_96_89 : _zz_dataOut_payload_96_91);
    _zz_dataOut_payload_97 <= (_zz_dataOut_payload_96_92 ? _zz_dataOut_payload_96_91 : _zz_dataOut_payload_96_89);
    _zz_dataOut_payload_98_3 <= (_zz_dataOut_payload_98_2 ? _zz_dataOut_payload_98 : _zz_dataOut_payload_98_1);
    _zz_dataOut_payload_99 <= (_zz_dataOut_payload_98_2 ? _zz_dataOut_payload_98_1 : _zz_dataOut_payload_98);
    _zz_dataOut_payload_100_9 <= (_zz_dataOut_payload_100_8 ? _zz_dataOut_payload_100_5 : _zz_dataOut_payload_100_7);
    _zz_dataOut_payload_101 <= (_zz_dataOut_payload_100_8 ? _zz_dataOut_payload_100_7 : _zz_dataOut_payload_100_5);
    _zz_dataOut_payload_102_3 <= (_zz_dataOut_payload_102_2 ? _zz_dataOut_payload_102 : _zz_dataOut_payload_102_1);
    _zz_dataOut_payload_103 <= (_zz_dataOut_payload_102_2 ? _zz_dataOut_payload_102_1 : _zz_dataOut_payload_102);
    _zz_dataOut_payload_96_94 <= _zz_dataOut_payload_96_93;
    _zz_dataOut_payload_97_1 <= _zz_dataOut_payload_97;
    _zz_dataOut_payload_98_4 <= _zz_dataOut_payload_98_3;
    _zz_dataOut_payload_99_1 <= _zz_dataOut_payload_99;
    _zz_dataOut_payload_100_10 <= _zz_dataOut_payload_100_9;
    _zz_dataOut_payload_101_1 <= _zz_dataOut_payload_101;
    _zz_dataOut_payload_102_4 <= _zz_dataOut_payload_102_3;
    _zz_dataOut_payload_103_1 <= _zz_dataOut_payload_103;
    _zz_dataOut_payload_104_21 <= (_zz_dataOut_payload_104_20 ? _zz_dataOut_payload_104_17 : _zz_dataOut_payload_104_19);
    _zz_dataOut_payload_105 <= (_zz_dataOut_payload_104_20 ? _zz_dataOut_payload_104_19 : _zz_dataOut_payload_104_17);
    _zz_dataOut_payload_106_3 <= (_zz_dataOut_payload_106_2 ? _zz_dataOut_payload_106 : _zz_dataOut_payload_106_1);
    _zz_dataOut_payload_107 <= (_zz_dataOut_payload_106_2 ? _zz_dataOut_payload_106_1 : _zz_dataOut_payload_106);
    _zz_dataOut_payload_108_9 <= (_zz_dataOut_payload_108_8 ? _zz_dataOut_payload_108_5 : _zz_dataOut_payload_108_7);
    _zz_dataOut_payload_109 <= (_zz_dataOut_payload_108_8 ? _zz_dataOut_payload_108_7 : _zz_dataOut_payload_108_5);
    _zz_dataOut_payload_110_3 <= (_zz_dataOut_payload_110_2 ? _zz_dataOut_payload_110 : _zz_dataOut_payload_110_1);
    _zz_dataOut_payload_111 <= (_zz_dataOut_payload_110_2 ? _zz_dataOut_payload_110_1 : _zz_dataOut_payload_110);
    _zz_dataOut_payload_104_22 <= _zz_dataOut_payload_104_21;
    _zz_dataOut_payload_105_1 <= _zz_dataOut_payload_105;
    _zz_dataOut_payload_106_4 <= _zz_dataOut_payload_106_3;
    _zz_dataOut_payload_107_1 <= _zz_dataOut_payload_107;
    _zz_dataOut_payload_108_10 <= _zz_dataOut_payload_108_9;
    _zz_dataOut_payload_109_1 <= _zz_dataOut_payload_109;
    _zz_dataOut_payload_110_4 <= _zz_dataOut_payload_110_3;
    _zz_dataOut_payload_111_1 <= _zz_dataOut_payload_111;
    _zz_dataOut_payload_96_95 <= _zz_dataOut_payload_96_94;
    _zz_dataOut_payload_97_2 <= _zz_dataOut_payload_97_1;
    _zz_dataOut_payload_98_5 <= _zz_dataOut_payload_98_4;
    _zz_dataOut_payload_99_2 <= _zz_dataOut_payload_99_1;
    _zz_dataOut_payload_100_11 <= _zz_dataOut_payload_100_10;
    _zz_dataOut_payload_101_2 <= _zz_dataOut_payload_101_1;
    _zz_dataOut_payload_102_5 <= _zz_dataOut_payload_102_4;
    _zz_dataOut_payload_103_2 <= _zz_dataOut_payload_103_1;
    _zz_dataOut_payload_104_23 <= _zz_dataOut_payload_104_22;
    _zz_dataOut_payload_105_2 <= _zz_dataOut_payload_105_1;
    _zz_dataOut_payload_106_5 <= _zz_dataOut_payload_106_4;
    _zz_dataOut_payload_107_2 <= _zz_dataOut_payload_107_1;
    _zz_dataOut_payload_108_11 <= _zz_dataOut_payload_108_10;
    _zz_dataOut_payload_109_2 <= _zz_dataOut_payload_109_1;
    _zz_dataOut_payload_110_5 <= _zz_dataOut_payload_110_4;
    _zz_dataOut_payload_111_2 <= _zz_dataOut_payload_111_1;
    _zz_dataOut_payload_112_45 <= (_zz_dataOut_payload_112_44 ? _zz_dataOut_payload_112_41 : _zz_dataOut_payload_112_43);
    _zz_dataOut_payload_113 <= (_zz_dataOut_payload_112_44 ? _zz_dataOut_payload_112_43 : _zz_dataOut_payload_112_41);
    _zz_dataOut_payload_114_3 <= (_zz_dataOut_payload_114_2 ? _zz_dataOut_payload_114 : _zz_dataOut_payload_114_1);
    _zz_dataOut_payload_115 <= (_zz_dataOut_payload_114_2 ? _zz_dataOut_payload_114_1 : _zz_dataOut_payload_114);
    _zz_dataOut_payload_116_9 <= (_zz_dataOut_payload_116_8 ? _zz_dataOut_payload_116_5 : _zz_dataOut_payload_116_7);
    _zz_dataOut_payload_117 <= (_zz_dataOut_payload_116_8 ? _zz_dataOut_payload_116_7 : _zz_dataOut_payload_116_5);
    _zz_dataOut_payload_118_3 <= (_zz_dataOut_payload_118_2 ? _zz_dataOut_payload_118 : _zz_dataOut_payload_118_1);
    _zz_dataOut_payload_119 <= (_zz_dataOut_payload_118_2 ? _zz_dataOut_payload_118_1 : _zz_dataOut_payload_118);
    _zz_dataOut_payload_112_46 <= _zz_dataOut_payload_112_45;
    _zz_dataOut_payload_113_1 <= _zz_dataOut_payload_113;
    _zz_dataOut_payload_114_4 <= _zz_dataOut_payload_114_3;
    _zz_dataOut_payload_115_1 <= _zz_dataOut_payload_115;
    _zz_dataOut_payload_116_10 <= _zz_dataOut_payload_116_9;
    _zz_dataOut_payload_117_1 <= _zz_dataOut_payload_117;
    _zz_dataOut_payload_118_4 <= _zz_dataOut_payload_118_3;
    _zz_dataOut_payload_119_1 <= _zz_dataOut_payload_119;
    _zz_dataOut_payload_120_21 <= (_zz_dataOut_payload_120_20 ? _zz_dataOut_payload_120_17 : _zz_dataOut_payload_120_19);
    _zz_dataOut_payload_121 <= (_zz_dataOut_payload_120_20 ? _zz_dataOut_payload_120_19 : _zz_dataOut_payload_120_17);
    _zz_dataOut_payload_122_3 <= (_zz_dataOut_payload_122_2 ? _zz_dataOut_payload_122 : _zz_dataOut_payload_122_1);
    _zz_dataOut_payload_123 <= (_zz_dataOut_payload_122_2 ? _zz_dataOut_payload_122_1 : _zz_dataOut_payload_122);
    _zz_dataOut_payload_124_9 <= (_zz_dataOut_payload_124_8 ? _zz_dataOut_payload_124_5 : _zz_dataOut_payload_124_7);
    _zz_dataOut_payload_125 <= (_zz_dataOut_payload_124_8 ? _zz_dataOut_payload_124_7 : _zz_dataOut_payload_124_5);
    _zz_dataOut_payload_126_3 <= (_zz_dataOut_payload_126_2 ? _zz_dataOut_payload_126 : _zz_dataOut_payload_126_1);
    _zz_dataOut_payload_127 <= (_zz_dataOut_payload_126_2 ? _zz_dataOut_payload_126_1 : _zz_dataOut_payload_126);
    _zz_dataOut_payload_120_22 <= _zz_dataOut_payload_120_21;
    _zz_dataOut_payload_121_1 <= _zz_dataOut_payload_121;
    _zz_dataOut_payload_122_4 <= _zz_dataOut_payload_122_3;
    _zz_dataOut_payload_123_1 <= _zz_dataOut_payload_123;
    _zz_dataOut_payload_124_10 <= _zz_dataOut_payload_124_9;
    _zz_dataOut_payload_125_1 <= _zz_dataOut_payload_125;
    _zz_dataOut_payload_126_4 <= _zz_dataOut_payload_126_3;
    _zz_dataOut_payload_127_1 <= _zz_dataOut_payload_127;
    _zz_dataOut_payload_112_47 <= _zz_dataOut_payload_112_46;
    _zz_dataOut_payload_113_2 <= _zz_dataOut_payload_113_1;
    _zz_dataOut_payload_114_5 <= _zz_dataOut_payload_114_4;
    _zz_dataOut_payload_115_2 <= _zz_dataOut_payload_115_1;
    _zz_dataOut_payload_116_11 <= _zz_dataOut_payload_116_10;
    _zz_dataOut_payload_117_2 <= _zz_dataOut_payload_117_1;
    _zz_dataOut_payload_118_5 <= _zz_dataOut_payload_118_4;
    _zz_dataOut_payload_119_2 <= _zz_dataOut_payload_119_1;
    _zz_dataOut_payload_120_23 <= _zz_dataOut_payload_120_22;
    _zz_dataOut_payload_121_2 <= _zz_dataOut_payload_121_1;
    _zz_dataOut_payload_122_5 <= _zz_dataOut_payload_122_4;
    _zz_dataOut_payload_123_2 <= _zz_dataOut_payload_123_1;
    _zz_dataOut_payload_124_11 <= _zz_dataOut_payload_124_10;
    _zz_dataOut_payload_125_2 <= _zz_dataOut_payload_125_1;
    _zz_dataOut_payload_126_5 <= _zz_dataOut_payload_126_4;
    _zz_dataOut_payload_127_2 <= _zz_dataOut_payload_127_1;
    _zz_dataOut_payload_96_96 <= _zz_dataOut_payload_96_95;
    _zz_dataOut_payload_97_3 <= _zz_dataOut_payload_97_2;
    _zz_dataOut_payload_98_6 <= _zz_dataOut_payload_98_5;
    _zz_dataOut_payload_99_3 <= _zz_dataOut_payload_99_2;
    _zz_dataOut_payload_100_12 <= _zz_dataOut_payload_100_11;
    _zz_dataOut_payload_101_3 <= _zz_dataOut_payload_101_2;
    _zz_dataOut_payload_102_6 <= _zz_dataOut_payload_102_5;
    _zz_dataOut_payload_103_3 <= _zz_dataOut_payload_103_2;
    _zz_dataOut_payload_104_24 <= _zz_dataOut_payload_104_23;
    _zz_dataOut_payload_105_3 <= _zz_dataOut_payload_105_2;
    _zz_dataOut_payload_106_6 <= _zz_dataOut_payload_106_5;
    _zz_dataOut_payload_107_3 <= _zz_dataOut_payload_107_2;
    _zz_dataOut_payload_108_12 <= _zz_dataOut_payload_108_11;
    _zz_dataOut_payload_109_3 <= _zz_dataOut_payload_109_2;
    _zz_dataOut_payload_110_6 <= _zz_dataOut_payload_110_5;
    _zz_dataOut_payload_111_3 <= _zz_dataOut_payload_111_2;
    _zz_dataOut_payload_112_48 <= _zz_dataOut_payload_112_47;
    _zz_dataOut_payload_113_3 <= _zz_dataOut_payload_113_2;
    _zz_dataOut_payload_114_6 <= _zz_dataOut_payload_114_5;
    _zz_dataOut_payload_115_3 <= _zz_dataOut_payload_115_2;
    _zz_dataOut_payload_116_12 <= _zz_dataOut_payload_116_11;
    _zz_dataOut_payload_117_3 <= _zz_dataOut_payload_117_2;
    _zz_dataOut_payload_118_6 <= _zz_dataOut_payload_118_5;
    _zz_dataOut_payload_119_3 <= _zz_dataOut_payload_119_2;
    _zz_dataOut_payload_120_24 <= _zz_dataOut_payload_120_23;
    _zz_dataOut_payload_121_3 <= _zz_dataOut_payload_121_2;
    _zz_dataOut_payload_122_6 <= _zz_dataOut_payload_122_5;
    _zz_dataOut_payload_123_3 <= _zz_dataOut_payload_123_2;
    _zz_dataOut_payload_124_12 <= _zz_dataOut_payload_124_11;
    _zz_dataOut_payload_125_3 <= _zz_dataOut_payload_125_2;
    _zz_dataOut_payload_126_6 <= _zz_dataOut_payload_126_5;
    _zz_dataOut_payload_127_3 <= _zz_dataOut_payload_127_2;
    _zz_dataOut_payload_64_193 <= _zz_dataOut_payload_64_192;
    _zz_dataOut_payload_65_4 <= _zz_dataOut_payload_65_3;
    _zz_dataOut_payload_66_7 <= _zz_dataOut_payload_66_6;
    _zz_dataOut_payload_67_4 <= _zz_dataOut_payload_67_3;
    _zz_dataOut_payload_68_13 <= _zz_dataOut_payload_68_12;
    _zz_dataOut_payload_69_4 <= _zz_dataOut_payload_69_3;
    _zz_dataOut_payload_70_7 <= _zz_dataOut_payload_70_6;
    _zz_dataOut_payload_71_4 <= _zz_dataOut_payload_71_3;
    _zz_dataOut_payload_72_25 <= _zz_dataOut_payload_72_24;
    _zz_dataOut_payload_73_4 <= _zz_dataOut_payload_73_3;
    _zz_dataOut_payload_74_7 <= _zz_dataOut_payload_74_6;
    _zz_dataOut_payload_75_4 <= _zz_dataOut_payload_75_3;
    _zz_dataOut_payload_76_13 <= _zz_dataOut_payload_76_12;
    _zz_dataOut_payload_77_4 <= _zz_dataOut_payload_77_3;
    _zz_dataOut_payload_78_7 <= _zz_dataOut_payload_78_6;
    _zz_dataOut_payload_79_4 <= _zz_dataOut_payload_79_3;
    _zz_dataOut_payload_80_49 <= _zz_dataOut_payload_80_48;
    _zz_dataOut_payload_81_4 <= _zz_dataOut_payload_81_3;
    _zz_dataOut_payload_82_7 <= _zz_dataOut_payload_82_6;
    _zz_dataOut_payload_83_4 <= _zz_dataOut_payload_83_3;
    _zz_dataOut_payload_84_13 <= _zz_dataOut_payload_84_12;
    _zz_dataOut_payload_85_4 <= _zz_dataOut_payload_85_3;
    _zz_dataOut_payload_86_7 <= _zz_dataOut_payload_86_6;
    _zz_dataOut_payload_87_4 <= _zz_dataOut_payload_87_3;
    _zz_dataOut_payload_88_25 <= _zz_dataOut_payload_88_24;
    _zz_dataOut_payload_89_4 <= _zz_dataOut_payload_89_3;
    _zz_dataOut_payload_90_7 <= _zz_dataOut_payload_90_6;
    _zz_dataOut_payload_91_4 <= _zz_dataOut_payload_91_3;
    _zz_dataOut_payload_92_13 <= _zz_dataOut_payload_92_12;
    _zz_dataOut_payload_93_4 <= _zz_dataOut_payload_93_3;
    _zz_dataOut_payload_94_7 <= _zz_dataOut_payload_94_6;
    _zz_dataOut_payload_95_4 <= _zz_dataOut_payload_95_3;
    _zz_dataOut_payload_96_97 <= _zz_dataOut_payload_96_96;
    _zz_dataOut_payload_97_4 <= _zz_dataOut_payload_97_3;
    _zz_dataOut_payload_98_7 <= _zz_dataOut_payload_98_6;
    _zz_dataOut_payload_99_4 <= _zz_dataOut_payload_99_3;
    _zz_dataOut_payload_100_13 <= _zz_dataOut_payload_100_12;
    _zz_dataOut_payload_101_4 <= _zz_dataOut_payload_101_3;
    _zz_dataOut_payload_102_7 <= _zz_dataOut_payload_102_6;
    _zz_dataOut_payload_103_4 <= _zz_dataOut_payload_103_3;
    _zz_dataOut_payload_104_25 <= _zz_dataOut_payload_104_24;
    _zz_dataOut_payload_105_4 <= _zz_dataOut_payload_105_3;
    _zz_dataOut_payload_106_7 <= _zz_dataOut_payload_106_6;
    _zz_dataOut_payload_107_4 <= _zz_dataOut_payload_107_3;
    _zz_dataOut_payload_108_13 <= _zz_dataOut_payload_108_12;
    _zz_dataOut_payload_109_4 <= _zz_dataOut_payload_109_3;
    _zz_dataOut_payload_110_7 <= _zz_dataOut_payload_110_6;
    _zz_dataOut_payload_111_4 <= _zz_dataOut_payload_111_3;
    _zz_dataOut_payload_112_49 <= _zz_dataOut_payload_112_48;
    _zz_dataOut_payload_113_4 <= _zz_dataOut_payload_113_3;
    _zz_dataOut_payload_114_7 <= _zz_dataOut_payload_114_6;
    _zz_dataOut_payload_115_4 <= _zz_dataOut_payload_115_3;
    _zz_dataOut_payload_116_13 <= _zz_dataOut_payload_116_12;
    _zz_dataOut_payload_117_4 <= _zz_dataOut_payload_117_3;
    _zz_dataOut_payload_118_7 <= _zz_dataOut_payload_118_6;
    _zz_dataOut_payload_119_4 <= _zz_dataOut_payload_119_3;
    _zz_dataOut_payload_120_25 <= _zz_dataOut_payload_120_24;
    _zz_dataOut_payload_121_4 <= _zz_dataOut_payload_121_3;
    _zz_dataOut_payload_122_7 <= _zz_dataOut_payload_122_6;
    _zz_dataOut_payload_123_4 <= _zz_dataOut_payload_123_3;
    _zz_dataOut_payload_124_13 <= _zz_dataOut_payload_124_12;
    _zz_dataOut_payload_125_4 <= _zz_dataOut_payload_125_3;
    _zz_dataOut_payload_126_7 <= _zz_dataOut_payload_126_6;
    _zz_dataOut_payload_127_4 <= _zz_dataOut_payload_127_3;
    _zz_dataOut_payload_0_16642 <= _zz_dataOut_payload_0_16641;
    _zz_dataOut_payload_1_5 <= _zz_dataOut_payload_1_4;
    _zz_dataOut_payload_2_8 <= _zz_dataOut_payload_2_7;
    _zz_dataOut_payload_3_5 <= _zz_dataOut_payload_3_4;
    _zz_dataOut_payload_4_14 <= _zz_dataOut_payload_4_13;
    _zz_dataOut_payload_5_5 <= _zz_dataOut_payload_5_4;
    _zz_dataOut_payload_6_8 <= _zz_dataOut_payload_6_7;
    _zz_dataOut_payload_7_5 <= _zz_dataOut_payload_7_4;
    _zz_dataOut_payload_8_26 <= _zz_dataOut_payload_8_25;
    _zz_dataOut_payload_9_5 <= _zz_dataOut_payload_9_4;
    _zz_dataOut_payload_10_8 <= _zz_dataOut_payload_10_7;
    _zz_dataOut_payload_11_5 <= _zz_dataOut_payload_11_4;
    _zz_dataOut_payload_12_14 <= _zz_dataOut_payload_12_13;
    _zz_dataOut_payload_13_5 <= _zz_dataOut_payload_13_4;
    _zz_dataOut_payload_14_8 <= _zz_dataOut_payload_14_7;
    _zz_dataOut_payload_15_5 <= _zz_dataOut_payload_15_4;
    _zz_dataOut_payload_16_50 <= _zz_dataOut_payload_16_49;
    _zz_dataOut_payload_17_5 <= _zz_dataOut_payload_17_4;
    _zz_dataOut_payload_18_8 <= _zz_dataOut_payload_18_7;
    _zz_dataOut_payload_19_5 <= _zz_dataOut_payload_19_4;
    _zz_dataOut_payload_20_14 <= _zz_dataOut_payload_20_13;
    _zz_dataOut_payload_21_5 <= _zz_dataOut_payload_21_4;
    _zz_dataOut_payload_22_8 <= _zz_dataOut_payload_22_7;
    _zz_dataOut_payload_23_5 <= _zz_dataOut_payload_23_4;
    _zz_dataOut_payload_24_26 <= _zz_dataOut_payload_24_25;
    _zz_dataOut_payload_25_5 <= _zz_dataOut_payload_25_4;
    _zz_dataOut_payload_26_8 <= _zz_dataOut_payload_26_7;
    _zz_dataOut_payload_27_5 <= _zz_dataOut_payload_27_4;
    _zz_dataOut_payload_28_14 <= _zz_dataOut_payload_28_13;
    _zz_dataOut_payload_29_5 <= _zz_dataOut_payload_29_4;
    _zz_dataOut_payload_30_8 <= _zz_dataOut_payload_30_7;
    _zz_dataOut_payload_31_5 <= _zz_dataOut_payload_31_4;
    _zz_dataOut_payload_32_98 <= _zz_dataOut_payload_32_97;
    _zz_dataOut_payload_33_5 <= _zz_dataOut_payload_33_4;
    _zz_dataOut_payload_34_8 <= _zz_dataOut_payload_34_7;
    _zz_dataOut_payload_35_5 <= _zz_dataOut_payload_35_4;
    _zz_dataOut_payload_36_14 <= _zz_dataOut_payload_36_13;
    _zz_dataOut_payload_37_5 <= _zz_dataOut_payload_37_4;
    _zz_dataOut_payload_38_8 <= _zz_dataOut_payload_38_7;
    _zz_dataOut_payload_39_5 <= _zz_dataOut_payload_39_4;
    _zz_dataOut_payload_40_26 <= _zz_dataOut_payload_40_25;
    _zz_dataOut_payload_41_5 <= _zz_dataOut_payload_41_4;
    _zz_dataOut_payload_42_8 <= _zz_dataOut_payload_42_7;
    _zz_dataOut_payload_43_5 <= _zz_dataOut_payload_43_4;
    _zz_dataOut_payload_44_14 <= _zz_dataOut_payload_44_13;
    _zz_dataOut_payload_45_5 <= _zz_dataOut_payload_45_4;
    _zz_dataOut_payload_46_8 <= _zz_dataOut_payload_46_7;
    _zz_dataOut_payload_47_5 <= _zz_dataOut_payload_47_4;
    _zz_dataOut_payload_48_50 <= _zz_dataOut_payload_48_49;
    _zz_dataOut_payload_49_5 <= _zz_dataOut_payload_49_4;
    _zz_dataOut_payload_50_8 <= _zz_dataOut_payload_50_7;
    _zz_dataOut_payload_51_5 <= _zz_dataOut_payload_51_4;
    _zz_dataOut_payload_52_14 <= _zz_dataOut_payload_52_13;
    _zz_dataOut_payload_53_5 <= _zz_dataOut_payload_53_4;
    _zz_dataOut_payload_54_8 <= _zz_dataOut_payload_54_7;
    _zz_dataOut_payload_55_5 <= _zz_dataOut_payload_55_4;
    _zz_dataOut_payload_56_26 <= _zz_dataOut_payload_56_25;
    _zz_dataOut_payload_57_5 <= _zz_dataOut_payload_57_4;
    _zz_dataOut_payload_58_8 <= _zz_dataOut_payload_58_7;
    _zz_dataOut_payload_59_5 <= _zz_dataOut_payload_59_4;
    _zz_dataOut_payload_60_14 <= _zz_dataOut_payload_60_13;
    _zz_dataOut_payload_61_5 <= _zz_dataOut_payload_61_4;
    _zz_dataOut_payload_62_8 <= _zz_dataOut_payload_62_7;
    _zz_dataOut_payload_63_5 <= _zz_dataOut_payload_63_4;
    _zz_dataOut_payload_64_194 <= _zz_dataOut_payload_64_193;
    _zz_dataOut_payload_65_5 <= _zz_dataOut_payload_65_4;
    _zz_dataOut_payload_66_8 <= _zz_dataOut_payload_66_7;
    _zz_dataOut_payload_67_5 <= _zz_dataOut_payload_67_4;
    _zz_dataOut_payload_68_14 <= _zz_dataOut_payload_68_13;
    _zz_dataOut_payload_69_5 <= _zz_dataOut_payload_69_4;
    _zz_dataOut_payload_70_8 <= _zz_dataOut_payload_70_7;
    _zz_dataOut_payload_71_5 <= _zz_dataOut_payload_71_4;
    _zz_dataOut_payload_72_26 <= _zz_dataOut_payload_72_25;
    _zz_dataOut_payload_73_5 <= _zz_dataOut_payload_73_4;
    _zz_dataOut_payload_74_8 <= _zz_dataOut_payload_74_7;
    _zz_dataOut_payload_75_5 <= _zz_dataOut_payload_75_4;
    _zz_dataOut_payload_76_14 <= _zz_dataOut_payload_76_13;
    _zz_dataOut_payload_77_5 <= _zz_dataOut_payload_77_4;
    _zz_dataOut_payload_78_8 <= _zz_dataOut_payload_78_7;
    _zz_dataOut_payload_79_5 <= _zz_dataOut_payload_79_4;
    _zz_dataOut_payload_80_50 <= _zz_dataOut_payload_80_49;
    _zz_dataOut_payload_81_5 <= _zz_dataOut_payload_81_4;
    _zz_dataOut_payload_82_8 <= _zz_dataOut_payload_82_7;
    _zz_dataOut_payload_83_5 <= _zz_dataOut_payload_83_4;
    _zz_dataOut_payload_84_14 <= _zz_dataOut_payload_84_13;
    _zz_dataOut_payload_85_5 <= _zz_dataOut_payload_85_4;
    _zz_dataOut_payload_86_8 <= _zz_dataOut_payload_86_7;
    _zz_dataOut_payload_87_5 <= _zz_dataOut_payload_87_4;
    _zz_dataOut_payload_88_26 <= _zz_dataOut_payload_88_25;
    _zz_dataOut_payload_89_5 <= _zz_dataOut_payload_89_4;
    _zz_dataOut_payload_90_8 <= _zz_dataOut_payload_90_7;
    _zz_dataOut_payload_91_5 <= _zz_dataOut_payload_91_4;
    _zz_dataOut_payload_92_14 <= _zz_dataOut_payload_92_13;
    _zz_dataOut_payload_93_5 <= _zz_dataOut_payload_93_4;
    _zz_dataOut_payload_94_8 <= _zz_dataOut_payload_94_7;
    _zz_dataOut_payload_95_5 <= _zz_dataOut_payload_95_4;
    _zz_dataOut_payload_96_98 <= _zz_dataOut_payload_96_97;
    _zz_dataOut_payload_97_5 <= _zz_dataOut_payload_97_4;
    _zz_dataOut_payload_98_8 <= _zz_dataOut_payload_98_7;
    _zz_dataOut_payload_99_5 <= _zz_dataOut_payload_99_4;
    _zz_dataOut_payload_100_14 <= _zz_dataOut_payload_100_13;
    _zz_dataOut_payload_101_5 <= _zz_dataOut_payload_101_4;
    _zz_dataOut_payload_102_8 <= _zz_dataOut_payload_102_7;
    _zz_dataOut_payload_103_5 <= _zz_dataOut_payload_103_4;
    _zz_dataOut_payload_104_26 <= _zz_dataOut_payload_104_25;
    _zz_dataOut_payload_105_5 <= _zz_dataOut_payload_105_4;
    _zz_dataOut_payload_106_8 <= _zz_dataOut_payload_106_7;
    _zz_dataOut_payload_107_5 <= _zz_dataOut_payload_107_4;
    _zz_dataOut_payload_108_14 <= _zz_dataOut_payload_108_13;
    _zz_dataOut_payload_109_5 <= _zz_dataOut_payload_109_4;
    _zz_dataOut_payload_110_8 <= _zz_dataOut_payload_110_7;
    _zz_dataOut_payload_111_5 <= _zz_dataOut_payload_111_4;
    _zz_dataOut_payload_112_50 <= _zz_dataOut_payload_112_49;
    _zz_dataOut_payload_113_5 <= _zz_dataOut_payload_113_4;
    _zz_dataOut_payload_114_8 <= _zz_dataOut_payload_114_7;
    _zz_dataOut_payload_115_5 <= _zz_dataOut_payload_115_4;
    _zz_dataOut_payload_116_14 <= _zz_dataOut_payload_116_13;
    _zz_dataOut_payload_117_5 <= _zz_dataOut_payload_117_4;
    _zz_dataOut_payload_118_8 <= _zz_dataOut_payload_118_7;
    _zz_dataOut_payload_119_5 <= _zz_dataOut_payload_119_4;
    _zz_dataOut_payload_120_26 <= _zz_dataOut_payload_120_25;
    _zz_dataOut_payload_121_5 <= _zz_dataOut_payload_121_4;
    _zz_dataOut_payload_122_8 <= _zz_dataOut_payload_122_7;
    _zz_dataOut_payload_123_5 <= _zz_dataOut_payload_123_4;
    _zz_dataOut_payload_124_14 <= _zz_dataOut_payload_124_13;
    _zz_dataOut_payload_125_5 <= _zz_dataOut_payload_125_4;
    _zz_dataOut_payload_126_8 <= _zz_dataOut_payload_126_7;
    _zz_dataOut_payload_127_5 <= _zz_dataOut_payload_127_4;
    _zz_dataOut_payload_128_381 <= (_zz_dataOut_payload_128_380 ? _zz_dataOut_payload_128_377 : _zz_dataOut_payload_128_379);
    _zz_dataOut_payload_129 <= (_zz_dataOut_payload_128_380 ? _zz_dataOut_payload_128_379 : _zz_dataOut_payload_128_377);
    _zz_dataOut_payload_130_3 <= (_zz_dataOut_payload_130_2 ? _zz_dataOut_payload_130 : _zz_dataOut_payload_130_1);
    _zz_dataOut_payload_131 <= (_zz_dataOut_payload_130_2 ? _zz_dataOut_payload_130_1 : _zz_dataOut_payload_130);
    _zz_dataOut_payload_132_9 <= (_zz_dataOut_payload_132_8 ? _zz_dataOut_payload_132_5 : _zz_dataOut_payload_132_7);
    _zz_dataOut_payload_133 <= (_zz_dataOut_payload_132_8 ? _zz_dataOut_payload_132_7 : _zz_dataOut_payload_132_5);
    _zz_dataOut_payload_134_3 <= (_zz_dataOut_payload_134_2 ? _zz_dataOut_payload_134 : _zz_dataOut_payload_134_1);
    _zz_dataOut_payload_135 <= (_zz_dataOut_payload_134_2 ? _zz_dataOut_payload_134_1 : _zz_dataOut_payload_134);
    _zz_dataOut_payload_128_382 <= _zz_dataOut_payload_128_381;
    _zz_dataOut_payload_129_1 <= _zz_dataOut_payload_129;
    _zz_dataOut_payload_130_4 <= _zz_dataOut_payload_130_3;
    _zz_dataOut_payload_131_1 <= _zz_dataOut_payload_131;
    _zz_dataOut_payload_132_10 <= _zz_dataOut_payload_132_9;
    _zz_dataOut_payload_133_1 <= _zz_dataOut_payload_133;
    _zz_dataOut_payload_134_4 <= _zz_dataOut_payload_134_3;
    _zz_dataOut_payload_135_1 <= _zz_dataOut_payload_135;
    _zz_dataOut_payload_136_21 <= (_zz_dataOut_payload_136_20 ? _zz_dataOut_payload_136_17 : _zz_dataOut_payload_136_19);
    _zz_dataOut_payload_137 <= (_zz_dataOut_payload_136_20 ? _zz_dataOut_payload_136_19 : _zz_dataOut_payload_136_17);
    _zz_dataOut_payload_138_3 <= (_zz_dataOut_payload_138_2 ? _zz_dataOut_payload_138 : _zz_dataOut_payload_138_1);
    _zz_dataOut_payload_139 <= (_zz_dataOut_payload_138_2 ? _zz_dataOut_payload_138_1 : _zz_dataOut_payload_138);
    _zz_dataOut_payload_140_9 <= (_zz_dataOut_payload_140_8 ? _zz_dataOut_payload_140_5 : _zz_dataOut_payload_140_7);
    _zz_dataOut_payload_141 <= (_zz_dataOut_payload_140_8 ? _zz_dataOut_payload_140_7 : _zz_dataOut_payload_140_5);
    _zz_dataOut_payload_142_3 <= (_zz_dataOut_payload_142_2 ? _zz_dataOut_payload_142 : _zz_dataOut_payload_142_1);
    _zz_dataOut_payload_143 <= (_zz_dataOut_payload_142_2 ? _zz_dataOut_payload_142_1 : _zz_dataOut_payload_142);
    _zz_dataOut_payload_136_22 <= _zz_dataOut_payload_136_21;
    _zz_dataOut_payload_137_1 <= _zz_dataOut_payload_137;
    _zz_dataOut_payload_138_4 <= _zz_dataOut_payload_138_3;
    _zz_dataOut_payload_139_1 <= _zz_dataOut_payload_139;
    _zz_dataOut_payload_140_10 <= _zz_dataOut_payload_140_9;
    _zz_dataOut_payload_141_1 <= _zz_dataOut_payload_141;
    _zz_dataOut_payload_142_4 <= _zz_dataOut_payload_142_3;
    _zz_dataOut_payload_143_1 <= _zz_dataOut_payload_143;
    _zz_dataOut_payload_128_383 <= _zz_dataOut_payload_128_382;
    _zz_dataOut_payload_129_2 <= _zz_dataOut_payload_129_1;
    _zz_dataOut_payload_130_5 <= _zz_dataOut_payload_130_4;
    _zz_dataOut_payload_131_2 <= _zz_dataOut_payload_131_1;
    _zz_dataOut_payload_132_11 <= _zz_dataOut_payload_132_10;
    _zz_dataOut_payload_133_2 <= _zz_dataOut_payload_133_1;
    _zz_dataOut_payload_134_5 <= _zz_dataOut_payload_134_4;
    _zz_dataOut_payload_135_2 <= _zz_dataOut_payload_135_1;
    _zz_dataOut_payload_136_23 <= _zz_dataOut_payload_136_22;
    _zz_dataOut_payload_137_2 <= _zz_dataOut_payload_137_1;
    _zz_dataOut_payload_138_5 <= _zz_dataOut_payload_138_4;
    _zz_dataOut_payload_139_2 <= _zz_dataOut_payload_139_1;
    _zz_dataOut_payload_140_11 <= _zz_dataOut_payload_140_10;
    _zz_dataOut_payload_141_2 <= _zz_dataOut_payload_141_1;
    _zz_dataOut_payload_142_5 <= _zz_dataOut_payload_142_4;
    _zz_dataOut_payload_143_2 <= _zz_dataOut_payload_143_1;
    _zz_dataOut_payload_144_45 <= (_zz_dataOut_payload_144_44 ? _zz_dataOut_payload_144_41 : _zz_dataOut_payload_144_43);
    _zz_dataOut_payload_145 <= (_zz_dataOut_payload_144_44 ? _zz_dataOut_payload_144_43 : _zz_dataOut_payload_144_41);
    _zz_dataOut_payload_146_3 <= (_zz_dataOut_payload_146_2 ? _zz_dataOut_payload_146 : _zz_dataOut_payload_146_1);
    _zz_dataOut_payload_147 <= (_zz_dataOut_payload_146_2 ? _zz_dataOut_payload_146_1 : _zz_dataOut_payload_146);
    _zz_dataOut_payload_148_9 <= (_zz_dataOut_payload_148_8 ? _zz_dataOut_payload_148_5 : _zz_dataOut_payload_148_7);
    _zz_dataOut_payload_149 <= (_zz_dataOut_payload_148_8 ? _zz_dataOut_payload_148_7 : _zz_dataOut_payload_148_5);
    _zz_dataOut_payload_150_3 <= (_zz_dataOut_payload_150_2 ? _zz_dataOut_payload_150 : _zz_dataOut_payload_150_1);
    _zz_dataOut_payload_151 <= (_zz_dataOut_payload_150_2 ? _zz_dataOut_payload_150_1 : _zz_dataOut_payload_150);
    _zz_dataOut_payload_144_46 <= _zz_dataOut_payload_144_45;
    _zz_dataOut_payload_145_1 <= _zz_dataOut_payload_145;
    _zz_dataOut_payload_146_4 <= _zz_dataOut_payload_146_3;
    _zz_dataOut_payload_147_1 <= _zz_dataOut_payload_147;
    _zz_dataOut_payload_148_10 <= _zz_dataOut_payload_148_9;
    _zz_dataOut_payload_149_1 <= _zz_dataOut_payload_149;
    _zz_dataOut_payload_150_4 <= _zz_dataOut_payload_150_3;
    _zz_dataOut_payload_151_1 <= _zz_dataOut_payload_151;
    _zz_dataOut_payload_152_21 <= (_zz_dataOut_payload_152_20 ? _zz_dataOut_payload_152_17 : _zz_dataOut_payload_152_19);
    _zz_dataOut_payload_153 <= (_zz_dataOut_payload_152_20 ? _zz_dataOut_payload_152_19 : _zz_dataOut_payload_152_17);
    _zz_dataOut_payload_154_3 <= (_zz_dataOut_payload_154_2 ? _zz_dataOut_payload_154 : _zz_dataOut_payload_154_1);
    _zz_dataOut_payload_155 <= (_zz_dataOut_payload_154_2 ? _zz_dataOut_payload_154_1 : _zz_dataOut_payload_154);
    _zz_dataOut_payload_156_9 <= (_zz_dataOut_payload_156_8 ? _zz_dataOut_payload_156_5 : _zz_dataOut_payload_156_7);
    _zz_dataOut_payload_157 <= (_zz_dataOut_payload_156_8 ? _zz_dataOut_payload_156_7 : _zz_dataOut_payload_156_5);
    _zz_dataOut_payload_158_3 <= (_zz_dataOut_payload_158_2 ? _zz_dataOut_payload_158 : _zz_dataOut_payload_158_1);
    _zz_dataOut_payload_159 <= (_zz_dataOut_payload_158_2 ? _zz_dataOut_payload_158_1 : _zz_dataOut_payload_158);
    _zz_dataOut_payload_152_22 <= _zz_dataOut_payload_152_21;
    _zz_dataOut_payload_153_1 <= _zz_dataOut_payload_153;
    _zz_dataOut_payload_154_4 <= _zz_dataOut_payload_154_3;
    _zz_dataOut_payload_155_1 <= _zz_dataOut_payload_155;
    _zz_dataOut_payload_156_10 <= _zz_dataOut_payload_156_9;
    _zz_dataOut_payload_157_1 <= _zz_dataOut_payload_157;
    _zz_dataOut_payload_158_4 <= _zz_dataOut_payload_158_3;
    _zz_dataOut_payload_159_1 <= _zz_dataOut_payload_159;
    _zz_dataOut_payload_144_47 <= _zz_dataOut_payload_144_46;
    _zz_dataOut_payload_145_2 <= _zz_dataOut_payload_145_1;
    _zz_dataOut_payload_146_5 <= _zz_dataOut_payload_146_4;
    _zz_dataOut_payload_147_2 <= _zz_dataOut_payload_147_1;
    _zz_dataOut_payload_148_11 <= _zz_dataOut_payload_148_10;
    _zz_dataOut_payload_149_2 <= _zz_dataOut_payload_149_1;
    _zz_dataOut_payload_150_5 <= _zz_dataOut_payload_150_4;
    _zz_dataOut_payload_151_2 <= _zz_dataOut_payload_151_1;
    _zz_dataOut_payload_152_23 <= _zz_dataOut_payload_152_22;
    _zz_dataOut_payload_153_2 <= _zz_dataOut_payload_153_1;
    _zz_dataOut_payload_154_5 <= _zz_dataOut_payload_154_4;
    _zz_dataOut_payload_155_2 <= _zz_dataOut_payload_155_1;
    _zz_dataOut_payload_156_11 <= _zz_dataOut_payload_156_10;
    _zz_dataOut_payload_157_2 <= _zz_dataOut_payload_157_1;
    _zz_dataOut_payload_158_5 <= _zz_dataOut_payload_158_4;
    _zz_dataOut_payload_159_2 <= _zz_dataOut_payload_159_1;
    _zz_dataOut_payload_128_384 <= _zz_dataOut_payload_128_383;
    _zz_dataOut_payload_129_3 <= _zz_dataOut_payload_129_2;
    _zz_dataOut_payload_130_6 <= _zz_dataOut_payload_130_5;
    _zz_dataOut_payload_131_3 <= _zz_dataOut_payload_131_2;
    _zz_dataOut_payload_132_12 <= _zz_dataOut_payload_132_11;
    _zz_dataOut_payload_133_3 <= _zz_dataOut_payload_133_2;
    _zz_dataOut_payload_134_6 <= _zz_dataOut_payload_134_5;
    _zz_dataOut_payload_135_3 <= _zz_dataOut_payload_135_2;
    _zz_dataOut_payload_136_24 <= _zz_dataOut_payload_136_23;
    _zz_dataOut_payload_137_3 <= _zz_dataOut_payload_137_2;
    _zz_dataOut_payload_138_6 <= _zz_dataOut_payload_138_5;
    _zz_dataOut_payload_139_3 <= _zz_dataOut_payload_139_2;
    _zz_dataOut_payload_140_12 <= _zz_dataOut_payload_140_11;
    _zz_dataOut_payload_141_3 <= _zz_dataOut_payload_141_2;
    _zz_dataOut_payload_142_6 <= _zz_dataOut_payload_142_5;
    _zz_dataOut_payload_143_3 <= _zz_dataOut_payload_143_2;
    _zz_dataOut_payload_144_48 <= _zz_dataOut_payload_144_47;
    _zz_dataOut_payload_145_3 <= _zz_dataOut_payload_145_2;
    _zz_dataOut_payload_146_6 <= _zz_dataOut_payload_146_5;
    _zz_dataOut_payload_147_3 <= _zz_dataOut_payload_147_2;
    _zz_dataOut_payload_148_12 <= _zz_dataOut_payload_148_11;
    _zz_dataOut_payload_149_3 <= _zz_dataOut_payload_149_2;
    _zz_dataOut_payload_150_6 <= _zz_dataOut_payload_150_5;
    _zz_dataOut_payload_151_3 <= _zz_dataOut_payload_151_2;
    _zz_dataOut_payload_152_24 <= _zz_dataOut_payload_152_23;
    _zz_dataOut_payload_153_3 <= _zz_dataOut_payload_153_2;
    _zz_dataOut_payload_154_6 <= _zz_dataOut_payload_154_5;
    _zz_dataOut_payload_155_3 <= _zz_dataOut_payload_155_2;
    _zz_dataOut_payload_156_12 <= _zz_dataOut_payload_156_11;
    _zz_dataOut_payload_157_3 <= _zz_dataOut_payload_157_2;
    _zz_dataOut_payload_158_6 <= _zz_dataOut_payload_158_5;
    _zz_dataOut_payload_159_3 <= _zz_dataOut_payload_159_2;
    _zz_dataOut_payload_160_93 <= (_zz_dataOut_payload_160_92 ? _zz_dataOut_payload_160_89 : _zz_dataOut_payload_160_91);
    _zz_dataOut_payload_161 <= (_zz_dataOut_payload_160_92 ? _zz_dataOut_payload_160_91 : _zz_dataOut_payload_160_89);
    _zz_dataOut_payload_162_3 <= (_zz_dataOut_payload_162_2 ? _zz_dataOut_payload_162 : _zz_dataOut_payload_162_1);
    _zz_dataOut_payload_163 <= (_zz_dataOut_payload_162_2 ? _zz_dataOut_payload_162_1 : _zz_dataOut_payload_162);
    _zz_dataOut_payload_164_9 <= (_zz_dataOut_payload_164_8 ? _zz_dataOut_payload_164_5 : _zz_dataOut_payload_164_7);
    _zz_dataOut_payload_165 <= (_zz_dataOut_payload_164_8 ? _zz_dataOut_payload_164_7 : _zz_dataOut_payload_164_5);
    _zz_dataOut_payload_166_3 <= (_zz_dataOut_payload_166_2 ? _zz_dataOut_payload_166 : _zz_dataOut_payload_166_1);
    _zz_dataOut_payload_167 <= (_zz_dataOut_payload_166_2 ? _zz_dataOut_payload_166_1 : _zz_dataOut_payload_166);
    _zz_dataOut_payload_160_94 <= _zz_dataOut_payload_160_93;
    _zz_dataOut_payload_161_1 <= _zz_dataOut_payload_161;
    _zz_dataOut_payload_162_4 <= _zz_dataOut_payload_162_3;
    _zz_dataOut_payload_163_1 <= _zz_dataOut_payload_163;
    _zz_dataOut_payload_164_10 <= _zz_dataOut_payload_164_9;
    _zz_dataOut_payload_165_1 <= _zz_dataOut_payload_165;
    _zz_dataOut_payload_166_4 <= _zz_dataOut_payload_166_3;
    _zz_dataOut_payload_167_1 <= _zz_dataOut_payload_167;
    _zz_dataOut_payload_168_21 <= (_zz_dataOut_payload_168_20 ? _zz_dataOut_payload_168_17 : _zz_dataOut_payload_168_19);
    _zz_dataOut_payload_169 <= (_zz_dataOut_payload_168_20 ? _zz_dataOut_payload_168_19 : _zz_dataOut_payload_168_17);
    _zz_dataOut_payload_170_3 <= (_zz_dataOut_payload_170_2 ? _zz_dataOut_payload_170 : _zz_dataOut_payload_170_1);
    _zz_dataOut_payload_171 <= (_zz_dataOut_payload_170_2 ? _zz_dataOut_payload_170_1 : _zz_dataOut_payload_170);
    _zz_dataOut_payload_172_9 <= (_zz_dataOut_payload_172_8 ? _zz_dataOut_payload_172_5 : _zz_dataOut_payload_172_7);
    _zz_dataOut_payload_173 <= (_zz_dataOut_payload_172_8 ? _zz_dataOut_payload_172_7 : _zz_dataOut_payload_172_5);
    _zz_dataOut_payload_174_3 <= (_zz_dataOut_payload_174_2 ? _zz_dataOut_payload_174 : _zz_dataOut_payload_174_1);
    _zz_dataOut_payload_175 <= (_zz_dataOut_payload_174_2 ? _zz_dataOut_payload_174_1 : _zz_dataOut_payload_174);
    _zz_dataOut_payload_168_22 <= _zz_dataOut_payload_168_21;
    _zz_dataOut_payload_169_1 <= _zz_dataOut_payload_169;
    _zz_dataOut_payload_170_4 <= _zz_dataOut_payload_170_3;
    _zz_dataOut_payload_171_1 <= _zz_dataOut_payload_171;
    _zz_dataOut_payload_172_10 <= _zz_dataOut_payload_172_9;
    _zz_dataOut_payload_173_1 <= _zz_dataOut_payload_173;
    _zz_dataOut_payload_174_4 <= _zz_dataOut_payload_174_3;
    _zz_dataOut_payload_175_1 <= _zz_dataOut_payload_175;
    _zz_dataOut_payload_160_95 <= _zz_dataOut_payload_160_94;
    _zz_dataOut_payload_161_2 <= _zz_dataOut_payload_161_1;
    _zz_dataOut_payload_162_5 <= _zz_dataOut_payload_162_4;
    _zz_dataOut_payload_163_2 <= _zz_dataOut_payload_163_1;
    _zz_dataOut_payload_164_11 <= _zz_dataOut_payload_164_10;
    _zz_dataOut_payload_165_2 <= _zz_dataOut_payload_165_1;
    _zz_dataOut_payload_166_5 <= _zz_dataOut_payload_166_4;
    _zz_dataOut_payload_167_2 <= _zz_dataOut_payload_167_1;
    _zz_dataOut_payload_168_23 <= _zz_dataOut_payload_168_22;
    _zz_dataOut_payload_169_2 <= _zz_dataOut_payload_169_1;
    _zz_dataOut_payload_170_5 <= _zz_dataOut_payload_170_4;
    _zz_dataOut_payload_171_2 <= _zz_dataOut_payload_171_1;
    _zz_dataOut_payload_172_11 <= _zz_dataOut_payload_172_10;
    _zz_dataOut_payload_173_2 <= _zz_dataOut_payload_173_1;
    _zz_dataOut_payload_174_5 <= _zz_dataOut_payload_174_4;
    _zz_dataOut_payload_175_2 <= _zz_dataOut_payload_175_1;
    _zz_dataOut_payload_176_45 <= (_zz_dataOut_payload_176_44 ? _zz_dataOut_payload_176_41 : _zz_dataOut_payload_176_43);
    _zz_dataOut_payload_177 <= (_zz_dataOut_payload_176_44 ? _zz_dataOut_payload_176_43 : _zz_dataOut_payload_176_41);
    _zz_dataOut_payload_178_3 <= (_zz_dataOut_payload_178_2 ? _zz_dataOut_payload_178 : _zz_dataOut_payload_178_1);
    _zz_dataOut_payload_179 <= (_zz_dataOut_payload_178_2 ? _zz_dataOut_payload_178_1 : _zz_dataOut_payload_178);
    _zz_dataOut_payload_180_9 <= (_zz_dataOut_payload_180_8 ? _zz_dataOut_payload_180_5 : _zz_dataOut_payload_180_7);
    _zz_dataOut_payload_181 <= (_zz_dataOut_payload_180_8 ? _zz_dataOut_payload_180_7 : _zz_dataOut_payload_180_5);
    _zz_dataOut_payload_182_3 <= (_zz_dataOut_payload_182_2 ? _zz_dataOut_payload_182 : _zz_dataOut_payload_182_1);
    _zz_dataOut_payload_183 <= (_zz_dataOut_payload_182_2 ? _zz_dataOut_payload_182_1 : _zz_dataOut_payload_182);
    _zz_dataOut_payload_176_46 <= _zz_dataOut_payload_176_45;
    _zz_dataOut_payload_177_1 <= _zz_dataOut_payload_177;
    _zz_dataOut_payload_178_4 <= _zz_dataOut_payload_178_3;
    _zz_dataOut_payload_179_1 <= _zz_dataOut_payload_179;
    _zz_dataOut_payload_180_10 <= _zz_dataOut_payload_180_9;
    _zz_dataOut_payload_181_1 <= _zz_dataOut_payload_181;
    _zz_dataOut_payload_182_4 <= _zz_dataOut_payload_182_3;
    _zz_dataOut_payload_183_1 <= _zz_dataOut_payload_183;
    _zz_dataOut_payload_184_21 <= (_zz_dataOut_payload_184_20 ? _zz_dataOut_payload_184_17 : _zz_dataOut_payload_184_19);
    _zz_dataOut_payload_185 <= (_zz_dataOut_payload_184_20 ? _zz_dataOut_payload_184_19 : _zz_dataOut_payload_184_17);
    _zz_dataOut_payload_186_3 <= (_zz_dataOut_payload_186_2 ? _zz_dataOut_payload_186 : _zz_dataOut_payload_186_1);
    _zz_dataOut_payload_187 <= (_zz_dataOut_payload_186_2 ? _zz_dataOut_payload_186_1 : _zz_dataOut_payload_186);
    _zz_dataOut_payload_188_9 <= (_zz_dataOut_payload_188_8 ? _zz_dataOut_payload_188_5 : _zz_dataOut_payload_188_7);
    _zz_dataOut_payload_189 <= (_zz_dataOut_payload_188_8 ? _zz_dataOut_payload_188_7 : _zz_dataOut_payload_188_5);
    _zz_dataOut_payload_190_3 <= (_zz_dataOut_payload_190_2 ? _zz_dataOut_payload_190 : _zz_dataOut_payload_190_1);
    _zz_dataOut_payload_191 <= (_zz_dataOut_payload_190_2 ? _zz_dataOut_payload_190_1 : _zz_dataOut_payload_190);
    _zz_dataOut_payload_184_22 <= _zz_dataOut_payload_184_21;
    _zz_dataOut_payload_185_1 <= _zz_dataOut_payload_185;
    _zz_dataOut_payload_186_4 <= _zz_dataOut_payload_186_3;
    _zz_dataOut_payload_187_1 <= _zz_dataOut_payload_187;
    _zz_dataOut_payload_188_10 <= _zz_dataOut_payload_188_9;
    _zz_dataOut_payload_189_1 <= _zz_dataOut_payload_189;
    _zz_dataOut_payload_190_4 <= _zz_dataOut_payload_190_3;
    _zz_dataOut_payload_191_1 <= _zz_dataOut_payload_191;
    _zz_dataOut_payload_176_47 <= _zz_dataOut_payload_176_46;
    _zz_dataOut_payload_177_2 <= _zz_dataOut_payload_177_1;
    _zz_dataOut_payload_178_5 <= _zz_dataOut_payload_178_4;
    _zz_dataOut_payload_179_2 <= _zz_dataOut_payload_179_1;
    _zz_dataOut_payload_180_11 <= _zz_dataOut_payload_180_10;
    _zz_dataOut_payload_181_2 <= _zz_dataOut_payload_181_1;
    _zz_dataOut_payload_182_5 <= _zz_dataOut_payload_182_4;
    _zz_dataOut_payload_183_2 <= _zz_dataOut_payload_183_1;
    _zz_dataOut_payload_184_23 <= _zz_dataOut_payload_184_22;
    _zz_dataOut_payload_185_2 <= _zz_dataOut_payload_185_1;
    _zz_dataOut_payload_186_5 <= _zz_dataOut_payload_186_4;
    _zz_dataOut_payload_187_2 <= _zz_dataOut_payload_187_1;
    _zz_dataOut_payload_188_11 <= _zz_dataOut_payload_188_10;
    _zz_dataOut_payload_189_2 <= _zz_dataOut_payload_189_1;
    _zz_dataOut_payload_190_5 <= _zz_dataOut_payload_190_4;
    _zz_dataOut_payload_191_2 <= _zz_dataOut_payload_191_1;
    _zz_dataOut_payload_160_96 <= _zz_dataOut_payload_160_95;
    _zz_dataOut_payload_161_3 <= _zz_dataOut_payload_161_2;
    _zz_dataOut_payload_162_6 <= _zz_dataOut_payload_162_5;
    _zz_dataOut_payload_163_3 <= _zz_dataOut_payload_163_2;
    _zz_dataOut_payload_164_12 <= _zz_dataOut_payload_164_11;
    _zz_dataOut_payload_165_3 <= _zz_dataOut_payload_165_2;
    _zz_dataOut_payload_166_6 <= _zz_dataOut_payload_166_5;
    _zz_dataOut_payload_167_3 <= _zz_dataOut_payload_167_2;
    _zz_dataOut_payload_168_24 <= _zz_dataOut_payload_168_23;
    _zz_dataOut_payload_169_3 <= _zz_dataOut_payload_169_2;
    _zz_dataOut_payload_170_6 <= _zz_dataOut_payload_170_5;
    _zz_dataOut_payload_171_3 <= _zz_dataOut_payload_171_2;
    _zz_dataOut_payload_172_12 <= _zz_dataOut_payload_172_11;
    _zz_dataOut_payload_173_3 <= _zz_dataOut_payload_173_2;
    _zz_dataOut_payload_174_6 <= _zz_dataOut_payload_174_5;
    _zz_dataOut_payload_175_3 <= _zz_dataOut_payload_175_2;
    _zz_dataOut_payload_176_48 <= _zz_dataOut_payload_176_47;
    _zz_dataOut_payload_177_3 <= _zz_dataOut_payload_177_2;
    _zz_dataOut_payload_178_6 <= _zz_dataOut_payload_178_5;
    _zz_dataOut_payload_179_3 <= _zz_dataOut_payload_179_2;
    _zz_dataOut_payload_180_12 <= _zz_dataOut_payload_180_11;
    _zz_dataOut_payload_181_3 <= _zz_dataOut_payload_181_2;
    _zz_dataOut_payload_182_6 <= _zz_dataOut_payload_182_5;
    _zz_dataOut_payload_183_3 <= _zz_dataOut_payload_183_2;
    _zz_dataOut_payload_184_24 <= _zz_dataOut_payload_184_23;
    _zz_dataOut_payload_185_3 <= _zz_dataOut_payload_185_2;
    _zz_dataOut_payload_186_6 <= _zz_dataOut_payload_186_5;
    _zz_dataOut_payload_187_3 <= _zz_dataOut_payload_187_2;
    _zz_dataOut_payload_188_12 <= _zz_dataOut_payload_188_11;
    _zz_dataOut_payload_189_3 <= _zz_dataOut_payload_189_2;
    _zz_dataOut_payload_190_6 <= _zz_dataOut_payload_190_5;
    _zz_dataOut_payload_191_3 <= _zz_dataOut_payload_191_2;
    _zz_dataOut_payload_128_385 <= _zz_dataOut_payload_128_384;
    _zz_dataOut_payload_129_4 <= _zz_dataOut_payload_129_3;
    _zz_dataOut_payload_130_7 <= _zz_dataOut_payload_130_6;
    _zz_dataOut_payload_131_4 <= _zz_dataOut_payload_131_3;
    _zz_dataOut_payload_132_13 <= _zz_dataOut_payload_132_12;
    _zz_dataOut_payload_133_4 <= _zz_dataOut_payload_133_3;
    _zz_dataOut_payload_134_7 <= _zz_dataOut_payload_134_6;
    _zz_dataOut_payload_135_4 <= _zz_dataOut_payload_135_3;
    _zz_dataOut_payload_136_25 <= _zz_dataOut_payload_136_24;
    _zz_dataOut_payload_137_4 <= _zz_dataOut_payload_137_3;
    _zz_dataOut_payload_138_7 <= _zz_dataOut_payload_138_6;
    _zz_dataOut_payload_139_4 <= _zz_dataOut_payload_139_3;
    _zz_dataOut_payload_140_13 <= _zz_dataOut_payload_140_12;
    _zz_dataOut_payload_141_4 <= _zz_dataOut_payload_141_3;
    _zz_dataOut_payload_142_7 <= _zz_dataOut_payload_142_6;
    _zz_dataOut_payload_143_4 <= _zz_dataOut_payload_143_3;
    _zz_dataOut_payload_144_49 <= _zz_dataOut_payload_144_48;
    _zz_dataOut_payload_145_4 <= _zz_dataOut_payload_145_3;
    _zz_dataOut_payload_146_7 <= _zz_dataOut_payload_146_6;
    _zz_dataOut_payload_147_4 <= _zz_dataOut_payload_147_3;
    _zz_dataOut_payload_148_13 <= _zz_dataOut_payload_148_12;
    _zz_dataOut_payload_149_4 <= _zz_dataOut_payload_149_3;
    _zz_dataOut_payload_150_7 <= _zz_dataOut_payload_150_6;
    _zz_dataOut_payload_151_4 <= _zz_dataOut_payload_151_3;
    _zz_dataOut_payload_152_25 <= _zz_dataOut_payload_152_24;
    _zz_dataOut_payload_153_4 <= _zz_dataOut_payload_153_3;
    _zz_dataOut_payload_154_7 <= _zz_dataOut_payload_154_6;
    _zz_dataOut_payload_155_4 <= _zz_dataOut_payload_155_3;
    _zz_dataOut_payload_156_13 <= _zz_dataOut_payload_156_12;
    _zz_dataOut_payload_157_4 <= _zz_dataOut_payload_157_3;
    _zz_dataOut_payload_158_7 <= _zz_dataOut_payload_158_6;
    _zz_dataOut_payload_159_4 <= _zz_dataOut_payload_159_3;
    _zz_dataOut_payload_160_97 <= _zz_dataOut_payload_160_96;
    _zz_dataOut_payload_161_4 <= _zz_dataOut_payload_161_3;
    _zz_dataOut_payload_162_7 <= _zz_dataOut_payload_162_6;
    _zz_dataOut_payload_163_4 <= _zz_dataOut_payload_163_3;
    _zz_dataOut_payload_164_13 <= _zz_dataOut_payload_164_12;
    _zz_dataOut_payload_165_4 <= _zz_dataOut_payload_165_3;
    _zz_dataOut_payload_166_7 <= _zz_dataOut_payload_166_6;
    _zz_dataOut_payload_167_4 <= _zz_dataOut_payload_167_3;
    _zz_dataOut_payload_168_25 <= _zz_dataOut_payload_168_24;
    _zz_dataOut_payload_169_4 <= _zz_dataOut_payload_169_3;
    _zz_dataOut_payload_170_7 <= _zz_dataOut_payload_170_6;
    _zz_dataOut_payload_171_4 <= _zz_dataOut_payload_171_3;
    _zz_dataOut_payload_172_13 <= _zz_dataOut_payload_172_12;
    _zz_dataOut_payload_173_4 <= _zz_dataOut_payload_173_3;
    _zz_dataOut_payload_174_7 <= _zz_dataOut_payload_174_6;
    _zz_dataOut_payload_175_4 <= _zz_dataOut_payload_175_3;
    _zz_dataOut_payload_176_49 <= _zz_dataOut_payload_176_48;
    _zz_dataOut_payload_177_4 <= _zz_dataOut_payload_177_3;
    _zz_dataOut_payload_178_7 <= _zz_dataOut_payload_178_6;
    _zz_dataOut_payload_179_4 <= _zz_dataOut_payload_179_3;
    _zz_dataOut_payload_180_13 <= _zz_dataOut_payload_180_12;
    _zz_dataOut_payload_181_4 <= _zz_dataOut_payload_181_3;
    _zz_dataOut_payload_182_7 <= _zz_dataOut_payload_182_6;
    _zz_dataOut_payload_183_4 <= _zz_dataOut_payload_183_3;
    _zz_dataOut_payload_184_25 <= _zz_dataOut_payload_184_24;
    _zz_dataOut_payload_185_4 <= _zz_dataOut_payload_185_3;
    _zz_dataOut_payload_186_7 <= _zz_dataOut_payload_186_6;
    _zz_dataOut_payload_187_4 <= _zz_dataOut_payload_187_3;
    _zz_dataOut_payload_188_13 <= _zz_dataOut_payload_188_12;
    _zz_dataOut_payload_189_4 <= _zz_dataOut_payload_189_3;
    _zz_dataOut_payload_190_7 <= _zz_dataOut_payload_190_6;
    _zz_dataOut_payload_191_4 <= _zz_dataOut_payload_191_3;
    _zz_dataOut_payload_192_189 <= (_zz_dataOut_payload_192_188 ? _zz_dataOut_payload_192_185 : _zz_dataOut_payload_192_187);
    _zz_dataOut_payload_193 <= (_zz_dataOut_payload_192_188 ? _zz_dataOut_payload_192_187 : _zz_dataOut_payload_192_185);
    _zz_dataOut_payload_194_3 <= (_zz_dataOut_payload_194_2 ? _zz_dataOut_payload_194 : _zz_dataOut_payload_194_1);
    _zz_dataOut_payload_195 <= (_zz_dataOut_payload_194_2 ? _zz_dataOut_payload_194_1 : _zz_dataOut_payload_194);
    _zz_dataOut_payload_196_9 <= (_zz_dataOut_payload_196_8 ? _zz_dataOut_payload_196_5 : _zz_dataOut_payload_196_7);
    _zz_dataOut_payload_197 <= (_zz_dataOut_payload_196_8 ? _zz_dataOut_payload_196_7 : _zz_dataOut_payload_196_5);
    _zz_dataOut_payload_198_3 <= (_zz_dataOut_payload_198_2 ? _zz_dataOut_payload_198 : _zz_dataOut_payload_198_1);
    _zz_dataOut_payload_199 <= (_zz_dataOut_payload_198_2 ? _zz_dataOut_payload_198_1 : _zz_dataOut_payload_198);
    _zz_dataOut_payload_192_190 <= _zz_dataOut_payload_192_189;
    _zz_dataOut_payload_193_1 <= _zz_dataOut_payload_193;
    _zz_dataOut_payload_194_4 <= _zz_dataOut_payload_194_3;
    _zz_dataOut_payload_195_1 <= _zz_dataOut_payload_195;
    _zz_dataOut_payload_196_10 <= _zz_dataOut_payload_196_9;
    _zz_dataOut_payload_197_1 <= _zz_dataOut_payload_197;
    _zz_dataOut_payload_198_4 <= _zz_dataOut_payload_198_3;
    _zz_dataOut_payload_199_1 <= _zz_dataOut_payload_199;
    _zz_dataOut_payload_200_21 <= (_zz_dataOut_payload_200_20 ? _zz_dataOut_payload_200_17 : _zz_dataOut_payload_200_19);
    _zz_dataOut_payload_201 <= (_zz_dataOut_payload_200_20 ? _zz_dataOut_payload_200_19 : _zz_dataOut_payload_200_17);
    _zz_dataOut_payload_202_3 <= (_zz_dataOut_payload_202_2 ? _zz_dataOut_payload_202 : _zz_dataOut_payload_202_1);
    _zz_dataOut_payload_203 <= (_zz_dataOut_payload_202_2 ? _zz_dataOut_payload_202_1 : _zz_dataOut_payload_202);
    _zz_dataOut_payload_204_9 <= (_zz_dataOut_payload_204_8 ? _zz_dataOut_payload_204_5 : _zz_dataOut_payload_204_7);
    _zz_dataOut_payload_205 <= (_zz_dataOut_payload_204_8 ? _zz_dataOut_payload_204_7 : _zz_dataOut_payload_204_5);
    _zz_dataOut_payload_206_3 <= (_zz_dataOut_payload_206_2 ? _zz_dataOut_payload_206 : _zz_dataOut_payload_206_1);
    _zz_dataOut_payload_207 <= (_zz_dataOut_payload_206_2 ? _zz_dataOut_payload_206_1 : _zz_dataOut_payload_206);
    _zz_dataOut_payload_200_22 <= _zz_dataOut_payload_200_21;
    _zz_dataOut_payload_201_1 <= _zz_dataOut_payload_201;
    _zz_dataOut_payload_202_4 <= _zz_dataOut_payload_202_3;
    _zz_dataOut_payload_203_1 <= _zz_dataOut_payload_203;
    _zz_dataOut_payload_204_10 <= _zz_dataOut_payload_204_9;
    _zz_dataOut_payload_205_1 <= _zz_dataOut_payload_205;
    _zz_dataOut_payload_206_4 <= _zz_dataOut_payload_206_3;
    _zz_dataOut_payload_207_1 <= _zz_dataOut_payload_207;
    _zz_dataOut_payload_192_191 <= _zz_dataOut_payload_192_190;
    _zz_dataOut_payload_193_2 <= _zz_dataOut_payload_193_1;
    _zz_dataOut_payload_194_5 <= _zz_dataOut_payload_194_4;
    _zz_dataOut_payload_195_2 <= _zz_dataOut_payload_195_1;
    _zz_dataOut_payload_196_11 <= _zz_dataOut_payload_196_10;
    _zz_dataOut_payload_197_2 <= _zz_dataOut_payload_197_1;
    _zz_dataOut_payload_198_5 <= _zz_dataOut_payload_198_4;
    _zz_dataOut_payload_199_2 <= _zz_dataOut_payload_199_1;
    _zz_dataOut_payload_200_23 <= _zz_dataOut_payload_200_22;
    _zz_dataOut_payload_201_2 <= _zz_dataOut_payload_201_1;
    _zz_dataOut_payload_202_5 <= _zz_dataOut_payload_202_4;
    _zz_dataOut_payload_203_2 <= _zz_dataOut_payload_203_1;
    _zz_dataOut_payload_204_11 <= _zz_dataOut_payload_204_10;
    _zz_dataOut_payload_205_2 <= _zz_dataOut_payload_205_1;
    _zz_dataOut_payload_206_5 <= _zz_dataOut_payload_206_4;
    _zz_dataOut_payload_207_2 <= _zz_dataOut_payload_207_1;
    _zz_dataOut_payload_208_45 <= (_zz_dataOut_payload_208_44 ? _zz_dataOut_payload_208_41 : _zz_dataOut_payload_208_43);
    _zz_dataOut_payload_209 <= (_zz_dataOut_payload_208_44 ? _zz_dataOut_payload_208_43 : _zz_dataOut_payload_208_41);
    _zz_dataOut_payload_210_3 <= (_zz_dataOut_payload_210_2 ? _zz_dataOut_payload_210 : _zz_dataOut_payload_210_1);
    _zz_dataOut_payload_211 <= (_zz_dataOut_payload_210_2 ? _zz_dataOut_payload_210_1 : _zz_dataOut_payload_210);
    _zz_dataOut_payload_212_9 <= (_zz_dataOut_payload_212_8 ? _zz_dataOut_payload_212_5 : _zz_dataOut_payload_212_7);
    _zz_dataOut_payload_213 <= (_zz_dataOut_payload_212_8 ? _zz_dataOut_payload_212_7 : _zz_dataOut_payload_212_5);
    _zz_dataOut_payload_214_3 <= (_zz_dataOut_payload_214_2 ? _zz_dataOut_payload_214 : _zz_dataOut_payload_214_1);
    _zz_dataOut_payload_215 <= (_zz_dataOut_payload_214_2 ? _zz_dataOut_payload_214_1 : _zz_dataOut_payload_214);
    _zz_dataOut_payload_208_46 <= _zz_dataOut_payload_208_45;
    _zz_dataOut_payload_209_1 <= _zz_dataOut_payload_209;
    _zz_dataOut_payload_210_4 <= _zz_dataOut_payload_210_3;
    _zz_dataOut_payload_211_1 <= _zz_dataOut_payload_211;
    _zz_dataOut_payload_212_10 <= _zz_dataOut_payload_212_9;
    _zz_dataOut_payload_213_1 <= _zz_dataOut_payload_213;
    _zz_dataOut_payload_214_4 <= _zz_dataOut_payload_214_3;
    _zz_dataOut_payload_215_1 <= _zz_dataOut_payload_215;
    _zz_dataOut_payload_216_21 <= (_zz_dataOut_payload_216_20 ? _zz_dataOut_payload_216_17 : _zz_dataOut_payload_216_19);
    _zz_dataOut_payload_217 <= (_zz_dataOut_payload_216_20 ? _zz_dataOut_payload_216_19 : _zz_dataOut_payload_216_17);
    _zz_dataOut_payload_218_3 <= (_zz_dataOut_payload_218_2 ? _zz_dataOut_payload_218 : _zz_dataOut_payload_218_1);
    _zz_dataOut_payload_219 <= (_zz_dataOut_payload_218_2 ? _zz_dataOut_payload_218_1 : _zz_dataOut_payload_218);
    _zz_dataOut_payload_220_9 <= (_zz_dataOut_payload_220_8 ? _zz_dataOut_payload_220_5 : _zz_dataOut_payload_220_7);
    _zz_dataOut_payload_221 <= (_zz_dataOut_payload_220_8 ? _zz_dataOut_payload_220_7 : _zz_dataOut_payload_220_5);
    _zz_dataOut_payload_222_3 <= (_zz_dataOut_payload_222_2 ? _zz_dataOut_payload_222 : _zz_dataOut_payload_222_1);
    _zz_dataOut_payload_223 <= (_zz_dataOut_payload_222_2 ? _zz_dataOut_payload_222_1 : _zz_dataOut_payload_222);
    _zz_dataOut_payload_216_22 <= _zz_dataOut_payload_216_21;
    _zz_dataOut_payload_217_1 <= _zz_dataOut_payload_217;
    _zz_dataOut_payload_218_4 <= _zz_dataOut_payload_218_3;
    _zz_dataOut_payload_219_1 <= _zz_dataOut_payload_219;
    _zz_dataOut_payload_220_10 <= _zz_dataOut_payload_220_9;
    _zz_dataOut_payload_221_1 <= _zz_dataOut_payload_221;
    _zz_dataOut_payload_222_4 <= _zz_dataOut_payload_222_3;
    _zz_dataOut_payload_223_1 <= _zz_dataOut_payload_223;
    _zz_dataOut_payload_208_47 <= _zz_dataOut_payload_208_46;
    _zz_dataOut_payload_209_2 <= _zz_dataOut_payload_209_1;
    _zz_dataOut_payload_210_5 <= _zz_dataOut_payload_210_4;
    _zz_dataOut_payload_211_2 <= _zz_dataOut_payload_211_1;
    _zz_dataOut_payload_212_11 <= _zz_dataOut_payload_212_10;
    _zz_dataOut_payload_213_2 <= _zz_dataOut_payload_213_1;
    _zz_dataOut_payload_214_5 <= _zz_dataOut_payload_214_4;
    _zz_dataOut_payload_215_2 <= _zz_dataOut_payload_215_1;
    _zz_dataOut_payload_216_23 <= _zz_dataOut_payload_216_22;
    _zz_dataOut_payload_217_2 <= _zz_dataOut_payload_217_1;
    _zz_dataOut_payload_218_5 <= _zz_dataOut_payload_218_4;
    _zz_dataOut_payload_219_2 <= _zz_dataOut_payload_219_1;
    _zz_dataOut_payload_220_11 <= _zz_dataOut_payload_220_10;
    _zz_dataOut_payload_221_2 <= _zz_dataOut_payload_221_1;
    _zz_dataOut_payload_222_5 <= _zz_dataOut_payload_222_4;
    _zz_dataOut_payload_223_2 <= _zz_dataOut_payload_223_1;
    _zz_dataOut_payload_192_192 <= _zz_dataOut_payload_192_191;
    _zz_dataOut_payload_193_3 <= _zz_dataOut_payload_193_2;
    _zz_dataOut_payload_194_6 <= _zz_dataOut_payload_194_5;
    _zz_dataOut_payload_195_3 <= _zz_dataOut_payload_195_2;
    _zz_dataOut_payload_196_12 <= _zz_dataOut_payload_196_11;
    _zz_dataOut_payload_197_3 <= _zz_dataOut_payload_197_2;
    _zz_dataOut_payload_198_6 <= _zz_dataOut_payload_198_5;
    _zz_dataOut_payload_199_3 <= _zz_dataOut_payload_199_2;
    _zz_dataOut_payload_200_24 <= _zz_dataOut_payload_200_23;
    _zz_dataOut_payload_201_3 <= _zz_dataOut_payload_201_2;
    _zz_dataOut_payload_202_6 <= _zz_dataOut_payload_202_5;
    _zz_dataOut_payload_203_3 <= _zz_dataOut_payload_203_2;
    _zz_dataOut_payload_204_12 <= _zz_dataOut_payload_204_11;
    _zz_dataOut_payload_205_3 <= _zz_dataOut_payload_205_2;
    _zz_dataOut_payload_206_6 <= _zz_dataOut_payload_206_5;
    _zz_dataOut_payload_207_3 <= _zz_dataOut_payload_207_2;
    _zz_dataOut_payload_208_48 <= _zz_dataOut_payload_208_47;
    _zz_dataOut_payload_209_3 <= _zz_dataOut_payload_209_2;
    _zz_dataOut_payload_210_6 <= _zz_dataOut_payload_210_5;
    _zz_dataOut_payload_211_3 <= _zz_dataOut_payload_211_2;
    _zz_dataOut_payload_212_12 <= _zz_dataOut_payload_212_11;
    _zz_dataOut_payload_213_3 <= _zz_dataOut_payload_213_2;
    _zz_dataOut_payload_214_6 <= _zz_dataOut_payload_214_5;
    _zz_dataOut_payload_215_3 <= _zz_dataOut_payload_215_2;
    _zz_dataOut_payload_216_24 <= _zz_dataOut_payload_216_23;
    _zz_dataOut_payload_217_3 <= _zz_dataOut_payload_217_2;
    _zz_dataOut_payload_218_6 <= _zz_dataOut_payload_218_5;
    _zz_dataOut_payload_219_3 <= _zz_dataOut_payload_219_2;
    _zz_dataOut_payload_220_12 <= _zz_dataOut_payload_220_11;
    _zz_dataOut_payload_221_3 <= _zz_dataOut_payload_221_2;
    _zz_dataOut_payload_222_6 <= _zz_dataOut_payload_222_5;
    _zz_dataOut_payload_223_3 <= _zz_dataOut_payload_223_2;
    _zz_dataOut_payload_224_93 <= (_zz_dataOut_payload_224_92 ? _zz_dataOut_payload_224_89 : _zz_dataOut_payload_224_91);
    _zz_dataOut_payload_225 <= (_zz_dataOut_payload_224_92 ? _zz_dataOut_payload_224_91 : _zz_dataOut_payload_224_89);
    _zz_dataOut_payload_226_3 <= (_zz_dataOut_payload_226_2 ? _zz_dataOut_payload_226 : _zz_dataOut_payload_226_1);
    _zz_dataOut_payload_227 <= (_zz_dataOut_payload_226_2 ? _zz_dataOut_payload_226_1 : _zz_dataOut_payload_226);
    _zz_dataOut_payload_228_9 <= (_zz_dataOut_payload_228_8 ? _zz_dataOut_payload_228_5 : _zz_dataOut_payload_228_7);
    _zz_dataOut_payload_229 <= (_zz_dataOut_payload_228_8 ? _zz_dataOut_payload_228_7 : _zz_dataOut_payload_228_5);
    _zz_dataOut_payload_230_3 <= (_zz_dataOut_payload_230_2 ? _zz_dataOut_payload_230 : _zz_dataOut_payload_230_1);
    _zz_dataOut_payload_231 <= (_zz_dataOut_payload_230_2 ? _zz_dataOut_payload_230_1 : _zz_dataOut_payload_230);
    _zz_dataOut_payload_224_94 <= _zz_dataOut_payload_224_93;
    _zz_dataOut_payload_225_1 <= _zz_dataOut_payload_225;
    _zz_dataOut_payload_226_4 <= _zz_dataOut_payload_226_3;
    _zz_dataOut_payload_227_1 <= _zz_dataOut_payload_227;
    _zz_dataOut_payload_228_10 <= _zz_dataOut_payload_228_9;
    _zz_dataOut_payload_229_1 <= _zz_dataOut_payload_229;
    _zz_dataOut_payload_230_4 <= _zz_dataOut_payload_230_3;
    _zz_dataOut_payload_231_1 <= _zz_dataOut_payload_231;
    _zz_dataOut_payload_232_21 <= (_zz_dataOut_payload_232_20 ? _zz_dataOut_payload_232_17 : _zz_dataOut_payload_232_19);
    _zz_dataOut_payload_233 <= (_zz_dataOut_payload_232_20 ? _zz_dataOut_payload_232_19 : _zz_dataOut_payload_232_17);
    _zz_dataOut_payload_234_3 <= (_zz_dataOut_payload_234_2 ? _zz_dataOut_payload_234 : _zz_dataOut_payload_234_1);
    _zz_dataOut_payload_235 <= (_zz_dataOut_payload_234_2 ? _zz_dataOut_payload_234_1 : _zz_dataOut_payload_234);
    _zz_dataOut_payload_236_9 <= (_zz_dataOut_payload_236_8 ? _zz_dataOut_payload_236_5 : _zz_dataOut_payload_236_7);
    _zz_dataOut_payload_237 <= (_zz_dataOut_payload_236_8 ? _zz_dataOut_payload_236_7 : _zz_dataOut_payload_236_5);
    _zz_dataOut_payload_238_3 <= (_zz_dataOut_payload_238_2 ? _zz_dataOut_payload_238 : _zz_dataOut_payload_238_1);
    _zz_dataOut_payload_239 <= (_zz_dataOut_payload_238_2 ? _zz_dataOut_payload_238_1 : _zz_dataOut_payload_238);
    _zz_dataOut_payload_232_22 <= _zz_dataOut_payload_232_21;
    _zz_dataOut_payload_233_1 <= _zz_dataOut_payload_233;
    _zz_dataOut_payload_234_4 <= _zz_dataOut_payload_234_3;
    _zz_dataOut_payload_235_1 <= _zz_dataOut_payload_235;
    _zz_dataOut_payload_236_10 <= _zz_dataOut_payload_236_9;
    _zz_dataOut_payload_237_1 <= _zz_dataOut_payload_237;
    _zz_dataOut_payload_238_4 <= _zz_dataOut_payload_238_3;
    _zz_dataOut_payload_239_1 <= _zz_dataOut_payload_239;
    _zz_dataOut_payload_224_95 <= _zz_dataOut_payload_224_94;
    _zz_dataOut_payload_225_2 <= _zz_dataOut_payload_225_1;
    _zz_dataOut_payload_226_5 <= _zz_dataOut_payload_226_4;
    _zz_dataOut_payload_227_2 <= _zz_dataOut_payload_227_1;
    _zz_dataOut_payload_228_11 <= _zz_dataOut_payload_228_10;
    _zz_dataOut_payload_229_2 <= _zz_dataOut_payload_229_1;
    _zz_dataOut_payload_230_5 <= _zz_dataOut_payload_230_4;
    _zz_dataOut_payload_231_2 <= _zz_dataOut_payload_231_1;
    _zz_dataOut_payload_232_23 <= _zz_dataOut_payload_232_22;
    _zz_dataOut_payload_233_2 <= _zz_dataOut_payload_233_1;
    _zz_dataOut_payload_234_5 <= _zz_dataOut_payload_234_4;
    _zz_dataOut_payload_235_2 <= _zz_dataOut_payload_235_1;
    _zz_dataOut_payload_236_11 <= _zz_dataOut_payload_236_10;
    _zz_dataOut_payload_237_2 <= _zz_dataOut_payload_237_1;
    _zz_dataOut_payload_238_5 <= _zz_dataOut_payload_238_4;
    _zz_dataOut_payload_239_2 <= _zz_dataOut_payload_239_1;
    _zz_dataOut_payload_240_45 <= (_zz_dataOut_payload_240_44 ? _zz_dataOut_payload_240_41 : _zz_dataOut_payload_240_43);
    _zz_dataOut_payload_241 <= (_zz_dataOut_payload_240_44 ? _zz_dataOut_payload_240_43 : _zz_dataOut_payload_240_41);
    _zz_dataOut_payload_242_3 <= (_zz_dataOut_payload_242_2 ? _zz_dataOut_payload_242 : _zz_dataOut_payload_242_1);
    _zz_dataOut_payload_243 <= (_zz_dataOut_payload_242_2 ? _zz_dataOut_payload_242_1 : _zz_dataOut_payload_242);
    _zz_dataOut_payload_244_9 <= (_zz_dataOut_payload_244_8 ? _zz_dataOut_payload_244_5 : _zz_dataOut_payload_244_7);
    _zz_dataOut_payload_245 <= (_zz_dataOut_payload_244_8 ? _zz_dataOut_payload_244_7 : _zz_dataOut_payload_244_5);
    _zz_dataOut_payload_246_3 <= (_zz_dataOut_payload_246_2 ? _zz_dataOut_payload_246 : _zz_dataOut_payload_246_1);
    _zz_dataOut_payload_247 <= (_zz_dataOut_payload_246_2 ? _zz_dataOut_payload_246_1 : _zz_dataOut_payload_246);
    _zz_dataOut_payload_240_46 <= _zz_dataOut_payload_240_45;
    _zz_dataOut_payload_241_1 <= _zz_dataOut_payload_241;
    _zz_dataOut_payload_242_4 <= _zz_dataOut_payload_242_3;
    _zz_dataOut_payload_243_1 <= _zz_dataOut_payload_243;
    _zz_dataOut_payload_244_10 <= _zz_dataOut_payload_244_9;
    _zz_dataOut_payload_245_1 <= _zz_dataOut_payload_245;
    _zz_dataOut_payload_246_4 <= _zz_dataOut_payload_246_3;
    _zz_dataOut_payload_247_1 <= _zz_dataOut_payload_247;
    _zz_dataOut_payload_248_21 <= (_zz_dataOut_payload_248_20 ? _zz_dataOut_payload_248_17 : _zz_dataOut_payload_248_19);
    _zz_dataOut_payload_249 <= (_zz_dataOut_payload_248_20 ? _zz_dataOut_payload_248_19 : _zz_dataOut_payload_248_17);
    _zz_dataOut_payload_250_3 <= (_zz_dataOut_payload_250_2 ? _zz_dataOut_payload_250 : _zz_dataOut_payload_250_1);
    _zz_dataOut_payload_251 <= (_zz_dataOut_payload_250_2 ? _zz_dataOut_payload_250_1 : _zz_dataOut_payload_250);
    _zz_dataOut_payload_252_9 <= (_zz_dataOut_payload_252_8 ? _zz_dataOut_payload_252_5 : _zz_dataOut_payload_252_7);
    _zz_dataOut_payload_253 <= (_zz_dataOut_payload_252_8 ? _zz_dataOut_payload_252_7 : _zz_dataOut_payload_252_5);
    _zz_dataOut_payload_254_3 <= (_zz_dataOut_payload_254_2 ? _zz_dataOut_payload_254 : _zz_dataOut_payload_254_1);
    _zz_dataOut_payload_255 <= (_zz_dataOut_payload_254_2 ? _zz_dataOut_payload_254_1 : _zz_dataOut_payload_254);
    _zz_dataOut_payload_248_22 <= _zz_dataOut_payload_248_21;
    _zz_dataOut_payload_249_1 <= _zz_dataOut_payload_249;
    _zz_dataOut_payload_250_4 <= _zz_dataOut_payload_250_3;
    _zz_dataOut_payload_251_1 <= _zz_dataOut_payload_251;
    _zz_dataOut_payload_252_10 <= _zz_dataOut_payload_252_9;
    _zz_dataOut_payload_253_1 <= _zz_dataOut_payload_253;
    _zz_dataOut_payload_254_4 <= _zz_dataOut_payload_254_3;
    _zz_dataOut_payload_255_1 <= _zz_dataOut_payload_255;
    _zz_dataOut_payload_240_47 <= _zz_dataOut_payload_240_46;
    _zz_dataOut_payload_241_2 <= _zz_dataOut_payload_241_1;
    _zz_dataOut_payload_242_5 <= _zz_dataOut_payload_242_4;
    _zz_dataOut_payload_243_2 <= _zz_dataOut_payload_243_1;
    _zz_dataOut_payload_244_11 <= _zz_dataOut_payload_244_10;
    _zz_dataOut_payload_245_2 <= _zz_dataOut_payload_245_1;
    _zz_dataOut_payload_246_5 <= _zz_dataOut_payload_246_4;
    _zz_dataOut_payload_247_2 <= _zz_dataOut_payload_247_1;
    _zz_dataOut_payload_248_23 <= _zz_dataOut_payload_248_22;
    _zz_dataOut_payload_249_2 <= _zz_dataOut_payload_249_1;
    _zz_dataOut_payload_250_5 <= _zz_dataOut_payload_250_4;
    _zz_dataOut_payload_251_2 <= _zz_dataOut_payload_251_1;
    _zz_dataOut_payload_252_11 <= _zz_dataOut_payload_252_10;
    _zz_dataOut_payload_253_2 <= _zz_dataOut_payload_253_1;
    _zz_dataOut_payload_254_5 <= _zz_dataOut_payload_254_4;
    _zz_dataOut_payload_255_2 <= _zz_dataOut_payload_255_1;
    _zz_dataOut_payload_224_96 <= _zz_dataOut_payload_224_95;
    _zz_dataOut_payload_225_3 <= _zz_dataOut_payload_225_2;
    _zz_dataOut_payload_226_6 <= _zz_dataOut_payload_226_5;
    _zz_dataOut_payload_227_3 <= _zz_dataOut_payload_227_2;
    _zz_dataOut_payload_228_12 <= _zz_dataOut_payload_228_11;
    _zz_dataOut_payload_229_3 <= _zz_dataOut_payload_229_2;
    _zz_dataOut_payload_230_6 <= _zz_dataOut_payload_230_5;
    _zz_dataOut_payload_231_3 <= _zz_dataOut_payload_231_2;
    _zz_dataOut_payload_232_24 <= _zz_dataOut_payload_232_23;
    _zz_dataOut_payload_233_3 <= _zz_dataOut_payload_233_2;
    _zz_dataOut_payload_234_6 <= _zz_dataOut_payload_234_5;
    _zz_dataOut_payload_235_3 <= _zz_dataOut_payload_235_2;
    _zz_dataOut_payload_236_12 <= _zz_dataOut_payload_236_11;
    _zz_dataOut_payload_237_3 <= _zz_dataOut_payload_237_2;
    _zz_dataOut_payload_238_6 <= _zz_dataOut_payload_238_5;
    _zz_dataOut_payload_239_3 <= _zz_dataOut_payload_239_2;
    _zz_dataOut_payload_240_48 <= _zz_dataOut_payload_240_47;
    _zz_dataOut_payload_241_3 <= _zz_dataOut_payload_241_2;
    _zz_dataOut_payload_242_6 <= _zz_dataOut_payload_242_5;
    _zz_dataOut_payload_243_3 <= _zz_dataOut_payload_243_2;
    _zz_dataOut_payload_244_12 <= _zz_dataOut_payload_244_11;
    _zz_dataOut_payload_245_3 <= _zz_dataOut_payload_245_2;
    _zz_dataOut_payload_246_6 <= _zz_dataOut_payload_246_5;
    _zz_dataOut_payload_247_3 <= _zz_dataOut_payload_247_2;
    _zz_dataOut_payload_248_24 <= _zz_dataOut_payload_248_23;
    _zz_dataOut_payload_249_3 <= _zz_dataOut_payload_249_2;
    _zz_dataOut_payload_250_6 <= _zz_dataOut_payload_250_5;
    _zz_dataOut_payload_251_3 <= _zz_dataOut_payload_251_2;
    _zz_dataOut_payload_252_12 <= _zz_dataOut_payload_252_11;
    _zz_dataOut_payload_253_3 <= _zz_dataOut_payload_253_2;
    _zz_dataOut_payload_254_6 <= _zz_dataOut_payload_254_5;
    _zz_dataOut_payload_255_3 <= _zz_dataOut_payload_255_2;
    _zz_dataOut_payload_192_193 <= _zz_dataOut_payload_192_192;
    _zz_dataOut_payload_193_4 <= _zz_dataOut_payload_193_3;
    _zz_dataOut_payload_194_7 <= _zz_dataOut_payload_194_6;
    _zz_dataOut_payload_195_4 <= _zz_dataOut_payload_195_3;
    _zz_dataOut_payload_196_13 <= _zz_dataOut_payload_196_12;
    _zz_dataOut_payload_197_4 <= _zz_dataOut_payload_197_3;
    _zz_dataOut_payload_198_7 <= _zz_dataOut_payload_198_6;
    _zz_dataOut_payload_199_4 <= _zz_dataOut_payload_199_3;
    _zz_dataOut_payload_200_25 <= _zz_dataOut_payload_200_24;
    _zz_dataOut_payload_201_4 <= _zz_dataOut_payload_201_3;
    _zz_dataOut_payload_202_7 <= _zz_dataOut_payload_202_6;
    _zz_dataOut_payload_203_4 <= _zz_dataOut_payload_203_3;
    _zz_dataOut_payload_204_13 <= _zz_dataOut_payload_204_12;
    _zz_dataOut_payload_205_4 <= _zz_dataOut_payload_205_3;
    _zz_dataOut_payload_206_7 <= _zz_dataOut_payload_206_6;
    _zz_dataOut_payload_207_4 <= _zz_dataOut_payload_207_3;
    _zz_dataOut_payload_208_49 <= _zz_dataOut_payload_208_48;
    _zz_dataOut_payload_209_4 <= _zz_dataOut_payload_209_3;
    _zz_dataOut_payload_210_7 <= _zz_dataOut_payload_210_6;
    _zz_dataOut_payload_211_4 <= _zz_dataOut_payload_211_3;
    _zz_dataOut_payload_212_13 <= _zz_dataOut_payload_212_12;
    _zz_dataOut_payload_213_4 <= _zz_dataOut_payload_213_3;
    _zz_dataOut_payload_214_7 <= _zz_dataOut_payload_214_6;
    _zz_dataOut_payload_215_4 <= _zz_dataOut_payload_215_3;
    _zz_dataOut_payload_216_25 <= _zz_dataOut_payload_216_24;
    _zz_dataOut_payload_217_4 <= _zz_dataOut_payload_217_3;
    _zz_dataOut_payload_218_7 <= _zz_dataOut_payload_218_6;
    _zz_dataOut_payload_219_4 <= _zz_dataOut_payload_219_3;
    _zz_dataOut_payload_220_13 <= _zz_dataOut_payload_220_12;
    _zz_dataOut_payload_221_4 <= _zz_dataOut_payload_221_3;
    _zz_dataOut_payload_222_7 <= _zz_dataOut_payload_222_6;
    _zz_dataOut_payload_223_4 <= _zz_dataOut_payload_223_3;
    _zz_dataOut_payload_224_97 <= _zz_dataOut_payload_224_96;
    _zz_dataOut_payload_225_4 <= _zz_dataOut_payload_225_3;
    _zz_dataOut_payload_226_7 <= _zz_dataOut_payload_226_6;
    _zz_dataOut_payload_227_4 <= _zz_dataOut_payload_227_3;
    _zz_dataOut_payload_228_13 <= _zz_dataOut_payload_228_12;
    _zz_dataOut_payload_229_4 <= _zz_dataOut_payload_229_3;
    _zz_dataOut_payload_230_7 <= _zz_dataOut_payload_230_6;
    _zz_dataOut_payload_231_4 <= _zz_dataOut_payload_231_3;
    _zz_dataOut_payload_232_25 <= _zz_dataOut_payload_232_24;
    _zz_dataOut_payload_233_4 <= _zz_dataOut_payload_233_3;
    _zz_dataOut_payload_234_7 <= _zz_dataOut_payload_234_6;
    _zz_dataOut_payload_235_4 <= _zz_dataOut_payload_235_3;
    _zz_dataOut_payload_236_13 <= _zz_dataOut_payload_236_12;
    _zz_dataOut_payload_237_4 <= _zz_dataOut_payload_237_3;
    _zz_dataOut_payload_238_7 <= _zz_dataOut_payload_238_6;
    _zz_dataOut_payload_239_4 <= _zz_dataOut_payload_239_3;
    _zz_dataOut_payload_240_49 <= _zz_dataOut_payload_240_48;
    _zz_dataOut_payload_241_4 <= _zz_dataOut_payload_241_3;
    _zz_dataOut_payload_242_7 <= _zz_dataOut_payload_242_6;
    _zz_dataOut_payload_243_4 <= _zz_dataOut_payload_243_3;
    _zz_dataOut_payload_244_13 <= _zz_dataOut_payload_244_12;
    _zz_dataOut_payload_245_4 <= _zz_dataOut_payload_245_3;
    _zz_dataOut_payload_246_7 <= _zz_dataOut_payload_246_6;
    _zz_dataOut_payload_247_4 <= _zz_dataOut_payload_247_3;
    _zz_dataOut_payload_248_25 <= _zz_dataOut_payload_248_24;
    _zz_dataOut_payload_249_4 <= _zz_dataOut_payload_249_3;
    _zz_dataOut_payload_250_7 <= _zz_dataOut_payload_250_6;
    _zz_dataOut_payload_251_4 <= _zz_dataOut_payload_251_3;
    _zz_dataOut_payload_252_13 <= _zz_dataOut_payload_252_12;
    _zz_dataOut_payload_253_4 <= _zz_dataOut_payload_253_3;
    _zz_dataOut_payload_254_7 <= _zz_dataOut_payload_254_6;
    _zz_dataOut_payload_255_4 <= _zz_dataOut_payload_255_3;
    _zz_dataOut_payload_128_386 <= _zz_dataOut_payload_128_385;
    _zz_dataOut_payload_129_5 <= _zz_dataOut_payload_129_4;
    _zz_dataOut_payload_130_8 <= _zz_dataOut_payload_130_7;
    _zz_dataOut_payload_131_5 <= _zz_dataOut_payload_131_4;
    _zz_dataOut_payload_132_14 <= _zz_dataOut_payload_132_13;
    _zz_dataOut_payload_133_5 <= _zz_dataOut_payload_133_4;
    _zz_dataOut_payload_134_8 <= _zz_dataOut_payload_134_7;
    _zz_dataOut_payload_135_5 <= _zz_dataOut_payload_135_4;
    _zz_dataOut_payload_136_26 <= _zz_dataOut_payload_136_25;
    _zz_dataOut_payload_137_5 <= _zz_dataOut_payload_137_4;
    _zz_dataOut_payload_138_8 <= _zz_dataOut_payload_138_7;
    _zz_dataOut_payload_139_5 <= _zz_dataOut_payload_139_4;
    _zz_dataOut_payload_140_14 <= _zz_dataOut_payload_140_13;
    _zz_dataOut_payload_141_5 <= _zz_dataOut_payload_141_4;
    _zz_dataOut_payload_142_8 <= _zz_dataOut_payload_142_7;
    _zz_dataOut_payload_143_5 <= _zz_dataOut_payload_143_4;
    _zz_dataOut_payload_144_50 <= _zz_dataOut_payload_144_49;
    _zz_dataOut_payload_145_5 <= _zz_dataOut_payload_145_4;
    _zz_dataOut_payload_146_8 <= _zz_dataOut_payload_146_7;
    _zz_dataOut_payload_147_5 <= _zz_dataOut_payload_147_4;
    _zz_dataOut_payload_148_14 <= _zz_dataOut_payload_148_13;
    _zz_dataOut_payload_149_5 <= _zz_dataOut_payload_149_4;
    _zz_dataOut_payload_150_8 <= _zz_dataOut_payload_150_7;
    _zz_dataOut_payload_151_5 <= _zz_dataOut_payload_151_4;
    _zz_dataOut_payload_152_26 <= _zz_dataOut_payload_152_25;
    _zz_dataOut_payload_153_5 <= _zz_dataOut_payload_153_4;
    _zz_dataOut_payload_154_8 <= _zz_dataOut_payload_154_7;
    _zz_dataOut_payload_155_5 <= _zz_dataOut_payload_155_4;
    _zz_dataOut_payload_156_14 <= _zz_dataOut_payload_156_13;
    _zz_dataOut_payload_157_5 <= _zz_dataOut_payload_157_4;
    _zz_dataOut_payload_158_8 <= _zz_dataOut_payload_158_7;
    _zz_dataOut_payload_159_5 <= _zz_dataOut_payload_159_4;
    _zz_dataOut_payload_160_98 <= _zz_dataOut_payload_160_97;
    _zz_dataOut_payload_161_5 <= _zz_dataOut_payload_161_4;
    _zz_dataOut_payload_162_8 <= _zz_dataOut_payload_162_7;
    _zz_dataOut_payload_163_5 <= _zz_dataOut_payload_163_4;
    _zz_dataOut_payload_164_14 <= _zz_dataOut_payload_164_13;
    _zz_dataOut_payload_165_5 <= _zz_dataOut_payload_165_4;
    _zz_dataOut_payload_166_8 <= _zz_dataOut_payload_166_7;
    _zz_dataOut_payload_167_5 <= _zz_dataOut_payload_167_4;
    _zz_dataOut_payload_168_26 <= _zz_dataOut_payload_168_25;
    _zz_dataOut_payload_169_5 <= _zz_dataOut_payload_169_4;
    _zz_dataOut_payload_170_8 <= _zz_dataOut_payload_170_7;
    _zz_dataOut_payload_171_5 <= _zz_dataOut_payload_171_4;
    _zz_dataOut_payload_172_14 <= _zz_dataOut_payload_172_13;
    _zz_dataOut_payload_173_5 <= _zz_dataOut_payload_173_4;
    _zz_dataOut_payload_174_8 <= _zz_dataOut_payload_174_7;
    _zz_dataOut_payload_175_5 <= _zz_dataOut_payload_175_4;
    _zz_dataOut_payload_176_50 <= _zz_dataOut_payload_176_49;
    _zz_dataOut_payload_177_5 <= _zz_dataOut_payload_177_4;
    _zz_dataOut_payload_178_8 <= _zz_dataOut_payload_178_7;
    _zz_dataOut_payload_179_5 <= _zz_dataOut_payload_179_4;
    _zz_dataOut_payload_180_14 <= _zz_dataOut_payload_180_13;
    _zz_dataOut_payload_181_5 <= _zz_dataOut_payload_181_4;
    _zz_dataOut_payload_182_8 <= _zz_dataOut_payload_182_7;
    _zz_dataOut_payload_183_5 <= _zz_dataOut_payload_183_4;
    _zz_dataOut_payload_184_26 <= _zz_dataOut_payload_184_25;
    _zz_dataOut_payload_185_5 <= _zz_dataOut_payload_185_4;
    _zz_dataOut_payload_186_8 <= _zz_dataOut_payload_186_7;
    _zz_dataOut_payload_187_5 <= _zz_dataOut_payload_187_4;
    _zz_dataOut_payload_188_14 <= _zz_dataOut_payload_188_13;
    _zz_dataOut_payload_189_5 <= _zz_dataOut_payload_189_4;
    _zz_dataOut_payload_190_8 <= _zz_dataOut_payload_190_7;
    _zz_dataOut_payload_191_5 <= _zz_dataOut_payload_191_4;
    _zz_dataOut_payload_192_194 <= _zz_dataOut_payload_192_193;
    _zz_dataOut_payload_193_5 <= _zz_dataOut_payload_193_4;
    _zz_dataOut_payload_194_8 <= _zz_dataOut_payload_194_7;
    _zz_dataOut_payload_195_5 <= _zz_dataOut_payload_195_4;
    _zz_dataOut_payload_196_14 <= _zz_dataOut_payload_196_13;
    _zz_dataOut_payload_197_5 <= _zz_dataOut_payload_197_4;
    _zz_dataOut_payload_198_8 <= _zz_dataOut_payload_198_7;
    _zz_dataOut_payload_199_5 <= _zz_dataOut_payload_199_4;
    _zz_dataOut_payload_200_26 <= _zz_dataOut_payload_200_25;
    _zz_dataOut_payload_201_5 <= _zz_dataOut_payload_201_4;
    _zz_dataOut_payload_202_8 <= _zz_dataOut_payload_202_7;
    _zz_dataOut_payload_203_5 <= _zz_dataOut_payload_203_4;
    _zz_dataOut_payload_204_14 <= _zz_dataOut_payload_204_13;
    _zz_dataOut_payload_205_5 <= _zz_dataOut_payload_205_4;
    _zz_dataOut_payload_206_8 <= _zz_dataOut_payload_206_7;
    _zz_dataOut_payload_207_5 <= _zz_dataOut_payload_207_4;
    _zz_dataOut_payload_208_50 <= _zz_dataOut_payload_208_49;
    _zz_dataOut_payload_209_5 <= _zz_dataOut_payload_209_4;
    _zz_dataOut_payload_210_8 <= _zz_dataOut_payload_210_7;
    _zz_dataOut_payload_211_5 <= _zz_dataOut_payload_211_4;
    _zz_dataOut_payload_212_14 <= _zz_dataOut_payload_212_13;
    _zz_dataOut_payload_213_5 <= _zz_dataOut_payload_213_4;
    _zz_dataOut_payload_214_8 <= _zz_dataOut_payload_214_7;
    _zz_dataOut_payload_215_5 <= _zz_dataOut_payload_215_4;
    _zz_dataOut_payload_216_26 <= _zz_dataOut_payload_216_25;
    _zz_dataOut_payload_217_5 <= _zz_dataOut_payload_217_4;
    _zz_dataOut_payload_218_8 <= _zz_dataOut_payload_218_7;
    _zz_dataOut_payload_219_5 <= _zz_dataOut_payload_219_4;
    _zz_dataOut_payload_220_14 <= _zz_dataOut_payload_220_13;
    _zz_dataOut_payload_221_5 <= _zz_dataOut_payload_221_4;
    _zz_dataOut_payload_222_8 <= _zz_dataOut_payload_222_7;
    _zz_dataOut_payload_223_5 <= _zz_dataOut_payload_223_4;
    _zz_dataOut_payload_224_98 <= _zz_dataOut_payload_224_97;
    _zz_dataOut_payload_225_5 <= _zz_dataOut_payload_225_4;
    _zz_dataOut_payload_226_8 <= _zz_dataOut_payload_226_7;
    _zz_dataOut_payload_227_5 <= _zz_dataOut_payload_227_4;
    _zz_dataOut_payload_228_14 <= _zz_dataOut_payload_228_13;
    _zz_dataOut_payload_229_5 <= _zz_dataOut_payload_229_4;
    _zz_dataOut_payload_230_8 <= _zz_dataOut_payload_230_7;
    _zz_dataOut_payload_231_5 <= _zz_dataOut_payload_231_4;
    _zz_dataOut_payload_232_26 <= _zz_dataOut_payload_232_25;
    _zz_dataOut_payload_233_5 <= _zz_dataOut_payload_233_4;
    _zz_dataOut_payload_234_8 <= _zz_dataOut_payload_234_7;
    _zz_dataOut_payload_235_5 <= _zz_dataOut_payload_235_4;
    _zz_dataOut_payload_236_14 <= _zz_dataOut_payload_236_13;
    _zz_dataOut_payload_237_5 <= _zz_dataOut_payload_237_4;
    _zz_dataOut_payload_238_8 <= _zz_dataOut_payload_238_7;
    _zz_dataOut_payload_239_5 <= _zz_dataOut_payload_239_4;
    _zz_dataOut_payload_240_50 <= _zz_dataOut_payload_240_49;
    _zz_dataOut_payload_241_5 <= _zz_dataOut_payload_241_4;
    _zz_dataOut_payload_242_8 <= _zz_dataOut_payload_242_7;
    _zz_dataOut_payload_243_5 <= _zz_dataOut_payload_243_4;
    _zz_dataOut_payload_244_14 <= _zz_dataOut_payload_244_13;
    _zz_dataOut_payload_245_5 <= _zz_dataOut_payload_245_4;
    _zz_dataOut_payload_246_8 <= _zz_dataOut_payload_246_7;
    _zz_dataOut_payload_247_5 <= _zz_dataOut_payload_247_4;
    _zz_dataOut_payload_248_26 <= _zz_dataOut_payload_248_25;
    _zz_dataOut_payload_249_5 <= _zz_dataOut_payload_249_4;
    _zz_dataOut_payload_250_8 <= _zz_dataOut_payload_250_7;
    _zz_dataOut_payload_251_5 <= _zz_dataOut_payload_251_4;
    _zz_dataOut_payload_252_14 <= _zz_dataOut_payload_252_13;
    _zz_dataOut_payload_253_5 <= _zz_dataOut_payload_253_4;
    _zz_dataOut_payload_254_8 <= _zz_dataOut_payload_254_7;
    _zz_dataOut_payload_255_5 <= _zz_dataOut_payload_255_4;
    _zz_dataOut_payload_0_16643 <= _zz_dataOut_payload_0_16642;
    _zz_dataOut_payload_1_6 <= _zz_dataOut_payload_1_5;
    _zz_dataOut_payload_2_9 <= _zz_dataOut_payload_2_8;
    _zz_dataOut_payload_3_6 <= _zz_dataOut_payload_3_5;
    _zz_dataOut_payload_4_15 <= _zz_dataOut_payload_4_14;
    _zz_dataOut_payload_5_6 <= _zz_dataOut_payload_5_5;
    _zz_dataOut_payload_6_9 <= _zz_dataOut_payload_6_8;
    _zz_dataOut_payload_7_6 <= _zz_dataOut_payload_7_5;
    _zz_dataOut_payload_8_27 <= _zz_dataOut_payload_8_26;
    _zz_dataOut_payload_9_6 <= _zz_dataOut_payload_9_5;
    _zz_dataOut_payload_10_9 <= _zz_dataOut_payload_10_8;
    _zz_dataOut_payload_11_6 <= _zz_dataOut_payload_11_5;
    _zz_dataOut_payload_12_15 <= _zz_dataOut_payload_12_14;
    _zz_dataOut_payload_13_6 <= _zz_dataOut_payload_13_5;
    _zz_dataOut_payload_14_9 <= _zz_dataOut_payload_14_8;
    _zz_dataOut_payload_15_6 <= _zz_dataOut_payload_15_5;
    _zz_dataOut_payload_16_51 <= _zz_dataOut_payload_16_50;
    _zz_dataOut_payload_17_6 <= _zz_dataOut_payload_17_5;
    _zz_dataOut_payload_18_9 <= _zz_dataOut_payload_18_8;
    _zz_dataOut_payload_19_6 <= _zz_dataOut_payload_19_5;
    _zz_dataOut_payload_20_15 <= _zz_dataOut_payload_20_14;
    _zz_dataOut_payload_21_6 <= _zz_dataOut_payload_21_5;
    _zz_dataOut_payload_22_9 <= _zz_dataOut_payload_22_8;
    _zz_dataOut_payload_23_6 <= _zz_dataOut_payload_23_5;
    _zz_dataOut_payload_24_27 <= _zz_dataOut_payload_24_26;
    _zz_dataOut_payload_25_6 <= _zz_dataOut_payload_25_5;
    _zz_dataOut_payload_26_9 <= _zz_dataOut_payload_26_8;
    _zz_dataOut_payload_27_6 <= _zz_dataOut_payload_27_5;
    _zz_dataOut_payload_28_15 <= _zz_dataOut_payload_28_14;
    _zz_dataOut_payload_29_6 <= _zz_dataOut_payload_29_5;
    _zz_dataOut_payload_30_9 <= _zz_dataOut_payload_30_8;
    _zz_dataOut_payload_31_6 <= _zz_dataOut_payload_31_5;
    _zz_dataOut_payload_32_99 <= _zz_dataOut_payload_32_98;
    _zz_dataOut_payload_33_6 <= _zz_dataOut_payload_33_5;
    _zz_dataOut_payload_34_9 <= _zz_dataOut_payload_34_8;
    _zz_dataOut_payload_35_6 <= _zz_dataOut_payload_35_5;
    _zz_dataOut_payload_36_15 <= _zz_dataOut_payload_36_14;
    _zz_dataOut_payload_37_6 <= _zz_dataOut_payload_37_5;
    _zz_dataOut_payload_38_9 <= _zz_dataOut_payload_38_8;
    _zz_dataOut_payload_39_6 <= _zz_dataOut_payload_39_5;
    _zz_dataOut_payload_40_27 <= _zz_dataOut_payload_40_26;
    _zz_dataOut_payload_41_6 <= _zz_dataOut_payload_41_5;
    _zz_dataOut_payload_42_9 <= _zz_dataOut_payload_42_8;
    _zz_dataOut_payload_43_6 <= _zz_dataOut_payload_43_5;
    _zz_dataOut_payload_44_15 <= _zz_dataOut_payload_44_14;
    _zz_dataOut_payload_45_6 <= _zz_dataOut_payload_45_5;
    _zz_dataOut_payload_46_9 <= _zz_dataOut_payload_46_8;
    _zz_dataOut_payload_47_6 <= _zz_dataOut_payload_47_5;
    _zz_dataOut_payload_48_51 <= _zz_dataOut_payload_48_50;
    _zz_dataOut_payload_49_6 <= _zz_dataOut_payload_49_5;
    _zz_dataOut_payload_50_9 <= _zz_dataOut_payload_50_8;
    _zz_dataOut_payload_51_6 <= _zz_dataOut_payload_51_5;
    _zz_dataOut_payload_52_15 <= _zz_dataOut_payload_52_14;
    _zz_dataOut_payload_53_6 <= _zz_dataOut_payload_53_5;
    _zz_dataOut_payload_54_9 <= _zz_dataOut_payload_54_8;
    _zz_dataOut_payload_55_6 <= _zz_dataOut_payload_55_5;
    _zz_dataOut_payload_56_27 <= _zz_dataOut_payload_56_26;
    _zz_dataOut_payload_57_6 <= _zz_dataOut_payload_57_5;
    _zz_dataOut_payload_58_9 <= _zz_dataOut_payload_58_8;
    _zz_dataOut_payload_59_6 <= _zz_dataOut_payload_59_5;
    _zz_dataOut_payload_60_15 <= _zz_dataOut_payload_60_14;
    _zz_dataOut_payload_61_6 <= _zz_dataOut_payload_61_5;
    _zz_dataOut_payload_62_9 <= _zz_dataOut_payload_62_8;
    _zz_dataOut_payload_63_6 <= _zz_dataOut_payload_63_5;
    _zz_dataOut_payload_64_195 <= _zz_dataOut_payload_64_194;
    _zz_dataOut_payload_65_6 <= _zz_dataOut_payload_65_5;
    _zz_dataOut_payload_66_9 <= _zz_dataOut_payload_66_8;
    _zz_dataOut_payload_67_6 <= _zz_dataOut_payload_67_5;
    _zz_dataOut_payload_68_15 <= _zz_dataOut_payload_68_14;
    _zz_dataOut_payload_69_6 <= _zz_dataOut_payload_69_5;
    _zz_dataOut_payload_70_9 <= _zz_dataOut_payload_70_8;
    _zz_dataOut_payload_71_6 <= _zz_dataOut_payload_71_5;
    _zz_dataOut_payload_72_27 <= _zz_dataOut_payload_72_26;
    _zz_dataOut_payload_73_6 <= _zz_dataOut_payload_73_5;
    _zz_dataOut_payload_74_9 <= _zz_dataOut_payload_74_8;
    _zz_dataOut_payload_75_6 <= _zz_dataOut_payload_75_5;
    _zz_dataOut_payload_76_15 <= _zz_dataOut_payload_76_14;
    _zz_dataOut_payload_77_6 <= _zz_dataOut_payload_77_5;
    _zz_dataOut_payload_78_9 <= _zz_dataOut_payload_78_8;
    _zz_dataOut_payload_79_6 <= _zz_dataOut_payload_79_5;
    _zz_dataOut_payload_80_51 <= _zz_dataOut_payload_80_50;
    _zz_dataOut_payload_81_6 <= _zz_dataOut_payload_81_5;
    _zz_dataOut_payload_82_9 <= _zz_dataOut_payload_82_8;
    _zz_dataOut_payload_83_6 <= _zz_dataOut_payload_83_5;
    _zz_dataOut_payload_84_15 <= _zz_dataOut_payload_84_14;
    _zz_dataOut_payload_85_6 <= _zz_dataOut_payload_85_5;
    _zz_dataOut_payload_86_9 <= _zz_dataOut_payload_86_8;
    _zz_dataOut_payload_87_6 <= _zz_dataOut_payload_87_5;
    _zz_dataOut_payload_88_27 <= _zz_dataOut_payload_88_26;
    _zz_dataOut_payload_89_6 <= _zz_dataOut_payload_89_5;
    _zz_dataOut_payload_90_9 <= _zz_dataOut_payload_90_8;
    _zz_dataOut_payload_91_6 <= _zz_dataOut_payload_91_5;
    _zz_dataOut_payload_92_15 <= _zz_dataOut_payload_92_14;
    _zz_dataOut_payload_93_6 <= _zz_dataOut_payload_93_5;
    _zz_dataOut_payload_94_9 <= _zz_dataOut_payload_94_8;
    _zz_dataOut_payload_95_6 <= _zz_dataOut_payload_95_5;
    _zz_dataOut_payload_96_99 <= _zz_dataOut_payload_96_98;
    _zz_dataOut_payload_97_6 <= _zz_dataOut_payload_97_5;
    _zz_dataOut_payload_98_9 <= _zz_dataOut_payload_98_8;
    _zz_dataOut_payload_99_6 <= _zz_dataOut_payload_99_5;
    _zz_dataOut_payload_100_15 <= _zz_dataOut_payload_100_14;
    _zz_dataOut_payload_101_6 <= _zz_dataOut_payload_101_5;
    _zz_dataOut_payload_102_9 <= _zz_dataOut_payload_102_8;
    _zz_dataOut_payload_103_6 <= _zz_dataOut_payload_103_5;
    _zz_dataOut_payload_104_27 <= _zz_dataOut_payload_104_26;
    _zz_dataOut_payload_105_6 <= _zz_dataOut_payload_105_5;
    _zz_dataOut_payload_106_9 <= _zz_dataOut_payload_106_8;
    _zz_dataOut_payload_107_6 <= _zz_dataOut_payload_107_5;
    _zz_dataOut_payload_108_15 <= _zz_dataOut_payload_108_14;
    _zz_dataOut_payload_109_6 <= _zz_dataOut_payload_109_5;
    _zz_dataOut_payload_110_9 <= _zz_dataOut_payload_110_8;
    _zz_dataOut_payload_111_6 <= _zz_dataOut_payload_111_5;
    _zz_dataOut_payload_112_51 <= _zz_dataOut_payload_112_50;
    _zz_dataOut_payload_113_6 <= _zz_dataOut_payload_113_5;
    _zz_dataOut_payload_114_9 <= _zz_dataOut_payload_114_8;
    _zz_dataOut_payload_115_6 <= _zz_dataOut_payload_115_5;
    _zz_dataOut_payload_116_15 <= _zz_dataOut_payload_116_14;
    _zz_dataOut_payload_117_6 <= _zz_dataOut_payload_117_5;
    _zz_dataOut_payload_118_9 <= _zz_dataOut_payload_118_8;
    _zz_dataOut_payload_119_6 <= _zz_dataOut_payload_119_5;
    _zz_dataOut_payload_120_27 <= _zz_dataOut_payload_120_26;
    _zz_dataOut_payload_121_6 <= _zz_dataOut_payload_121_5;
    _zz_dataOut_payload_122_9 <= _zz_dataOut_payload_122_8;
    _zz_dataOut_payload_123_6 <= _zz_dataOut_payload_123_5;
    _zz_dataOut_payload_124_15 <= _zz_dataOut_payload_124_14;
    _zz_dataOut_payload_125_6 <= _zz_dataOut_payload_125_5;
    _zz_dataOut_payload_126_9 <= _zz_dataOut_payload_126_8;
    _zz_dataOut_payload_127_6 <= _zz_dataOut_payload_127_5;
    _zz_dataOut_payload_128_387 <= _zz_dataOut_payload_128_386;
    _zz_dataOut_payload_129_6 <= _zz_dataOut_payload_129_5;
    _zz_dataOut_payload_130_9 <= _zz_dataOut_payload_130_8;
    _zz_dataOut_payload_131_6 <= _zz_dataOut_payload_131_5;
    _zz_dataOut_payload_132_15 <= _zz_dataOut_payload_132_14;
    _zz_dataOut_payload_133_6 <= _zz_dataOut_payload_133_5;
    _zz_dataOut_payload_134_9 <= _zz_dataOut_payload_134_8;
    _zz_dataOut_payload_135_6 <= _zz_dataOut_payload_135_5;
    _zz_dataOut_payload_136_27 <= _zz_dataOut_payload_136_26;
    _zz_dataOut_payload_137_6 <= _zz_dataOut_payload_137_5;
    _zz_dataOut_payload_138_9 <= _zz_dataOut_payload_138_8;
    _zz_dataOut_payload_139_6 <= _zz_dataOut_payload_139_5;
    _zz_dataOut_payload_140_15 <= _zz_dataOut_payload_140_14;
    _zz_dataOut_payload_141_6 <= _zz_dataOut_payload_141_5;
    _zz_dataOut_payload_142_9 <= _zz_dataOut_payload_142_8;
    _zz_dataOut_payload_143_6 <= _zz_dataOut_payload_143_5;
    _zz_dataOut_payload_144_51 <= _zz_dataOut_payload_144_50;
    _zz_dataOut_payload_145_6 <= _zz_dataOut_payload_145_5;
    _zz_dataOut_payload_146_9 <= _zz_dataOut_payload_146_8;
    _zz_dataOut_payload_147_6 <= _zz_dataOut_payload_147_5;
    _zz_dataOut_payload_148_15 <= _zz_dataOut_payload_148_14;
    _zz_dataOut_payload_149_6 <= _zz_dataOut_payload_149_5;
    _zz_dataOut_payload_150_9 <= _zz_dataOut_payload_150_8;
    _zz_dataOut_payload_151_6 <= _zz_dataOut_payload_151_5;
    _zz_dataOut_payload_152_27 <= _zz_dataOut_payload_152_26;
    _zz_dataOut_payload_153_6 <= _zz_dataOut_payload_153_5;
    _zz_dataOut_payload_154_9 <= _zz_dataOut_payload_154_8;
    _zz_dataOut_payload_155_6 <= _zz_dataOut_payload_155_5;
    _zz_dataOut_payload_156_15 <= _zz_dataOut_payload_156_14;
    _zz_dataOut_payload_157_6 <= _zz_dataOut_payload_157_5;
    _zz_dataOut_payload_158_9 <= _zz_dataOut_payload_158_8;
    _zz_dataOut_payload_159_6 <= _zz_dataOut_payload_159_5;
    _zz_dataOut_payload_160_99 <= _zz_dataOut_payload_160_98;
    _zz_dataOut_payload_161_6 <= _zz_dataOut_payload_161_5;
    _zz_dataOut_payload_162_9 <= _zz_dataOut_payload_162_8;
    _zz_dataOut_payload_163_6 <= _zz_dataOut_payload_163_5;
    _zz_dataOut_payload_164_15 <= _zz_dataOut_payload_164_14;
    _zz_dataOut_payload_165_6 <= _zz_dataOut_payload_165_5;
    _zz_dataOut_payload_166_9 <= _zz_dataOut_payload_166_8;
    _zz_dataOut_payload_167_6 <= _zz_dataOut_payload_167_5;
    _zz_dataOut_payload_168_27 <= _zz_dataOut_payload_168_26;
    _zz_dataOut_payload_169_6 <= _zz_dataOut_payload_169_5;
    _zz_dataOut_payload_170_9 <= _zz_dataOut_payload_170_8;
    _zz_dataOut_payload_171_6 <= _zz_dataOut_payload_171_5;
    _zz_dataOut_payload_172_15 <= _zz_dataOut_payload_172_14;
    _zz_dataOut_payload_173_6 <= _zz_dataOut_payload_173_5;
    _zz_dataOut_payload_174_9 <= _zz_dataOut_payload_174_8;
    _zz_dataOut_payload_175_6 <= _zz_dataOut_payload_175_5;
    _zz_dataOut_payload_176_51 <= _zz_dataOut_payload_176_50;
    _zz_dataOut_payload_177_6 <= _zz_dataOut_payload_177_5;
    _zz_dataOut_payload_178_9 <= _zz_dataOut_payload_178_8;
    _zz_dataOut_payload_179_6 <= _zz_dataOut_payload_179_5;
    _zz_dataOut_payload_180_15 <= _zz_dataOut_payload_180_14;
    _zz_dataOut_payload_181_6 <= _zz_dataOut_payload_181_5;
    _zz_dataOut_payload_182_9 <= _zz_dataOut_payload_182_8;
    _zz_dataOut_payload_183_6 <= _zz_dataOut_payload_183_5;
    _zz_dataOut_payload_184_27 <= _zz_dataOut_payload_184_26;
    _zz_dataOut_payload_185_6 <= _zz_dataOut_payload_185_5;
    _zz_dataOut_payload_186_9 <= _zz_dataOut_payload_186_8;
    _zz_dataOut_payload_187_6 <= _zz_dataOut_payload_187_5;
    _zz_dataOut_payload_188_15 <= _zz_dataOut_payload_188_14;
    _zz_dataOut_payload_189_6 <= _zz_dataOut_payload_189_5;
    _zz_dataOut_payload_190_9 <= _zz_dataOut_payload_190_8;
    _zz_dataOut_payload_191_6 <= _zz_dataOut_payload_191_5;
    _zz_dataOut_payload_192_195 <= _zz_dataOut_payload_192_194;
    _zz_dataOut_payload_193_6 <= _zz_dataOut_payload_193_5;
    _zz_dataOut_payload_194_9 <= _zz_dataOut_payload_194_8;
    _zz_dataOut_payload_195_6 <= _zz_dataOut_payload_195_5;
    _zz_dataOut_payload_196_15 <= _zz_dataOut_payload_196_14;
    _zz_dataOut_payload_197_6 <= _zz_dataOut_payload_197_5;
    _zz_dataOut_payload_198_9 <= _zz_dataOut_payload_198_8;
    _zz_dataOut_payload_199_6 <= _zz_dataOut_payload_199_5;
    _zz_dataOut_payload_200_27 <= _zz_dataOut_payload_200_26;
    _zz_dataOut_payload_201_6 <= _zz_dataOut_payload_201_5;
    _zz_dataOut_payload_202_9 <= _zz_dataOut_payload_202_8;
    _zz_dataOut_payload_203_6 <= _zz_dataOut_payload_203_5;
    _zz_dataOut_payload_204_15 <= _zz_dataOut_payload_204_14;
    _zz_dataOut_payload_205_6 <= _zz_dataOut_payload_205_5;
    _zz_dataOut_payload_206_9 <= _zz_dataOut_payload_206_8;
    _zz_dataOut_payload_207_6 <= _zz_dataOut_payload_207_5;
    _zz_dataOut_payload_208_51 <= _zz_dataOut_payload_208_50;
    _zz_dataOut_payload_209_6 <= _zz_dataOut_payload_209_5;
    _zz_dataOut_payload_210_9 <= _zz_dataOut_payload_210_8;
    _zz_dataOut_payload_211_6 <= _zz_dataOut_payload_211_5;
    _zz_dataOut_payload_212_15 <= _zz_dataOut_payload_212_14;
    _zz_dataOut_payload_213_6 <= _zz_dataOut_payload_213_5;
    _zz_dataOut_payload_214_9 <= _zz_dataOut_payload_214_8;
    _zz_dataOut_payload_215_6 <= _zz_dataOut_payload_215_5;
    _zz_dataOut_payload_216_27 <= _zz_dataOut_payload_216_26;
    _zz_dataOut_payload_217_6 <= _zz_dataOut_payload_217_5;
    _zz_dataOut_payload_218_9 <= _zz_dataOut_payload_218_8;
    _zz_dataOut_payload_219_6 <= _zz_dataOut_payload_219_5;
    _zz_dataOut_payload_220_15 <= _zz_dataOut_payload_220_14;
    _zz_dataOut_payload_221_6 <= _zz_dataOut_payload_221_5;
    _zz_dataOut_payload_222_9 <= _zz_dataOut_payload_222_8;
    _zz_dataOut_payload_223_6 <= _zz_dataOut_payload_223_5;
    _zz_dataOut_payload_224_99 <= _zz_dataOut_payload_224_98;
    _zz_dataOut_payload_225_6 <= _zz_dataOut_payload_225_5;
    _zz_dataOut_payload_226_9 <= _zz_dataOut_payload_226_8;
    _zz_dataOut_payload_227_6 <= _zz_dataOut_payload_227_5;
    _zz_dataOut_payload_228_15 <= _zz_dataOut_payload_228_14;
    _zz_dataOut_payload_229_6 <= _zz_dataOut_payload_229_5;
    _zz_dataOut_payload_230_9 <= _zz_dataOut_payload_230_8;
    _zz_dataOut_payload_231_6 <= _zz_dataOut_payload_231_5;
    _zz_dataOut_payload_232_27 <= _zz_dataOut_payload_232_26;
    _zz_dataOut_payload_233_6 <= _zz_dataOut_payload_233_5;
    _zz_dataOut_payload_234_9 <= _zz_dataOut_payload_234_8;
    _zz_dataOut_payload_235_6 <= _zz_dataOut_payload_235_5;
    _zz_dataOut_payload_236_15 <= _zz_dataOut_payload_236_14;
    _zz_dataOut_payload_237_6 <= _zz_dataOut_payload_237_5;
    _zz_dataOut_payload_238_9 <= _zz_dataOut_payload_238_8;
    _zz_dataOut_payload_239_6 <= _zz_dataOut_payload_239_5;
    _zz_dataOut_payload_240_51 <= _zz_dataOut_payload_240_50;
    _zz_dataOut_payload_241_6 <= _zz_dataOut_payload_241_5;
    _zz_dataOut_payload_242_9 <= _zz_dataOut_payload_242_8;
    _zz_dataOut_payload_243_6 <= _zz_dataOut_payload_243_5;
    _zz_dataOut_payload_244_15 <= _zz_dataOut_payload_244_14;
    _zz_dataOut_payload_245_6 <= _zz_dataOut_payload_245_5;
    _zz_dataOut_payload_246_9 <= _zz_dataOut_payload_246_8;
    _zz_dataOut_payload_247_6 <= _zz_dataOut_payload_247_5;
    _zz_dataOut_payload_248_27 <= _zz_dataOut_payload_248_26;
    _zz_dataOut_payload_249_6 <= _zz_dataOut_payload_249_5;
    _zz_dataOut_payload_250_9 <= _zz_dataOut_payload_250_8;
    _zz_dataOut_payload_251_6 <= _zz_dataOut_payload_251_5;
    _zz_dataOut_payload_252_15 <= _zz_dataOut_payload_252_14;
    _zz_dataOut_payload_253_6 <= _zz_dataOut_payload_253_5;
    _zz_dataOut_payload_254_9 <= _zz_dataOut_payload_254_8;
    _zz_dataOut_payload_255_6 <= _zz_dataOut_payload_255_5;
    _zz_dataOut_payload_0_16644 <= _zz_dataOut_payload_0_16643;
    _zz_dataOut_payload_1_7 <= _zz_dataOut_payload_1_6;
    _zz_dataOut_payload_2_10 <= _zz_dataOut_payload_2_9;
    _zz_dataOut_payload_3_7 <= _zz_dataOut_payload_3_6;
    _zz_dataOut_payload_4_16 <= _zz_dataOut_payload_4_15;
    _zz_dataOut_payload_5_7 <= _zz_dataOut_payload_5_6;
    _zz_dataOut_payload_6_10 <= _zz_dataOut_payload_6_9;
    _zz_dataOut_payload_7_7 <= _zz_dataOut_payload_7_6;
    _zz_dataOut_payload_8_28 <= _zz_dataOut_payload_8_27;
    _zz_dataOut_payload_9_7 <= _zz_dataOut_payload_9_6;
    _zz_dataOut_payload_10_10 <= _zz_dataOut_payload_10_9;
    _zz_dataOut_payload_11_7 <= _zz_dataOut_payload_11_6;
    _zz_dataOut_payload_12_16 <= _zz_dataOut_payload_12_15;
    _zz_dataOut_payload_13_7 <= _zz_dataOut_payload_13_6;
    _zz_dataOut_payload_14_10 <= _zz_dataOut_payload_14_9;
    _zz_dataOut_payload_15_7 <= _zz_dataOut_payload_15_6;
    _zz_dataOut_payload_16_52 <= _zz_dataOut_payload_16_51;
    _zz_dataOut_payload_17_7 <= _zz_dataOut_payload_17_6;
    _zz_dataOut_payload_18_10 <= _zz_dataOut_payload_18_9;
    _zz_dataOut_payload_19_7 <= _zz_dataOut_payload_19_6;
    _zz_dataOut_payload_20_16 <= _zz_dataOut_payload_20_15;
    _zz_dataOut_payload_21_7 <= _zz_dataOut_payload_21_6;
    _zz_dataOut_payload_22_10 <= _zz_dataOut_payload_22_9;
    _zz_dataOut_payload_23_7 <= _zz_dataOut_payload_23_6;
    _zz_dataOut_payload_24_28 <= _zz_dataOut_payload_24_27;
    _zz_dataOut_payload_25_7 <= _zz_dataOut_payload_25_6;
    _zz_dataOut_payload_26_10 <= _zz_dataOut_payload_26_9;
    _zz_dataOut_payload_27_7 <= _zz_dataOut_payload_27_6;
    _zz_dataOut_payload_28_16 <= _zz_dataOut_payload_28_15;
    _zz_dataOut_payload_29_7 <= _zz_dataOut_payload_29_6;
    _zz_dataOut_payload_30_10 <= _zz_dataOut_payload_30_9;
    _zz_dataOut_payload_31_7 <= _zz_dataOut_payload_31_6;
    _zz_dataOut_payload_32_100 <= _zz_dataOut_payload_32_99;
    _zz_dataOut_payload_33_7 <= _zz_dataOut_payload_33_6;
    _zz_dataOut_payload_34_10 <= _zz_dataOut_payload_34_9;
    _zz_dataOut_payload_35_7 <= _zz_dataOut_payload_35_6;
    _zz_dataOut_payload_36_16 <= _zz_dataOut_payload_36_15;
    _zz_dataOut_payload_37_7 <= _zz_dataOut_payload_37_6;
    _zz_dataOut_payload_38_10 <= _zz_dataOut_payload_38_9;
    _zz_dataOut_payload_39_7 <= _zz_dataOut_payload_39_6;
    _zz_dataOut_payload_40_28 <= _zz_dataOut_payload_40_27;
    _zz_dataOut_payload_41_7 <= _zz_dataOut_payload_41_6;
    _zz_dataOut_payload_42_10 <= _zz_dataOut_payload_42_9;
    _zz_dataOut_payload_43_7 <= _zz_dataOut_payload_43_6;
    _zz_dataOut_payload_44_16 <= _zz_dataOut_payload_44_15;
    _zz_dataOut_payload_45_7 <= _zz_dataOut_payload_45_6;
    _zz_dataOut_payload_46_10 <= _zz_dataOut_payload_46_9;
    _zz_dataOut_payload_47_7 <= _zz_dataOut_payload_47_6;
    _zz_dataOut_payload_48_52 <= _zz_dataOut_payload_48_51;
    _zz_dataOut_payload_49_7 <= _zz_dataOut_payload_49_6;
    _zz_dataOut_payload_50_10 <= _zz_dataOut_payload_50_9;
    _zz_dataOut_payload_51_7 <= _zz_dataOut_payload_51_6;
    _zz_dataOut_payload_52_16 <= _zz_dataOut_payload_52_15;
    _zz_dataOut_payload_53_7 <= _zz_dataOut_payload_53_6;
    _zz_dataOut_payload_54_10 <= _zz_dataOut_payload_54_9;
    _zz_dataOut_payload_55_7 <= _zz_dataOut_payload_55_6;
    _zz_dataOut_payload_56_28 <= _zz_dataOut_payload_56_27;
    _zz_dataOut_payload_57_7 <= _zz_dataOut_payload_57_6;
    _zz_dataOut_payload_58_10 <= _zz_dataOut_payload_58_9;
    _zz_dataOut_payload_59_7 <= _zz_dataOut_payload_59_6;
    _zz_dataOut_payload_60_16 <= _zz_dataOut_payload_60_15;
    _zz_dataOut_payload_61_7 <= _zz_dataOut_payload_61_6;
    _zz_dataOut_payload_62_10 <= _zz_dataOut_payload_62_9;
    _zz_dataOut_payload_63_7 <= _zz_dataOut_payload_63_6;
    _zz_dataOut_payload_64_196 <= _zz_dataOut_payload_64_195;
    _zz_dataOut_payload_65_7 <= _zz_dataOut_payload_65_6;
    _zz_dataOut_payload_66_10 <= _zz_dataOut_payload_66_9;
    _zz_dataOut_payload_67_7 <= _zz_dataOut_payload_67_6;
    _zz_dataOut_payload_68_16 <= _zz_dataOut_payload_68_15;
    _zz_dataOut_payload_69_7 <= _zz_dataOut_payload_69_6;
    _zz_dataOut_payload_70_10 <= _zz_dataOut_payload_70_9;
    _zz_dataOut_payload_71_7 <= _zz_dataOut_payload_71_6;
    _zz_dataOut_payload_72_28 <= _zz_dataOut_payload_72_27;
    _zz_dataOut_payload_73_7 <= _zz_dataOut_payload_73_6;
    _zz_dataOut_payload_74_10 <= _zz_dataOut_payload_74_9;
    _zz_dataOut_payload_75_7 <= _zz_dataOut_payload_75_6;
    _zz_dataOut_payload_76_16 <= _zz_dataOut_payload_76_15;
    _zz_dataOut_payload_77_7 <= _zz_dataOut_payload_77_6;
    _zz_dataOut_payload_78_10 <= _zz_dataOut_payload_78_9;
    _zz_dataOut_payload_79_7 <= _zz_dataOut_payload_79_6;
    _zz_dataOut_payload_80_52 <= _zz_dataOut_payload_80_51;
    _zz_dataOut_payload_81_7 <= _zz_dataOut_payload_81_6;
    _zz_dataOut_payload_82_10 <= _zz_dataOut_payload_82_9;
    _zz_dataOut_payload_83_7 <= _zz_dataOut_payload_83_6;
    _zz_dataOut_payload_84_16 <= _zz_dataOut_payload_84_15;
    _zz_dataOut_payload_85_7 <= _zz_dataOut_payload_85_6;
    _zz_dataOut_payload_86_10 <= _zz_dataOut_payload_86_9;
    _zz_dataOut_payload_87_7 <= _zz_dataOut_payload_87_6;
    _zz_dataOut_payload_88_28 <= _zz_dataOut_payload_88_27;
    _zz_dataOut_payload_89_7 <= _zz_dataOut_payload_89_6;
    _zz_dataOut_payload_90_10 <= _zz_dataOut_payload_90_9;
    _zz_dataOut_payload_91_7 <= _zz_dataOut_payload_91_6;
    _zz_dataOut_payload_92_16 <= _zz_dataOut_payload_92_15;
    _zz_dataOut_payload_93_7 <= _zz_dataOut_payload_93_6;
    _zz_dataOut_payload_94_10 <= _zz_dataOut_payload_94_9;
    _zz_dataOut_payload_95_7 <= _zz_dataOut_payload_95_6;
    _zz_dataOut_payload_96_100 <= _zz_dataOut_payload_96_99;
    _zz_dataOut_payload_97_7 <= _zz_dataOut_payload_97_6;
    _zz_dataOut_payload_98_10 <= _zz_dataOut_payload_98_9;
    _zz_dataOut_payload_99_7 <= _zz_dataOut_payload_99_6;
    _zz_dataOut_payload_100_16 <= _zz_dataOut_payload_100_15;
    _zz_dataOut_payload_101_7 <= _zz_dataOut_payload_101_6;
    _zz_dataOut_payload_102_10 <= _zz_dataOut_payload_102_9;
    _zz_dataOut_payload_103_7 <= _zz_dataOut_payload_103_6;
    _zz_dataOut_payload_104_28 <= _zz_dataOut_payload_104_27;
    _zz_dataOut_payload_105_7 <= _zz_dataOut_payload_105_6;
    _zz_dataOut_payload_106_10 <= _zz_dataOut_payload_106_9;
    _zz_dataOut_payload_107_7 <= _zz_dataOut_payload_107_6;
    _zz_dataOut_payload_108_16 <= _zz_dataOut_payload_108_15;
    _zz_dataOut_payload_109_7 <= _zz_dataOut_payload_109_6;
    _zz_dataOut_payload_110_10 <= _zz_dataOut_payload_110_9;
    _zz_dataOut_payload_111_7 <= _zz_dataOut_payload_111_6;
    _zz_dataOut_payload_112_52 <= _zz_dataOut_payload_112_51;
    _zz_dataOut_payload_113_7 <= _zz_dataOut_payload_113_6;
    _zz_dataOut_payload_114_10 <= _zz_dataOut_payload_114_9;
    _zz_dataOut_payload_115_7 <= _zz_dataOut_payload_115_6;
    _zz_dataOut_payload_116_16 <= _zz_dataOut_payload_116_15;
    _zz_dataOut_payload_117_7 <= _zz_dataOut_payload_117_6;
    _zz_dataOut_payload_118_10 <= _zz_dataOut_payload_118_9;
    _zz_dataOut_payload_119_7 <= _zz_dataOut_payload_119_6;
    _zz_dataOut_payload_120_28 <= _zz_dataOut_payload_120_27;
    _zz_dataOut_payload_121_7 <= _zz_dataOut_payload_121_6;
    _zz_dataOut_payload_122_10 <= _zz_dataOut_payload_122_9;
    _zz_dataOut_payload_123_7 <= _zz_dataOut_payload_123_6;
    _zz_dataOut_payload_124_16 <= _zz_dataOut_payload_124_15;
    _zz_dataOut_payload_125_7 <= _zz_dataOut_payload_125_6;
    _zz_dataOut_payload_126_10 <= _zz_dataOut_payload_126_9;
    _zz_dataOut_payload_127_7 <= _zz_dataOut_payload_127_6;
    _zz_dataOut_payload_128_388 <= _zz_dataOut_payload_128_387;
    _zz_dataOut_payload_129_7 <= _zz_dataOut_payload_129_6;
    _zz_dataOut_payload_130_10 <= _zz_dataOut_payload_130_9;
    _zz_dataOut_payload_131_7 <= _zz_dataOut_payload_131_6;
    _zz_dataOut_payload_132_16 <= _zz_dataOut_payload_132_15;
    _zz_dataOut_payload_133_7 <= _zz_dataOut_payload_133_6;
    _zz_dataOut_payload_134_10 <= _zz_dataOut_payload_134_9;
    _zz_dataOut_payload_135_7 <= _zz_dataOut_payload_135_6;
    _zz_dataOut_payload_136_28 <= _zz_dataOut_payload_136_27;
    _zz_dataOut_payload_137_7 <= _zz_dataOut_payload_137_6;
    _zz_dataOut_payload_138_10 <= _zz_dataOut_payload_138_9;
    _zz_dataOut_payload_139_7 <= _zz_dataOut_payload_139_6;
    _zz_dataOut_payload_140_16 <= _zz_dataOut_payload_140_15;
    _zz_dataOut_payload_141_7 <= _zz_dataOut_payload_141_6;
    _zz_dataOut_payload_142_10 <= _zz_dataOut_payload_142_9;
    _zz_dataOut_payload_143_7 <= _zz_dataOut_payload_143_6;
    _zz_dataOut_payload_144_52 <= _zz_dataOut_payload_144_51;
    _zz_dataOut_payload_145_7 <= _zz_dataOut_payload_145_6;
    _zz_dataOut_payload_146_10 <= _zz_dataOut_payload_146_9;
    _zz_dataOut_payload_147_7 <= _zz_dataOut_payload_147_6;
    _zz_dataOut_payload_148_16 <= _zz_dataOut_payload_148_15;
    _zz_dataOut_payload_149_7 <= _zz_dataOut_payload_149_6;
    _zz_dataOut_payload_150_10 <= _zz_dataOut_payload_150_9;
    _zz_dataOut_payload_151_7 <= _zz_dataOut_payload_151_6;
    _zz_dataOut_payload_152_28 <= _zz_dataOut_payload_152_27;
    _zz_dataOut_payload_153_7 <= _zz_dataOut_payload_153_6;
    _zz_dataOut_payload_154_10 <= _zz_dataOut_payload_154_9;
    _zz_dataOut_payload_155_7 <= _zz_dataOut_payload_155_6;
    _zz_dataOut_payload_156_16 <= _zz_dataOut_payload_156_15;
    _zz_dataOut_payload_157_7 <= _zz_dataOut_payload_157_6;
    _zz_dataOut_payload_158_10 <= _zz_dataOut_payload_158_9;
    _zz_dataOut_payload_159_7 <= _zz_dataOut_payload_159_6;
    _zz_dataOut_payload_160_100 <= _zz_dataOut_payload_160_99;
    _zz_dataOut_payload_161_7 <= _zz_dataOut_payload_161_6;
    _zz_dataOut_payload_162_10 <= _zz_dataOut_payload_162_9;
    _zz_dataOut_payload_163_7 <= _zz_dataOut_payload_163_6;
    _zz_dataOut_payload_164_16 <= _zz_dataOut_payload_164_15;
    _zz_dataOut_payload_165_7 <= _zz_dataOut_payload_165_6;
    _zz_dataOut_payload_166_10 <= _zz_dataOut_payload_166_9;
    _zz_dataOut_payload_167_7 <= _zz_dataOut_payload_167_6;
    _zz_dataOut_payload_168_28 <= _zz_dataOut_payload_168_27;
    _zz_dataOut_payload_169_7 <= _zz_dataOut_payload_169_6;
    _zz_dataOut_payload_170_10 <= _zz_dataOut_payload_170_9;
    _zz_dataOut_payload_171_7 <= _zz_dataOut_payload_171_6;
    _zz_dataOut_payload_172_16 <= _zz_dataOut_payload_172_15;
    _zz_dataOut_payload_173_7 <= _zz_dataOut_payload_173_6;
    _zz_dataOut_payload_174_10 <= _zz_dataOut_payload_174_9;
    _zz_dataOut_payload_175_7 <= _zz_dataOut_payload_175_6;
    _zz_dataOut_payload_176_52 <= _zz_dataOut_payload_176_51;
    _zz_dataOut_payload_177_7 <= _zz_dataOut_payload_177_6;
    _zz_dataOut_payload_178_10 <= _zz_dataOut_payload_178_9;
    _zz_dataOut_payload_179_7 <= _zz_dataOut_payload_179_6;
    _zz_dataOut_payload_180_16 <= _zz_dataOut_payload_180_15;
    _zz_dataOut_payload_181_7 <= _zz_dataOut_payload_181_6;
    _zz_dataOut_payload_182_10 <= _zz_dataOut_payload_182_9;
    _zz_dataOut_payload_183_7 <= _zz_dataOut_payload_183_6;
    _zz_dataOut_payload_184_28 <= _zz_dataOut_payload_184_27;
    _zz_dataOut_payload_185_7 <= _zz_dataOut_payload_185_6;
    _zz_dataOut_payload_186_10 <= _zz_dataOut_payload_186_9;
    _zz_dataOut_payload_187_7 <= _zz_dataOut_payload_187_6;
    _zz_dataOut_payload_188_16 <= _zz_dataOut_payload_188_15;
    _zz_dataOut_payload_189_7 <= _zz_dataOut_payload_189_6;
    _zz_dataOut_payload_190_10 <= _zz_dataOut_payload_190_9;
    _zz_dataOut_payload_191_7 <= _zz_dataOut_payload_191_6;
    _zz_dataOut_payload_192_196 <= _zz_dataOut_payload_192_195;
    _zz_dataOut_payload_193_7 <= _zz_dataOut_payload_193_6;
    _zz_dataOut_payload_194_10 <= _zz_dataOut_payload_194_9;
    _zz_dataOut_payload_195_7 <= _zz_dataOut_payload_195_6;
    _zz_dataOut_payload_196_16 <= _zz_dataOut_payload_196_15;
    _zz_dataOut_payload_197_7 <= _zz_dataOut_payload_197_6;
    _zz_dataOut_payload_198_10 <= _zz_dataOut_payload_198_9;
    _zz_dataOut_payload_199_7 <= _zz_dataOut_payload_199_6;
    _zz_dataOut_payload_200_28 <= _zz_dataOut_payload_200_27;
    _zz_dataOut_payload_201_7 <= _zz_dataOut_payload_201_6;
    _zz_dataOut_payload_202_10 <= _zz_dataOut_payload_202_9;
    _zz_dataOut_payload_203_7 <= _zz_dataOut_payload_203_6;
    _zz_dataOut_payload_204_16 <= _zz_dataOut_payload_204_15;
    _zz_dataOut_payload_205_7 <= _zz_dataOut_payload_205_6;
    _zz_dataOut_payload_206_10 <= _zz_dataOut_payload_206_9;
    _zz_dataOut_payload_207_7 <= _zz_dataOut_payload_207_6;
    _zz_dataOut_payload_208_52 <= _zz_dataOut_payload_208_51;
    _zz_dataOut_payload_209_7 <= _zz_dataOut_payload_209_6;
    _zz_dataOut_payload_210_10 <= _zz_dataOut_payload_210_9;
    _zz_dataOut_payload_211_7 <= _zz_dataOut_payload_211_6;
    _zz_dataOut_payload_212_16 <= _zz_dataOut_payload_212_15;
    _zz_dataOut_payload_213_7 <= _zz_dataOut_payload_213_6;
    _zz_dataOut_payload_214_10 <= _zz_dataOut_payload_214_9;
    _zz_dataOut_payload_215_7 <= _zz_dataOut_payload_215_6;
    _zz_dataOut_payload_216_28 <= _zz_dataOut_payload_216_27;
    _zz_dataOut_payload_217_7 <= _zz_dataOut_payload_217_6;
    _zz_dataOut_payload_218_10 <= _zz_dataOut_payload_218_9;
    _zz_dataOut_payload_219_7 <= _zz_dataOut_payload_219_6;
    _zz_dataOut_payload_220_16 <= _zz_dataOut_payload_220_15;
    _zz_dataOut_payload_221_7 <= _zz_dataOut_payload_221_6;
    _zz_dataOut_payload_222_10 <= _zz_dataOut_payload_222_9;
    _zz_dataOut_payload_223_7 <= _zz_dataOut_payload_223_6;
    _zz_dataOut_payload_224_100 <= _zz_dataOut_payload_224_99;
    _zz_dataOut_payload_225_7 <= _zz_dataOut_payload_225_6;
    _zz_dataOut_payload_226_10 <= _zz_dataOut_payload_226_9;
    _zz_dataOut_payload_227_7 <= _zz_dataOut_payload_227_6;
    _zz_dataOut_payload_228_16 <= _zz_dataOut_payload_228_15;
    _zz_dataOut_payload_229_7 <= _zz_dataOut_payload_229_6;
    _zz_dataOut_payload_230_10 <= _zz_dataOut_payload_230_9;
    _zz_dataOut_payload_231_7 <= _zz_dataOut_payload_231_6;
    _zz_dataOut_payload_232_28 <= _zz_dataOut_payload_232_27;
    _zz_dataOut_payload_233_7 <= _zz_dataOut_payload_233_6;
    _zz_dataOut_payload_234_10 <= _zz_dataOut_payload_234_9;
    _zz_dataOut_payload_235_7 <= _zz_dataOut_payload_235_6;
    _zz_dataOut_payload_236_16 <= _zz_dataOut_payload_236_15;
    _zz_dataOut_payload_237_7 <= _zz_dataOut_payload_237_6;
    _zz_dataOut_payload_238_10 <= _zz_dataOut_payload_238_9;
    _zz_dataOut_payload_239_7 <= _zz_dataOut_payload_239_6;
    _zz_dataOut_payload_240_52 <= _zz_dataOut_payload_240_51;
    _zz_dataOut_payload_241_7 <= _zz_dataOut_payload_241_6;
    _zz_dataOut_payload_242_10 <= _zz_dataOut_payload_242_9;
    _zz_dataOut_payload_243_7 <= _zz_dataOut_payload_243_6;
    _zz_dataOut_payload_244_16 <= _zz_dataOut_payload_244_15;
    _zz_dataOut_payload_245_7 <= _zz_dataOut_payload_245_6;
    _zz_dataOut_payload_246_10 <= _zz_dataOut_payload_246_9;
    _zz_dataOut_payload_247_7 <= _zz_dataOut_payload_247_6;
    _zz_dataOut_payload_248_28 <= _zz_dataOut_payload_248_27;
    _zz_dataOut_payload_249_7 <= _zz_dataOut_payload_249_6;
    _zz_dataOut_payload_250_10 <= _zz_dataOut_payload_250_9;
    _zz_dataOut_payload_251_7 <= _zz_dataOut_payload_251_6;
    _zz_dataOut_payload_252_16 <= _zz_dataOut_payload_252_15;
    _zz_dataOut_payload_253_7 <= _zz_dataOut_payload_253_6;
    _zz_dataOut_payload_254_10 <= _zz_dataOut_payload_254_9;
    _zz_dataOut_payload_255_7 <= _zz_dataOut_payload_255_6;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      dataIn_valid_delay_1 <= 1'b0;
      dataIn_valid_delay_2 <= 1'b0;
      dataIn_valid_delay_3 <= 1'b0;
      dataIn_valid_delay_4 <= 1'b0;
      dataIn_valid_delay_5 <= 1'b0;
      dataIn_valid_delay_6 <= 1'b0;
      dataIn_valid_delay_7 <= 1'b0;
      dataIn_valid_delay_8 <= 1'b0;
      dataIn_valid_delay_9 <= 1'b0;
      dataIn_valid_delay_10 <= 1'b0;
      dataIn_valid_delay_11 <= 1'b0;
      dataIn_valid_delay_12 <= 1'b0;
      dataIn_valid_delay_13 <= 1'b0;
      dataIn_valid_delay_14 <= 1'b0;
      dataIn_valid_delay_15 <= 1'b0;
      dataIn_valid_delay_16 <= 1'b0;
      dataIn_valid_delay_17 <= 1'b0;
      dataIn_valid_delay_18 <= 1'b0;
      dataIn_valid_delay_19 <= 1'b0;
      dataIn_valid_delay_20 <= 1'b0;
      dataIn_valid_delay_21 <= 1'b0;
      dataIn_valid_delay_22 <= 1'b0;
      dataIn_valid_delay_23 <= 1'b0;
      dataIn_valid_delay_24 <= 1'b0;
      dataIn_valid_delay_25 <= 1'b0;
      dataIn_valid_delay_26 <= 1'b0;
      dataIn_valid_delay_27 <= 1'b0;
      dataIn_valid_delay_28 <= 1'b0;
      dataIn_valid_delay_29 <= 1'b0;
      dataIn_valid_delay_30 <= 1'b0;
      dataIn_valid_delay_31 <= 1'b0;
      dataIn_valid_delay_32 <= 1'b0;
      dataIn_valid_delay_33 <= 1'b0;
      dataIn_valid_delay_34 <= 1'b0;
      dataIn_valid_delay_35 <= 1'b0;
      dataIn_valid_delay_36 <= 1'b0;
    end else begin
      dataIn_valid_delay_1 <= dataIn_valid;
      dataIn_valid_delay_2 <= dataIn_valid_delay_1;
      dataIn_valid_delay_3 <= dataIn_valid_delay_2;
      dataIn_valid_delay_4 <= dataIn_valid_delay_3;
      dataIn_valid_delay_5 <= dataIn_valid_delay_4;
      dataIn_valid_delay_6 <= dataIn_valid_delay_5;
      dataIn_valid_delay_7 <= dataIn_valid_delay_6;
      dataIn_valid_delay_8 <= dataIn_valid_delay_7;
      dataIn_valid_delay_9 <= dataIn_valid_delay_8;
      dataIn_valid_delay_10 <= dataIn_valid_delay_9;
      dataIn_valid_delay_11 <= dataIn_valid_delay_10;
      dataIn_valid_delay_12 <= dataIn_valid_delay_11;
      dataIn_valid_delay_13 <= dataIn_valid_delay_12;
      dataIn_valid_delay_14 <= dataIn_valid_delay_13;
      dataIn_valid_delay_15 <= dataIn_valid_delay_14;
      dataIn_valid_delay_16 <= dataIn_valid_delay_15;
      dataIn_valid_delay_17 <= dataIn_valid_delay_16;
      dataIn_valid_delay_18 <= dataIn_valid_delay_17;
      dataIn_valid_delay_19 <= dataIn_valid_delay_18;
      dataIn_valid_delay_20 <= dataIn_valid_delay_19;
      dataIn_valid_delay_21 <= dataIn_valid_delay_20;
      dataIn_valid_delay_22 <= dataIn_valid_delay_21;
      dataIn_valid_delay_23 <= dataIn_valid_delay_22;
      dataIn_valid_delay_24 <= dataIn_valid_delay_23;
      dataIn_valid_delay_25 <= dataIn_valid_delay_24;
      dataIn_valid_delay_26 <= dataIn_valid_delay_25;
      dataIn_valid_delay_27 <= dataIn_valid_delay_26;
      dataIn_valid_delay_28 <= dataIn_valid_delay_27;
      dataIn_valid_delay_29 <= dataIn_valid_delay_28;
      dataIn_valid_delay_30 <= dataIn_valid_delay_29;
      dataIn_valid_delay_31 <= dataIn_valid_delay_30;
      dataIn_valid_delay_32 <= dataIn_valid_delay_31;
      dataIn_valid_delay_33 <= dataIn_valid_delay_32;
      dataIn_valid_delay_34 <= dataIn_valid_delay_33;
      dataIn_valid_delay_35 <= dataIn_valid_delay_34;
      dataIn_valid_delay_36 <= dataIn_valid_delay_35;
    end
  end


endmodule
